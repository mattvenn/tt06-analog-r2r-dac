magic
tech sky130A
magscale 1 2
timestamp 1708507682
<< viali >>
rect 4905 15113 4939 15147
rect 8861 15113 8895 15147
rect 2513 15045 2547 15079
rect 1225 14977 1259 15011
rect 1041 14909 1075 14943
rect 2329 14909 2363 14943
rect 3525 14909 3559 14943
rect 4905 14909 4939 14943
rect 5181 14909 5215 14943
rect 5273 14909 5307 14943
rect 6101 14909 6135 14943
rect 7389 14909 7423 14943
rect 8677 14909 8711 14943
rect 8953 14909 8987 14943
rect 9045 14909 9079 14943
rect 9965 14909 9999 14943
rect 11253 14909 11287 14943
rect 12725 14909 12759 14943
rect 13829 14909 13863 14943
rect 3709 14773 3743 14807
rect 4629 14773 4663 14807
rect 5457 14773 5491 14807
rect 6285 14773 6319 14807
rect 7573 14773 7607 14807
rect 8401 14773 8435 14807
rect 9229 14773 9263 14807
rect 10149 14773 10183 14807
rect 11437 14773 11471 14807
rect 12541 14773 12575 14807
rect 12817 14773 12851 14807
rect 14013 14773 14047 14807
rect 5825 14569 5859 14603
rect 8125 14569 8159 14603
rect 12725 14501 12759 14535
rect 4833 14433 4867 14467
rect 5089 14433 5123 14467
rect 5457 14433 5491 14467
rect 6938 14433 6972 14467
rect 7205 14433 7239 14467
rect 7573 14433 7607 14467
rect 7849 14433 7883 14467
rect 9238 14433 9272 14467
rect 10793 14433 10827 14467
rect 12090 14433 12124 14467
rect 12357 14433 12391 14467
rect 12449 14433 12483 14467
rect 14381 14433 14415 14467
rect 9505 14365 9539 14399
rect 10149 14365 10183 14399
rect 10517 14365 10551 14399
rect 10609 14365 10643 14399
rect 14473 14365 14507 14399
rect 3709 14229 3743 14263
rect 5273 14229 5307 14263
rect 7297 14229 7331 14263
rect 7481 14229 7515 14263
rect 10977 14229 11011 14263
rect 14197 14229 14231 14263
rect 4997 14025 5031 14059
rect 7021 14025 7055 14059
rect 9229 14025 9263 14059
rect 10425 14025 10459 14059
rect 10885 14025 10919 14059
rect 11253 14025 11287 14059
rect 12909 13957 12943 13991
rect 4353 13889 4387 13923
rect 6377 13889 6411 13923
rect 8585 13889 8619 13923
rect 4721 13821 4755 13855
rect 4813 13821 4847 13855
rect 6745 13821 6779 13855
rect 6837 13821 6871 13855
rect 8953 13821 8987 13855
rect 9045 13821 9079 13855
rect 10609 13821 10643 13855
rect 10971 13821 11005 13855
rect 11897 13821 11931 13855
rect 12081 13821 12115 13855
rect 12173 13821 12207 13855
rect 12357 13821 12391 13855
rect 12633 13821 12667 13855
rect 14473 13821 14507 13855
rect 14565 13821 14599 13855
rect 11529 13753 11563 13787
rect 11989 13753 12023 13787
rect 12725 13753 12759 13787
rect 12909 13753 12943 13787
rect 12265 13685 12299 13719
rect 13829 13685 13863 13719
rect 14657 13685 14691 13719
rect 12173 13481 12207 13515
rect 12725 13481 12759 13515
rect 14933 13481 14967 13515
rect 4353 13345 4387 13379
rect 6101 13345 6135 13379
rect 8329 13345 8363 13379
rect 9312 13345 9346 13379
rect 11667 13345 11701 13379
rect 11805 13345 11839 13379
rect 11897 13345 11931 13379
rect 11989 13345 12023 13379
rect 12449 13345 12483 13379
rect 13369 13345 13403 13379
rect 3893 13277 3927 13311
rect 4261 13277 4295 13311
rect 6009 13277 6043 13311
rect 6469 13277 6503 13311
rect 8585 13277 8619 13311
rect 9045 13277 9079 13311
rect 11529 13277 11563 13311
rect 12725 13277 12759 13311
rect 13645 13277 13679 13311
rect 4537 13141 4571 13175
rect 5825 13141 5859 13175
rect 7205 13141 7239 13175
rect 10425 13141 10459 13175
rect 12541 13141 12575 13175
rect 6745 12937 6779 12971
rect 7113 12937 7147 12971
rect 7757 12937 7791 12971
rect 9045 12937 9079 12971
rect 9965 12937 9999 12971
rect 10885 12937 10919 12971
rect 12725 12869 12759 12903
rect 4629 12801 4663 12835
rect 5273 12801 5307 12835
rect 7021 12801 7055 12835
rect 7941 12801 7975 12835
rect 8769 12801 8803 12835
rect 10241 12801 10275 12835
rect 4373 12733 4407 12767
rect 5540 12733 5574 12767
rect 7107 12733 7141 12767
rect 7205 12733 7239 12767
rect 7665 12733 7699 12767
rect 8861 12733 8895 12767
rect 10149 12733 10183 12767
rect 10885 12733 10919 12767
rect 11253 12733 11287 12767
rect 11345 12733 11379 12767
rect 11529 12733 11563 12767
rect 11805 12733 11839 12767
rect 11989 12733 12023 12767
rect 12081 12733 12115 12767
rect 12173 12733 12207 12767
rect 12449 12733 12483 12767
rect 12541 12733 12575 12767
rect 13185 12733 13219 12767
rect 13829 12733 13863 12767
rect 13921 12733 13955 12767
rect 14013 12733 14047 12767
rect 14197 12733 14231 12767
rect 11713 12665 11747 12699
rect 12357 12665 12391 12699
rect 12817 12665 12851 12699
rect 13001 12665 13035 12699
rect 3249 12597 3283 12631
rect 6653 12597 6687 12631
rect 7297 12597 7331 12631
rect 8217 12597 8251 12631
rect 8401 12597 8435 12631
rect 10609 12597 10643 12631
rect 10701 12597 10735 12631
rect 11897 12597 11931 12631
rect 13553 12597 13587 12631
rect 4261 12393 4295 12427
rect 12633 12393 12667 12427
rect 15025 12325 15059 12359
rect 4537 12257 4571 12291
rect 4813 12257 4847 12291
rect 7849 12257 7883 12291
rect 8125 12257 8159 12291
rect 8217 12257 8251 12291
rect 12449 12257 12483 12291
rect 13369 12257 13403 12291
rect 13645 12257 13679 12291
rect 7941 12189 7975 12223
rect 8493 12189 8527 12223
rect 9505 12189 9539 12223
rect 12265 12189 12299 12223
rect 8769 12121 8803 12155
rect 9873 12121 9907 12155
rect 4721 12053 4755 12087
rect 8401 12053 8435 12087
rect 8953 12053 8987 12087
rect 9965 12053 9999 12087
rect 12725 11849 12759 11883
rect 12909 11849 12943 11883
rect 6653 11781 6687 11815
rect 3893 11713 3927 11747
rect 4353 11713 4387 11747
rect 8125 11713 8159 11747
rect 9689 11713 9723 11747
rect 11713 11713 11747 11747
rect 3985 11645 4019 11679
rect 5089 11645 5123 11679
rect 5273 11645 5307 11679
rect 5365 11645 5399 11679
rect 5457 11645 5491 11679
rect 6837 11645 6871 11679
rect 6985 11645 7019 11679
rect 7113 11645 7147 11679
rect 7343 11645 7377 11679
rect 7757 11645 7791 11679
rect 7849 11645 7883 11679
rect 8723 11645 8757 11679
rect 9136 11645 9170 11679
rect 9229 11645 9263 11679
rect 12081 11645 12115 11679
rect 12265 11645 12299 11679
rect 13829 11645 13863 11679
rect 13921 11645 13955 11679
rect 14013 11645 14047 11679
rect 14197 11645 14231 11679
rect 6285 11577 6319 11611
rect 7205 11577 7239 11611
rect 8217 11577 8251 11611
rect 8861 11577 8895 11611
rect 8953 11577 8987 11611
rect 9934 11577 9968 11611
rect 13093 11577 13127 11611
rect 5733 11509 5767 11543
rect 6745 11509 6779 11543
rect 7481 11509 7515 11543
rect 7573 11509 7607 11543
rect 8585 11509 8619 11543
rect 11069 11509 11103 11543
rect 11161 11509 11195 11543
rect 12173 11509 12207 11543
rect 12893 11509 12927 11543
rect 13553 11509 13587 11543
rect 4261 11305 4295 11339
rect 4813 11305 4847 11339
rect 7757 11305 7791 11339
rect 8953 11305 8987 11339
rect 9689 11305 9723 11339
rect 11897 11305 11931 11339
rect 13001 11305 13035 11339
rect 10517 11237 10551 11271
rect 3801 11169 3835 11203
rect 4353 11169 4387 11203
rect 4905 11169 4939 11203
rect 5917 11169 5951 11203
rect 6009 11169 6043 11203
rect 6193 11169 6227 11203
rect 6653 11169 6687 11203
rect 6745 11169 6779 11203
rect 7021 11169 7055 11203
rect 7389 11169 7423 11203
rect 7849 11169 7883 11203
rect 8493 11169 8527 11203
rect 9873 11169 9907 11203
rect 10149 11169 10183 11203
rect 10333 11169 10367 11203
rect 10609 11169 10643 11203
rect 12357 11169 12391 11203
rect 12450 11169 12484 11203
rect 12633 11169 12667 11203
rect 12725 11169 12759 11203
rect 12822 11169 12856 11203
rect 13369 11169 13403 11203
rect 13645 11169 13679 11203
rect 5181 11101 5215 11135
rect 11621 11101 11655 11135
rect 11805 11101 11839 11135
rect 5457 11033 5491 11067
rect 6101 11033 6135 11067
rect 6469 11033 6503 11067
rect 6929 11033 6963 11067
rect 7481 11033 7515 11067
rect 9965 11033 9999 11067
rect 10057 11033 10091 11067
rect 3893 10965 3927 10999
rect 4629 10965 4663 10999
rect 4997 10965 5031 10999
rect 6377 10965 6411 10999
rect 7113 10965 7147 10999
rect 7573 10965 7607 10999
rect 8769 10965 8803 10999
rect 12265 10965 12299 10999
rect 14933 10965 14967 10999
rect 4997 10761 5031 10795
rect 5549 10761 5583 10795
rect 10333 10761 10367 10795
rect 12633 10761 12667 10795
rect 13277 10761 13311 10795
rect 4813 10693 4847 10727
rect 4537 10625 4571 10659
rect 9965 10625 9999 10659
rect 10057 10625 10091 10659
rect 9873 10557 9907 10591
rect 10149 10557 10183 10591
rect 12817 10557 12851 10591
rect 13093 10557 13127 10591
rect 13185 10557 13219 10591
rect 13369 10557 13403 10591
rect 7021 10489 7055 10523
rect 10425 10489 10459 10523
rect 12173 10489 12207 10523
rect 13001 10421 13035 10455
rect 7389 10217 7423 10251
rect 7665 10217 7699 10251
rect 8585 10217 8619 10251
rect 9873 10217 9907 10251
rect 11437 10217 11471 10251
rect 5917 10149 5951 10183
rect 6469 10149 6503 10183
rect 11345 10149 11379 10183
rect 5181 10081 5215 10115
rect 5365 10081 5399 10115
rect 6561 10081 6595 10115
rect 7481 10081 7515 10115
rect 7757 10081 7791 10115
rect 8493 10081 8527 10115
rect 8769 10081 8803 10115
rect 9045 10081 9079 10115
rect 9229 10081 9263 10115
rect 9321 10081 9355 10115
rect 9413 10081 9447 10115
rect 9781 10081 9815 10115
rect 10057 10081 10091 10115
rect 12265 10081 12299 10115
rect 12449 10081 12483 10115
rect 12817 10081 12851 10115
rect 13081 10081 13115 10115
rect 13185 10081 13219 10115
rect 13277 10081 13311 10115
rect 8953 10013 8987 10047
rect 12541 10013 12575 10047
rect 12633 10013 12667 10047
rect 13369 10013 13403 10047
rect 13645 10013 13679 10047
rect 9689 9945 9723 9979
rect 13001 9945 13035 9979
rect 5365 9877 5399 9911
rect 6193 9877 6227 9911
rect 10057 9877 10091 9911
rect 14933 9877 14967 9911
rect 6745 9673 6779 9707
rect 7573 9673 7607 9707
rect 7757 9673 7791 9707
rect 8585 9673 8619 9707
rect 9321 9673 9355 9707
rect 11345 9673 11379 9707
rect 13369 9673 13403 9707
rect 6285 9605 6319 9639
rect 8769 9605 8803 9639
rect 13093 9605 13127 9639
rect 4905 9537 4939 9571
rect 7113 9537 7147 9571
rect 10701 9537 10735 9571
rect 5172 9469 5206 9503
rect 6929 9469 6963 9503
rect 7021 9469 7055 9503
rect 7205 9469 7239 9503
rect 7389 9469 7423 9503
rect 10434 9469 10468 9503
rect 10793 9469 10827 9503
rect 10977 9469 11011 9503
rect 11161 9469 11195 9503
rect 12449 9469 12483 9503
rect 12597 9469 12631 9503
rect 12725 9469 12759 9503
rect 12817 9469 12851 9503
rect 12914 9469 12948 9503
rect 13185 9469 13219 9503
rect 13369 9469 13403 9503
rect 13829 9469 13863 9503
rect 13921 9469 13955 9503
rect 14013 9469 14047 9503
rect 14197 9469 14231 9503
rect 7941 9401 7975 9435
rect 8401 9401 8435 9435
rect 7731 9333 7765 9367
rect 8611 9333 8645 9367
rect 10977 9333 11011 9367
rect 13553 9333 13587 9367
rect 6837 9129 6871 9163
rect 7665 9129 7699 9163
rect 11621 9129 11655 9163
rect 7297 9061 7331 9095
rect 10241 9061 10275 9095
rect 12725 9061 12759 9095
rect 4925 8993 4959 9027
rect 5181 8993 5215 9027
rect 5273 8993 5307 9027
rect 5457 8993 5491 9027
rect 6193 8993 6227 9027
rect 6377 8993 6411 9027
rect 6653 8993 6687 9027
rect 6745 8993 6779 9027
rect 7113 8993 7147 9027
rect 7389 8993 7423 9027
rect 7573 8993 7607 9027
rect 11252 8993 11286 9027
rect 11345 8993 11379 9027
rect 11897 8993 11931 9027
rect 11989 8993 12023 9027
rect 12357 8993 12391 9027
rect 12541 8993 12575 9027
rect 13369 8993 13403 9027
rect 13645 8993 13679 9027
rect 5365 8925 5399 8959
rect 6009 8925 6043 8959
rect 6469 8925 6503 8959
rect 11069 8925 11103 8959
rect 11161 8925 11195 8959
rect 6285 8857 6319 8891
rect 7113 8857 7147 8891
rect 3801 8789 3835 8823
rect 8953 8789 8987 8823
rect 11529 8789 11563 8823
rect 11805 8789 11839 8823
rect 14933 8789 14967 8823
rect 6193 8585 6227 8619
rect 11805 8585 11839 8619
rect 11989 8585 12023 8619
rect 12173 8585 12207 8619
rect 13277 8585 13311 8619
rect 9413 8517 9447 8551
rect 7757 8449 7791 8483
rect 12725 8449 12759 8483
rect 4537 8381 4571 8415
rect 5917 8381 5951 8415
rect 6193 8381 6227 8415
rect 7113 8381 7147 8415
rect 7297 8381 7331 8415
rect 7389 8381 7423 8415
rect 7573 8381 7607 8415
rect 8401 8381 8435 8415
rect 8559 8381 8593 8415
rect 8861 8381 8895 8415
rect 9137 8381 9171 8415
rect 9321 8381 9355 8415
rect 10793 8381 10827 8415
rect 11529 8381 11563 8415
rect 11621 8381 11655 8415
rect 13737 8381 13771 8415
rect 14013 8381 14047 8415
rect 14197 8381 14231 8415
rect 14381 8381 14415 8415
rect 14933 8381 14967 8415
rect 7849 8313 7883 8347
rect 8033 8313 8067 8347
rect 8677 8313 8711 8347
rect 8769 8313 8803 8347
rect 9229 8313 9263 8347
rect 10526 8313 10560 8347
rect 11805 8313 11839 8347
rect 12357 8313 12391 8347
rect 12909 8313 12943 8347
rect 5181 8245 5215 8279
rect 6009 8245 6043 8279
rect 7297 8245 7331 8279
rect 8217 8245 8251 8279
rect 9045 8245 9079 8279
rect 12157 8245 12191 8279
rect 13001 8245 13035 8279
rect 13093 8245 13127 8279
rect 13553 8245 13587 8279
rect 3525 8041 3559 8075
rect 6929 8041 6963 8075
rect 9689 8041 9723 8075
rect 4660 7973 4694 8007
rect 5181 7973 5215 8007
rect 5457 7973 5491 8007
rect 6745 7973 6779 8007
rect 7021 7973 7055 8007
rect 11621 7973 11655 8007
rect 12173 7973 12207 8007
rect 4997 7905 5031 7939
rect 5273 7905 5307 7939
rect 5365 7905 5399 7939
rect 5549 7905 5583 7939
rect 6009 7905 6043 7939
rect 6101 7905 6135 7939
rect 6285 7905 6319 7939
rect 6377 7905 6411 7939
rect 6469 7905 6503 7939
rect 6653 7905 6687 7939
rect 7113 7905 7147 7939
rect 9229 7905 9263 7939
rect 9413 7905 9447 7939
rect 9505 7905 9539 7939
rect 11437 7905 11471 7939
rect 11713 7905 11747 7939
rect 11805 7905 11839 7939
rect 12081 7905 12115 7939
rect 12265 7905 12299 7939
rect 13645 7905 13679 7939
rect 4905 7837 4939 7871
rect 5825 7837 5859 7871
rect 6561 7837 6595 7871
rect 9045 7837 9079 7871
rect 13369 7837 13403 7871
rect 4997 7769 5031 7803
rect 7297 7701 7331 7735
rect 11989 7701 12023 7735
rect 14933 7701 14967 7735
rect 7941 7497 7975 7531
rect 12449 7429 12483 7463
rect 9045 7361 9079 7395
rect 7665 7293 7699 7327
rect 7757 7293 7791 7327
rect 8585 7293 8619 7327
rect 8887 7293 8921 7327
rect 11989 7293 12023 7327
rect 12173 7293 12207 7327
rect 12265 7293 12299 7327
rect 12547 7293 12581 7327
rect 12725 7293 12759 7327
rect 8677 7225 8711 7259
rect 8769 7225 8803 7259
rect 9229 7225 9263 7259
rect 9597 7225 9631 7259
rect 12449 7225 12483 7259
rect 12633 7225 12667 7259
rect 8401 7157 8435 7191
rect 11345 7157 11379 7191
rect 6561 6953 6595 6987
rect 6729 6953 6763 6987
rect 8125 6953 8159 6987
rect 8677 6953 8711 6987
rect 10793 6953 10827 6987
rect 12357 6953 12391 6987
rect 6929 6885 6963 6919
rect 7573 6885 7607 6919
rect 11222 6885 11256 6919
rect 4629 6817 4663 6851
rect 4813 6817 4847 6851
rect 6009 6817 6043 6851
rect 6193 6817 6227 6851
rect 6285 6817 6319 6851
rect 6469 6817 6503 6851
rect 7205 6817 7239 6851
rect 7481 6817 7515 6851
rect 7665 6817 7699 6851
rect 7757 6817 7791 6851
rect 7941 6817 7975 6851
rect 8401 6817 8435 6851
rect 9790 6817 9824 6851
rect 10057 6817 10091 6851
rect 10333 6817 10367 6851
rect 10609 6817 10643 6851
rect 10977 6817 11011 6851
rect 12633 6817 12667 6851
rect 12725 6817 12759 6851
rect 13001 6817 13035 6851
rect 13093 6817 13127 6851
rect 13369 6817 13403 6851
rect 5825 6749 5859 6783
rect 7389 6749 7423 6783
rect 8217 6749 8251 6783
rect 10425 6749 10459 6783
rect 12449 6749 12483 6783
rect 13277 6749 13311 6783
rect 13645 6749 13679 6783
rect 6101 6681 6135 6715
rect 7021 6681 7055 6715
rect 4629 6613 4663 6647
rect 6745 6613 6779 6647
rect 8585 6613 8619 6647
rect 12541 6613 12575 6647
rect 13185 6613 13219 6647
rect 14933 6613 14967 6647
rect 6377 6409 6411 6443
rect 7389 6409 7423 6443
rect 9137 6409 9171 6443
rect 10609 6409 10643 6443
rect 12265 6409 12299 6443
rect 13553 6409 13587 6443
rect 5549 6341 5583 6375
rect 7205 6341 7239 6375
rect 12725 6341 12759 6375
rect 8769 6273 8803 6307
rect 4169 6205 4203 6239
rect 6285 6205 6319 6239
rect 7665 6205 7699 6239
rect 7849 6205 7883 6239
rect 8953 6205 8987 6239
rect 10885 6205 10919 6239
rect 12163 6205 12197 6239
rect 12357 6205 12391 6239
rect 12449 6205 12483 6239
rect 12541 6205 12575 6239
rect 12725 6205 12759 6239
rect 13553 6205 13587 6239
rect 13829 6205 13863 6239
rect 7343 6171 7377 6205
rect 4436 6137 4470 6171
rect 7573 6137 7607 6171
rect 8493 6137 8527 6171
rect 10609 6137 10643 6171
rect 7757 6069 7791 6103
rect 10793 6069 10827 6103
rect 13737 6069 13771 6103
rect 7573 5797 7607 5831
rect 10977 5797 11011 5831
rect 4528 5729 4562 5763
rect 7849 5729 7883 5763
rect 12725 5729 12759 5763
rect 12817 5729 12851 5763
rect 4261 5661 4295 5695
rect 13093 5661 13127 5695
rect 6285 5593 6319 5627
rect 5641 5525 5675 5559
rect 8033 5525 8067 5559
rect 14381 5525 14415 5559
rect 6009 5321 6043 5355
rect 13369 5253 13403 5287
rect 6929 5185 6963 5219
rect 7297 5185 7331 5219
rect 8677 5185 8711 5219
rect 10149 5185 10183 5219
rect 10517 5185 10551 5219
rect 10609 5185 10643 5219
rect 11989 5185 12023 5219
rect 12081 5185 12115 5219
rect 13001 5185 13035 5219
rect 5825 5117 5859 5151
rect 6009 5117 6043 5151
rect 6285 5117 6319 5151
rect 6377 5117 6411 5151
rect 7481 5117 7515 5151
rect 8401 5117 8435 5151
rect 8585 5117 8619 5151
rect 10333 5117 10367 5151
rect 10425 5117 10459 5151
rect 10793 5117 10827 5151
rect 10885 5117 10919 5151
rect 11805 5117 11839 5151
rect 11897 5117 11931 5151
rect 12265 5117 12299 5151
rect 12357 5117 12391 5151
rect 13093 5117 13127 5151
rect 13553 5117 13587 5151
rect 7849 5049 7883 5083
rect 8493 5049 8527 5083
rect 8922 5049 8956 5083
rect 13369 5049 13403 5083
rect 6193 4981 6227 5015
rect 7573 4981 7607 5015
rect 7665 4981 7699 5015
rect 10057 4981 10091 5015
rect 11529 4981 11563 5015
rect 11621 4981 11655 5015
rect 13185 4981 13219 5015
rect 13645 4981 13679 5015
rect 6193 4777 6227 4811
rect 7573 4777 7607 4811
rect 8217 4777 8251 4811
rect 10425 4777 10459 4811
rect 11253 4777 11287 4811
rect 11345 4777 11379 4811
rect 13369 4777 13403 4811
rect 5457 4709 5491 4743
rect 7849 4709 7883 4743
rect 10593 4709 10627 4743
rect 10793 4709 10827 4743
rect 11161 4709 11195 4743
rect 12234 4709 12268 4743
rect 5273 4641 5307 4675
rect 5549 4641 5583 4675
rect 6377 4641 6411 4675
rect 6653 4641 6687 4675
rect 6837 4641 6871 4675
rect 7205 4641 7239 4675
rect 7481 4641 7515 4675
rect 7757 4641 7791 4675
rect 7941 4641 7975 4675
rect 8401 4641 8435 4675
rect 10149 4641 10183 4675
rect 10333 4641 10367 4675
rect 11713 4641 11747 4675
rect 11989 4641 12023 4675
rect 6561 4573 6595 4607
rect 8125 4573 8159 4607
rect 8585 4573 8619 4607
rect 10977 4573 11011 4607
rect 6469 4505 6503 4539
rect 10333 4505 10367 4539
rect 11529 4505 11563 4539
rect 11805 4505 11839 4539
rect 5273 4437 5307 4471
rect 6929 4437 6963 4471
rect 7205 4437 7239 4471
rect 10609 4437 10643 4471
rect 6653 4233 6687 4267
rect 6929 4233 6963 4267
rect 11713 4233 11747 4267
rect 5641 4165 5675 4199
rect 8953 4165 8987 4199
rect 5917 4097 5951 4131
rect 7389 4097 7423 4131
rect 11069 4097 11103 4131
rect 4261 4029 4295 4063
rect 4528 4029 4562 4063
rect 6469 4029 6503 4063
rect 6561 4029 6595 4063
rect 6736 4029 6770 4063
rect 7113 4029 7147 4063
rect 7205 4029 7239 4063
rect 7297 4029 7331 4063
rect 9229 4029 9263 4063
rect 9321 4029 9355 4063
rect 9505 4029 9539 4063
rect 10977 4029 11011 4063
rect 11713 4029 11747 4063
rect 11897 4029 11931 4063
rect 8953 3961 8987 3995
rect 9137 3893 9171 3927
rect 9413 3893 9447 3927
rect 11345 3893 11379 3927
rect 8125 3689 8159 3723
rect 9597 3689 9631 3723
rect 9965 3689 9999 3723
rect 11161 3689 11195 3723
rect 7757 3621 7791 3655
rect 10057 3621 10091 3655
rect 7665 3553 7699 3587
rect 7857 3553 7891 3587
rect 8033 3553 8067 3587
rect 8217 3553 8251 3587
rect 8309 3553 8343 3587
rect 9045 3553 9079 3587
rect 9413 3553 9447 3587
rect 11102 3553 11136 3587
rect 11529 3553 11563 3587
rect 8861 3485 8895 3519
rect 11621 3485 11655 3519
rect 9137 3349 9171 3383
rect 10977 3349 11011 3383
rect 8401 3145 8435 3179
rect 11345 3145 11379 3179
rect 5457 3009 5491 3043
rect 7481 3009 7515 3043
rect 7665 3009 7699 3043
rect 7941 3009 7975 3043
rect 7054 2941 7088 2975
rect 7573 2941 7607 2975
rect 8033 2941 8067 2975
rect 9514 2941 9548 2975
rect 9781 2941 9815 2975
rect 9965 2941 9999 2975
rect 5724 2873 5758 2907
rect 10232 2873 10266 2907
rect 6837 2805 6871 2839
rect 6929 2805 6963 2839
rect 7113 2805 7147 2839
rect 5917 2601 5951 2635
rect 10333 2601 10367 2635
rect 5825 2465 5859 2499
rect 6009 2465 6043 2499
rect 10241 2465 10275 2499
rect 10425 2465 10459 2499
<< metal1 >>
rect 552 15258 15364 15280
rect 552 15206 2249 15258
rect 2301 15206 2313 15258
rect 2365 15206 2377 15258
rect 2429 15206 2441 15258
rect 2493 15206 2505 15258
rect 2557 15206 5951 15258
rect 6003 15206 6015 15258
rect 6067 15206 6079 15258
rect 6131 15206 6143 15258
rect 6195 15206 6207 15258
rect 6259 15206 9653 15258
rect 9705 15206 9717 15258
rect 9769 15206 9781 15258
rect 9833 15206 9845 15258
rect 9897 15206 9909 15258
rect 9961 15206 13355 15258
rect 13407 15206 13419 15258
rect 13471 15206 13483 15258
rect 13535 15206 13547 15258
rect 13599 15206 13611 15258
rect 13663 15206 15364 15258
rect 552 15184 15364 15206
rect 4890 15104 4896 15156
rect 4948 15104 4954 15156
rect 8849 15147 8907 15153
rect 8849 15113 8861 15147
rect 8895 15144 8907 15147
rect 10870 15144 10876 15156
rect 8895 15116 10876 15144
rect 8895 15113 8907 15116
rect 8849 15107 8907 15113
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 2501 15079 2559 15085
rect 2501 15045 2513 15079
rect 2547 15076 2559 15079
rect 5534 15076 5540 15088
rect 2547 15048 5540 15076
rect 2547 15045 2559 15048
rect 2501 15039 2559 15045
rect 5534 15036 5540 15048
rect 5592 15036 5598 15088
rect 1213 15011 1271 15017
rect 1213 14977 1225 15011
rect 1259 15008 1271 15011
rect 1259 14980 4752 15008
rect 1259 14977 1271 14980
rect 1213 14971 1271 14977
rect 842 14900 848 14952
rect 900 14940 906 14952
rect 1029 14943 1087 14949
rect 1029 14940 1041 14943
rect 900 14912 1041 14940
rect 900 14900 906 14912
rect 1029 14909 1041 14912
rect 1075 14909 1087 14943
rect 1029 14903 1087 14909
rect 2130 14900 2136 14952
rect 2188 14940 2194 14952
rect 2317 14943 2375 14949
rect 2317 14940 2329 14943
rect 2188 14912 2329 14940
rect 2188 14900 2194 14912
rect 2317 14909 2329 14912
rect 2363 14909 2375 14943
rect 2317 14903 2375 14909
rect 3418 14900 3424 14952
rect 3476 14940 3482 14952
rect 3513 14943 3571 14949
rect 3513 14940 3525 14943
rect 3476 14912 3525 14940
rect 3476 14900 3482 14912
rect 3513 14909 3525 14912
rect 3559 14909 3571 14943
rect 4724 14940 4752 14980
rect 4798 14968 4804 15020
rect 4856 15008 4862 15020
rect 4856 14980 5212 15008
rect 4856 14968 4862 14980
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4724 14912 4905 14940
rect 3513 14903 3571 14909
rect 4893 14909 4905 14912
rect 4939 14940 4951 14943
rect 5074 14940 5080 14952
rect 4939 14912 5080 14940
rect 4939 14909 4951 14912
rect 4893 14903 4951 14909
rect 5074 14900 5080 14912
rect 5132 14900 5138 14952
rect 5184 14949 5212 14980
rect 8570 14968 8576 15020
rect 8628 15008 8634 15020
rect 8628 14980 9076 15008
rect 8628 14968 8634 14980
rect 5169 14943 5227 14949
rect 5169 14909 5181 14943
rect 5215 14909 5227 14943
rect 5169 14903 5227 14909
rect 5261 14943 5319 14949
rect 5261 14909 5273 14943
rect 5307 14909 5319 14943
rect 5261 14903 5319 14909
rect 4706 14832 4712 14884
rect 4764 14872 4770 14884
rect 5276 14872 5304 14903
rect 5810 14900 5816 14952
rect 5868 14940 5874 14952
rect 6089 14943 6147 14949
rect 6089 14940 6101 14943
rect 5868 14912 6101 14940
rect 5868 14900 5874 14912
rect 6089 14909 6101 14912
rect 6135 14909 6147 14943
rect 6089 14903 6147 14909
rect 7282 14900 7288 14952
rect 7340 14940 7346 14952
rect 7377 14943 7435 14949
rect 7377 14940 7389 14943
rect 7340 14912 7389 14940
rect 7340 14900 7346 14912
rect 7377 14909 7389 14912
rect 7423 14909 7435 14943
rect 7377 14903 7435 14909
rect 7558 14900 7564 14952
rect 7616 14940 7622 14952
rect 8665 14943 8723 14949
rect 8665 14940 8677 14943
rect 7616 14912 8677 14940
rect 7616 14900 7622 14912
rect 8665 14909 8677 14912
rect 8711 14909 8723 14943
rect 8665 14903 8723 14909
rect 8938 14900 8944 14952
rect 8996 14900 9002 14952
rect 9048 14949 9076 14980
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14909 9091 14943
rect 9033 14903 9091 14909
rect 9953 14943 10011 14949
rect 9953 14909 9965 14943
rect 9999 14940 10011 14943
rect 10042 14940 10048 14952
rect 9999 14912 10048 14940
rect 9999 14909 10011 14912
rect 9953 14903 10011 14909
rect 10042 14900 10048 14912
rect 10100 14900 10106 14952
rect 11146 14900 11152 14952
rect 11204 14940 11210 14952
rect 11241 14943 11299 14949
rect 11241 14940 11253 14943
rect 11204 14912 11253 14940
rect 11204 14900 11210 14912
rect 11241 14909 11253 14912
rect 11287 14909 11299 14943
rect 11241 14903 11299 14909
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 12713 14943 12771 14949
rect 12713 14940 12725 14943
rect 12492 14912 12725 14940
rect 12492 14900 12498 14912
rect 12713 14909 12725 14912
rect 12759 14909 12771 14943
rect 12713 14903 12771 14909
rect 13722 14900 13728 14952
rect 13780 14940 13786 14952
rect 13817 14943 13875 14949
rect 13817 14940 13829 14943
rect 13780 14912 13829 14940
rect 13780 14900 13786 14912
rect 13817 14909 13829 14912
rect 13863 14909 13875 14943
rect 13817 14903 13875 14909
rect 4764 14844 5304 14872
rect 4764 14832 4770 14844
rect 10502 14832 10508 14884
rect 10560 14872 10566 14884
rect 10560 14844 12572 14872
rect 10560 14832 10566 14844
rect 3697 14807 3755 14813
rect 3697 14773 3709 14807
rect 3743 14804 3755 14807
rect 4430 14804 4436 14816
rect 3743 14776 4436 14804
rect 3743 14773 3755 14776
rect 3697 14767 3755 14773
rect 4430 14764 4436 14776
rect 4488 14764 4494 14816
rect 4614 14764 4620 14816
rect 4672 14764 4678 14816
rect 5442 14764 5448 14816
rect 5500 14764 5506 14816
rect 6270 14764 6276 14816
rect 6328 14764 6334 14816
rect 7561 14807 7619 14813
rect 7561 14773 7573 14807
rect 7607 14804 7619 14807
rect 7650 14804 7656 14816
rect 7607 14776 7656 14804
rect 7607 14773 7619 14776
rect 7561 14767 7619 14773
rect 7650 14764 7656 14776
rect 7708 14764 7714 14816
rect 8386 14764 8392 14816
rect 8444 14764 8450 14816
rect 9030 14764 9036 14816
rect 9088 14804 9094 14816
rect 9217 14807 9275 14813
rect 9217 14804 9229 14807
rect 9088 14776 9229 14804
rect 9088 14764 9094 14776
rect 9217 14773 9229 14776
rect 9263 14773 9275 14807
rect 9217 14767 9275 14773
rect 10137 14807 10195 14813
rect 10137 14773 10149 14807
rect 10183 14804 10195 14807
rect 10778 14804 10784 14816
rect 10183 14776 10784 14804
rect 10183 14773 10195 14776
rect 10137 14767 10195 14773
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 11330 14764 11336 14816
rect 11388 14804 11394 14816
rect 12544 14813 12572 14844
rect 11425 14807 11483 14813
rect 11425 14804 11437 14807
rect 11388 14776 11437 14804
rect 11388 14764 11394 14776
rect 11425 14773 11437 14776
rect 11471 14773 11483 14807
rect 11425 14767 11483 14773
rect 12529 14807 12587 14813
rect 12529 14773 12541 14807
rect 12575 14773 12587 14807
rect 12529 14767 12587 14773
rect 12802 14764 12808 14816
rect 12860 14764 12866 14816
rect 13998 14764 14004 14816
rect 14056 14764 14062 14816
rect 552 14714 15520 14736
rect 552 14662 4100 14714
rect 4152 14662 4164 14714
rect 4216 14662 4228 14714
rect 4280 14662 4292 14714
rect 4344 14662 4356 14714
rect 4408 14662 7802 14714
rect 7854 14662 7866 14714
rect 7918 14662 7930 14714
rect 7982 14662 7994 14714
rect 8046 14662 8058 14714
rect 8110 14662 11504 14714
rect 11556 14662 11568 14714
rect 11620 14662 11632 14714
rect 11684 14662 11696 14714
rect 11748 14662 11760 14714
rect 11812 14662 15206 14714
rect 15258 14662 15270 14714
rect 15322 14662 15334 14714
rect 15386 14662 15398 14714
rect 15450 14662 15462 14714
rect 15514 14662 15520 14714
rect 552 14640 15520 14662
rect 5813 14603 5871 14609
rect 5813 14569 5825 14603
rect 5859 14600 5871 14603
rect 7466 14600 7472 14612
rect 5859 14572 7472 14600
rect 5859 14569 5871 14572
rect 5813 14563 5871 14569
rect 7466 14560 7472 14572
rect 7524 14600 7530 14612
rect 8113 14603 8171 14609
rect 7524 14572 7880 14600
rect 7524 14560 7530 14572
rect 5258 14532 5264 14544
rect 5092 14504 5264 14532
rect 4821 14467 4879 14473
rect 4821 14433 4833 14467
rect 4867 14464 4879 14467
rect 4982 14464 4988 14476
rect 4867 14436 4988 14464
rect 4867 14433 4879 14436
rect 4821 14427 4879 14433
rect 4982 14424 4988 14436
rect 5040 14424 5046 14476
rect 5092 14473 5120 14504
rect 5258 14492 5264 14504
rect 5316 14532 5322 14544
rect 5316 14504 7788 14532
rect 5316 14492 5322 14504
rect 5077 14467 5135 14473
rect 5077 14433 5089 14467
rect 5123 14433 5135 14467
rect 5077 14427 5135 14433
rect 5166 14424 5172 14476
rect 5224 14464 5230 14476
rect 5445 14467 5503 14473
rect 5445 14464 5457 14467
rect 5224 14436 5457 14464
rect 5224 14424 5230 14436
rect 5445 14433 5457 14436
rect 5491 14433 5503 14467
rect 5445 14427 5503 14433
rect 3697 14263 3755 14269
rect 3697 14229 3709 14263
rect 3743 14260 3755 14263
rect 4798 14260 4804 14272
rect 3743 14232 4804 14260
rect 3743 14229 3755 14232
rect 3697 14223 3755 14229
rect 4798 14220 4804 14232
rect 4856 14220 4862 14272
rect 5166 14220 5172 14272
rect 5224 14260 5230 14272
rect 5261 14263 5319 14269
rect 5261 14260 5273 14263
rect 5224 14232 5273 14260
rect 5224 14220 5230 14232
rect 5261 14229 5273 14232
rect 5307 14229 5319 14263
rect 5261 14223 5319 14229
rect 5350 14220 5356 14272
rect 5408 14260 5414 14272
rect 5460 14260 5488 14427
rect 6914 14424 6920 14476
rect 6972 14473 6978 14476
rect 7208 14473 7236 14504
rect 6972 14427 6984 14473
rect 7193 14467 7251 14473
rect 7193 14433 7205 14467
rect 7239 14433 7251 14467
rect 7193 14427 7251 14433
rect 6972 14424 6978 14427
rect 7558 14424 7564 14476
rect 7616 14424 7622 14476
rect 7576 14328 7604 14424
rect 7760 14396 7788 14504
rect 7852 14473 7880 14572
rect 8113 14569 8125 14603
rect 8159 14600 8171 14603
rect 8202 14600 8208 14612
rect 8159 14572 8208 14600
rect 8159 14569 8171 14572
rect 8113 14563 8171 14569
rect 8202 14560 8208 14572
rect 8260 14600 8266 14612
rect 8938 14600 8944 14612
rect 8260 14572 8944 14600
rect 8260 14560 8266 14572
rect 8938 14560 8944 14572
rect 8996 14560 9002 14612
rect 13998 14560 14004 14612
rect 14056 14560 14062 14612
rect 12713 14535 12771 14541
rect 9508 14504 12388 14532
rect 7837 14467 7895 14473
rect 7837 14433 7849 14467
rect 7883 14433 7895 14467
rect 7837 14427 7895 14433
rect 9214 14424 9220 14476
rect 9272 14473 9278 14476
rect 9272 14427 9284 14473
rect 9272 14424 9278 14427
rect 9508 14408 9536 14504
rect 12360 14473 12388 14504
rect 12713 14501 12725 14535
rect 12759 14532 12771 14535
rect 12802 14532 12808 14544
rect 12759 14504 12808 14532
rect 12759 14501 12771 14504
rect 12713 14495 12771 14501
rect 12802 14492 12808 14504
rect 12860 14492 12866 14544
rect 10781 14467 10839 14473
rect 10781 14433 10793 14467
rect 10827 14464 10839 14467
rect 12078 14467 12136 14473
rect 12078 14464 12090 14467
rect 10827 14436 12090 14464
rect 10827 14433 10839 14436
rect 10781 14427 10839 14433
rect 12078 14433 12090 14436
rect 12124 14433 12136 14467
rect 12078 14427 12136 14433
rect 12345 14467 12403 14473
rect 12345 14433 12357 14467
rect 12391 14464 12403 14467
rect 12434 14464 12440 14476
rect 12391 14436 12440 14464
rect 12391 14433 12403 14436
rect 12345 14427 12403 14433
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 14016 14464 14044 14560
rect 14369 14467 14427 14473
rect 14369 14464 14381 14467
rect 8478 14396 8484 14408
rect 7760 14368 8484 14396
rect 8478 14356 8484 14368
rect 8536 14356 8542 14408
rect 9490 14356 9496 14408
rect 9548 14356 9554 14408
rect 10134 14356 10140 14408
rect 10192 14356 10198 14408
rect 10226 14356 10232 14408
rect 10284 14396 10290 14408
rect 10505 14399 10563 14405
rect 10505 14396 10517 14399
rect 10284 14368 10517 14396
rect 10284 14356 10290 14368
rect 10505 14365 10517 14368
rect 10551 14365 10563 14399
rect 10505 14359 10563 14365
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14396 10655 14399
rect 11330 14396 11336 14408
rect 10643 14368 11336 14396
rect 10643 14365 10655 14368
rect 10597 14359 10655 14365
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 13832 14396 13860 14450
rect 14016 14436 14381 14464
rect 14369 14433 14381 14436
rect 14415 14433 14427 14467
rect 14369 14427 14427 14433
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 13832 14368 14473 14396
rect 14461 14365 14473 14368
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 7208 14300 7604 14328
rect 7208 14260 7236 14300
rect 5408 14232 7236 14260
rect 5408 14220 5414 14232
rect 7282 14220 7288 14272
rect 7340 14220 7346 14272
rect 7374 14220 7380 14272
rect 7432 14260 7438 14272
rect 7469 14263 7527 14269
rect 7469 14260 7481 14263
rect 7432 14232 7481 14260
rect 7432 14220 7438 14232
rect 7469 14229 7481 14232
rect 7515 14229 7527 14263
rect 7469 14223 7527 14229
rect 9122 14220 9128 14272
rect 9180 14260 9186 14272
rect 10962 14260 10968 14272
rect 9180 14232 10968 14260
rect 9180 14220 9186 14232
rect 10962 14220 10968 14232
rect 11020 14220 11026 14272
rect 14182 14220 14188 14272
rect 14240 14220 14246 14272
rect 552 14170 15364 14192
rect 552 14118 2249 14170
rect 2301 14118 2313 14170
rect 2365 14118 2377 14170
rect 2429 14118 2441 14170
rect 2493 14118 2505 14170
rect 2557 14118 5951 14170
rect 6003 14118 6015 14170
rect 6067 14118 6079 14170
rect 6131 14118 6143 14170
rect 6195 14118 6207 14170
rect 6259 14118 9653 14170
rect 9705 14118 9717 14170
rect 9769 14118 9781 14170
rect 9833 14118 9845 14170
rect 9897 14118 9909 14170
rect 9961 14118 13355 14170
rect 13407 14118 13419 14170
rect 13471 14118 13483 14170
rect 13535 14118 13547 14170
rect 13599 14118 13611 14170
rect 13663 14118 15364 14170
rect 552 14096 15364 14118
rect 4890 14016 4896 14068
rect 4948 14016 4954 14068
rect 4982 14016 4988 14068
rect 5040 14016 5046 14068
rect 6914 14016 6920 14068
rect 6972 14056 6978 14068
rect 7009 14059 7067 14065
rect 7009 14056 7021 14059
rect 6972 14028 7021 14056
rect 6972 14016 6978 14028
rect 7009 14025 7021 14028
rect 7055 14025 7067 14059
rect 7009 14019 7067 14025
rect 9214 14016 9220 14068
rect 9272 14016 9278 14068
rect 10134 14016 10140 14068
rect 10192 14056 10198 14068
rect 10413 14059 10471 14065
rect 10413 14056 10425 14059
rect 10192 14028 10425 14056
rect 10192 14016 10198 14028
rect 10413 14025 10425 14028
rect 10459 14025 10471 14059
rect 10413 14019 10471 14025
rect 10870 14016 10876 14068
rect 10928 14056 10934 14068
rect 11054 14056 11060 14068
rect 10928 14028 11060 14056
rect 10928 14016 10934 14028
rect 11054 14016 11060 14028
rect 11112 14056 11118 14068
rect 11241 14059 11299 14065
rect 11241 14056 11253 14059
rect 11112 14028 11253 14056
rect 11112 14016 11118 14028
rect 11241 14025 11253 14028
rect 11287 14025 11299 14059
rect 11241 14019 11299 14025
rect 12066 14016 12072 14068
rect 12124 14056 12130 14068
rect 13906 14056 13912 14068
rect 12124 14028 13912 14056
rect 12124 14016 12130 14028
rect 13906 14016 13912 14028
rect 13964 14016 13970 14068
rect 4908 13988 4936 14016
rect 6178 13988 6184 14000
rect 4908 13960 6184 13988
rect 6178 13948 6184 13960
rect 6236 13948 6242 14000
rect 8754 13988 8760 14000
rect 6288 13960 8760 13988
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 4614 13920 4620 13932
rect 4387 13892 4620 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 4614 13880 4620 13892
rect 4672 13880 4678 13932
rect 5166 13920 5172 13932
rect 4724 13892 5172 13920
rect 4522 13812 4528 13864
rect 4580 13852 4586 13864
rect 4724 13861 4752 13892
rect 5166 13880 5172 13892
rect 5224 13920 5230 13932
rect 5224 13892 5534 13920
rect 5224 13880 5230 13892
rect 4709 13855 4767 13861
rect 4709 13852 4721 13855
rect 4580 13824 4721 13852
rect 4580 13812 4586 13824
rect 4709 13821 4721 13824
rect 4755 13821 4767 13855
rect 4709 13815 4767 13821
rect 4801 13855 4859 13861
rect 4801 13821 4813 13855
rect 4847 13821 4859 13855
rect 5506 13852 5534 13892
rect 6288 13852 6316 13960
rect 8754 13948 8760 13960
rect 8812 13988 8818 14000
rect 10778 13988 10784 14000
rect 8812 13960 8984 13988
rect 8812 13948 8818 13960
rect 6365 13923 6423 13929
rect 6365 13889 6377 13923
rect 6411 13920 6423 13923
rect 7282 13920 7288 13932
rect 6411 13892 7288 13920
rect 6411 13889 6423 13892
rect 6365 13883 6423 13889
rect 7282 13880 7288 13892
rect 7340 13880 7346 13932
rect 8386 13880 8392 13932
rect 8444 13920 8450 13932
rect 8573 13923 8631 13929
rect 8573 13920 8585 13923
rect 8444 13892 8585 13920
rect 8444 13880 8450 13892
rect 8573 13889 8585 13892
rect 8619 13889 8631 13923
rect 8573 13883 8631 13889
rect 6733 13855 6791 13861
rect 6733 13852 6745 13855
rect 5506 13824 6745 13852
rect 4801 13815 4859 13821
rect 6733 13821 6745 13824
rect 6779 13821 6791 13855
rect 6733 13815 6791 13821
rect 6825 13855 6883 13861
rect 6825 13821 6837 13855
rect 6871 13852 6883 13855
rect 7650 13852 7656 13864
rect 6871 13824 7656 13852
rect 6871 13821 6883 13824
rect 6825 13815 6883 13821
rect 4816 13784 4844 13815
rect 7650 13812 7656 13824
rect 7708 13852 7714 13864
rect 8846 13852 8852 13864
rect 7708 13824 8852 13852
rect 7708 13812 7714 13824
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 8956 13861 8984 13960
rect 9048 13960 10784 13988
rect 9048 13861 9076 13960
rect 10778 13948 10784 13960
rect 10836 13948 10842 14000
rect 12894 13948 12900 14000
rect 12952 13948 12958 14000
rect 14182 13920 14188 13932
rect 11532 13892 14188 13920
rect 8941 13855 8999 13861
rect 8941 13821 8953 13855
rect 8987 13821 8999 13855
rect 8941 13815 8999 13821
rect 9033 13855 9091 13861
rect 9033 13821 9045 13855
rect 9079 13821 9091 13855
rect 9033 13815 9091 13821
rect 10226 13812 10232 13864
rect 10284 13852 10290 13864
rect 10962 13861 10968 13864
rect 10597 13855 10655 13861
rect 10597 13852 10609 13855
rect 10284 13824 10609 13852
rect 10284 13812 10290 13824
rect 10597 13821 10609 13824
rect 10643 13821 10655 13855
rect 10959 13852 10968 13861
rect 10923 13824 10968 13852
rect 10597 13815 10655 13821
rect 10959 13815 10968 13824
rect 10962 13812 10968 13815
rect 11020 13812 11026 13864
rect 5442 13784 5448 13796
rect 4816 13756 5448 13784
rect 5442 13744 5448 13756
rect 5500 13784 5506 13796
rect 11422 13784 11428 13796
rect 5500 13756 11428 13784
rect 5500 13744 5506 13756
rect 11422 13744 11428 13756
rect 11480 13744 11486 13796
rect 11532 13793 11560 13892
rect 14182 13880 14188 13892
rect 14240 13920 14246 13932
rect 14240 13892 14596 13920
rect 14240 13880 14246 13892
rect 11882 13812 11888 13864
rect 11940 13812 11946 13864
rect 12066 13812 12072 13864
rect 12124 13812 12130 13864
rect 12158 13812 12164 13864
rect 12216 13812 12222 13864
rect 12342 13812 12348 13864
rect 12400 13812 12406 13864
rect 12618 13812 12624 13864
rect 12676 13812 12682 13864
rect 14458 13812 14464 13864
rect 14516 13812 14522 13864
rect 14568 13861 14596 13892
rect 14553 13855 14611 13861
rect 14553 13821 14565 13855
rect 14599 13821 14611 13855
rect 14553 13815 14611 13821
rect 15102 13812 15108 13864
rect 15160 13812 15166 13864
rect 11517 13787 11575 13793
rect 11517 13753 11529 13787
rect 11563 13753 11575 13787
rect 11517 13747 11575 13753
rect 11977 13787 12035 13793
rect 11977 13753 11989 13787
rect 12023 13784 12035 13787
rect 12713 13787 12771 13793
rect 12713 13784 12725 13787
rect 12023 13756 12725 13784
rect 12023 13753 12035 13756
rect 11977 13747 12035 13753
rect 12713 13753 12725 13756
rect 12759 13753 12771 13787
rect 12713 13747 12771 13753
rect 12897 13787 12955 13793
rect 12897 13753 12909 13787
rect 12943 13784 12955 13787
rect 12986 13784 12992 13796
rect 12943 13756 12992 13784
rect 12943 13753 12955 13756
rect 12897 13747 12955 13753
rect 6178 13676 6184 13728
rect 6236 13716 6242 13728
rect 7374 13716 7380 13728
rect 6236 13688 7380 13716
rect 6236 13676 6242 13688
rect 7374 13676 7380 13688
rect 7432 13716 7438 13728
rect 7650 13716 7656 13728
rect 7432 13688 7656 13716
rect 7432 13676 7438 13688
rect 7650 13676 7656 13688
rect 7708 13716 7714 13728
rect 11532 13716 11560 13747
rect 12986 13744 12992 13756
rect 13044 13744 13050 13796
rect 14476 13784 14504 13812
rect 15120 13784 15148 13812
rect 14476 13756 15148 13784
rect 7708 13688 11560 13716
rect 7708 13676 7714 13688
rect 12250 13676 12256 13728
rect 12308 13676 12314 13728
rect 12802 13676 12808 13728
rect 12860 13716 12866 13728
rect 13817 13719 13875 13725
rect 13817 13716 13829 13719
rect 12860 13688 13829 13716
rect 12860 13676 12866 13688
rect 13817 13685 13829 13688
rect 13863 13685 13875 13719
rect 13817 13679 13875 13685
rect 14642 13676 14648 13728
rect 14700 13676 14706 13728
rect 552 13626 15520 13648
rect 552 13574 4100 13626
rect 4152 13574 4164 13626
rect 4216 13574 4228 13626
rect 4280 13574 4292 13626
rect 4344 13574 4356 13626
rect 4408 13574 7802 13626
rect 7854 13574 7866 13626
rect 7918 13574 7930 13626
rect 7982 13574 7994 13626
rect 8046 13574 8058 13626
rect 8110 13574 11504 13626
rect 11556 13574 11568 13626
rect 11620 13574 11632 13626
rect 11684 13574 11696 13626
rect 11748 13574 11760 13626
rect 11812 13574 15206 13626
rect 15258 13574 15270 13626
rect 15322 13574 15334 13626
rect 15386 13574 15398 13626
rect 15450 13574 15462 13626
rect 15514 13574 15520 13626
rect 552 13552 15520 13574
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 12161 13515 12219 13521
rect 12161 13512 12173 13515
rect 11940 13484 12173 13512
rect 11940 13472 11946 13484
rect 12161 13481 12173 13484
rect 12207 13481 12219 13515
rect 12161 13475 12219 13481
rect 12250 13472 12256 13524
rect 12308 13472 12314 13524
rect 12434 13472 12440 13524
rect 12492 13472 12498 13524
rect 12618 13472 12624 13524
rect 12676 13512 12682 13524
rect 12713 13515 12771 13521
rect 12713 13512 12725 13515
rect 12676 13484 12725 13512
rect 12676 13472 12682 13484
rect 12713 13481 12725 13484
rect 12759 13481 12771 13515
rect 12713 13475 12771 13481
rect 14921 13515 14979 13521
rect 14921 13481 14933 13515
rect 14967 13512 14979 13515
rect 15102 13512 15108 13524
rect 14967 13484 15108 13512
rect 14967 13481 14979 13484
rect 14921 13475 14979 13481
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 12066 13444 12072 13456
rect 8220 13416 12072 13444
rect 4341 13379 4399 13385
rect 4341 13345 4353 13379
rect 4387 13376 4399 13379
rect 4522 13376 4528 13388
rect 4387 13348 4528 13376
rect 4387 13345 4399 13348
rect 4341 13339 4399 13345
rect 4522 13336 4528 13348
rect 4580 13336 4586 13388
rect 6089 13379 6147 13385
rect 6089 13376 6101 13379
rect 5506 13348 6101 13376
rect 3881 13311 3939 13317
rect 3881 13277 3893 13311
rect 3927 13308 3939 13311
rect 4154 13308 4160 13320
rect 3927 13280 4160 13308
rect 3927 13277 3939 13280
rect 3881 13271 3939 13277
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13277 4307 13311
rect 4540 13308 4568 13336
rect 5506 13308 5534 13348
rect 6089 13345 6101 13348
rect 6135 13345 6147 13379
rect 8220 13376 8248 13416
rect 12066 13404 12072 13416
rect 12124 13404 12130 13456
rect 6089 13339 6147 13345
rect 6380 13348 8248 13376
rect 8317 13379 8375 13385
rect 4540 13280 5534 13308
rect 5997 13311 6055 13317
rect 4249 13271 4307 13277
rect 5997 13277 6009 13311
rect 6043 13300 6055 13311
rect 6270 13308 6276 13320
rect 6196 13300 6276 13308
rect 6043 13280 6276 13300
rect 6043 13277 6224 13280
rect 5997 13272 6224 13277
rect 5997 13271 6055 13272
rect 4264 13240 4292 13271
rect 6270 13268 6276 13280
rect 6328 13308 6334 13320
rect 6380 13308 6408 13348
rect 8317 13345 8329 13379
rect 8363 13376 8375 13379
rect 8662 13376 8668 13388
rect 8363 13348 8668 13376
rect 8363 13345 8375 13348
rect 8317 13339 8375 13345
rect 8662 13336 8668 13348
rect 8720 13336 8726 13388
rect 9306 13385 9312 13388
rect 9300 13339 9312 13385
rect 9306 13336 9312 13339
rect 9364 13336 9370 13388
rect 11655 13379 11713 13385
rect 11655 13376 11667 13379
rect 10060 13348 11667 13376
rect 6328 13280 6408 13308
rect 6328 13268 6334 13280
rect 6454 13268 6460 13320
rect 6512 13268 6518 13320
rect 8570 13268 8576 13320
rect 8628 13308 8634 13320
rect 9033 13311 9091 13317
rect 9033 13308 9045 13311
rect 8628 13280 9045 13308
rect 8628 13268 8634 13280
rect 9033 13277 9045 13280
rect 9079 13277 9091 13311
rect 9033 13271 9091 13277
rect 4338 13240 4344 13252
rect 4264 13212 4344 13240
rect 4338 13200 4344 13212
rect 4396 13240 4402 13252
rect 4396 13212 7696 13240
rect 4396 13200 4402 13212
rect 4522 13132 4528 13184
rect 4580 13132 4586 13184
rect 5810 13132 5816 13184
rect 5868 13132 5874 13184
rect 7193 13175 7251 13181
rect 7193 13141 7205 13175
rect 7239 13172 7251 13175
rect 7374 13172 7380 13184
rect 7239 13144 7380 13172
rect 7239 13141 7251 13144
rect 7193 13135 7251 13141
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 7668 13172 7696 13212
rect 10060 13172 10088 13348
rect 11655 13345 11667 13348
rect 11701 13345 11713 13379
rect 11655 13339 11713 13345
rect 11790 13336 11796 13388
rect 11848 13336 11854 13388
rect 11882 13336 11888 13388
rect 11940 13336 11946 13388
rect 11977 13379 12035 13385
rect 11977 13345 11989 13379
rect 12023 13376 12035 13379
rect 12268 13376 12296 13472
rect 12452 13444 12480 13472
rect 13262 13444 13268 13456
rect 12452 13416 13268 13444
rect 13262 13404 13268 13416
rect 13320 13444 13326 13456
rect 13320 13416 13400 13444
rect 13320 13404 13326 13416
rect 12023 13348 12296 13376
rect 12023 13345 12035 13348
rect 11977 13339 12035 13345
rect 12342 13336 12348 13388
rect 12400 13376 12406 13388
rect 12437 13379 12495 13385
rect 12437 13376 12449 13379
rect 12400 13348 12449 13376
rect 12400 13336 12406 13348
rect 12437 13345 12449 13348
rect 12483 13345 12495 13379
rect 12437 13339 12495 13345
rect 12802 13336 12808 13388
rect 12860 13336 12866 13388
rect 12894 13336 12900 13388
rect 12952 13336 12958 13388
rect 13372 13385 13400 13416
rect 13357 13379 13415 13385
rect 13357 13345 13369 13379
rect 13403 13345 13415 13379
rect 13357 13339 13415 13345
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 11296 13280 11529 13308
rect 11296 13268 11302 13280
rect 11517 13277 11529 13280
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 12713 13311 12771 13317
rect 12713 13277 12725 13311
rect 12759 13308 12771 13311
rect 12820 13308 12848 13336
rect 12759 13280 12848 13308
rect 12912 13308 12940 13336
rect 13633 13311 13691 13317
rect 13633 13308 13645 13311
rect 12912 13280 13645 13308
rect 12759 13277 12771 13280
rect 12713 13271 12771 13277
rect 13633 13277 13645 13280
rect 13679 13277 13691 13311
rect 13633 13271 13691 13277
rect 7668 13144 10088 13172
rect 10410 13132 10416 13184
rect 10468 13132 10474 13184
rect 12526 13132 12532 13184
rect 12584 13132 12590 13184
rect 552 13082 15364 13104
rect 552 13030 2249 13082
rect 2301 13030 2313 13082
rect 2365 13030 2377 13082
rect 2429 13030 2441 13082
rect 2493 13030 2505 13082
rect 2557 13030 5951 13082
rect 6003 13030 6015 13082
rect 6067 13030 6079 13082
rect 6131 13030 6143 13082
rect 6195 13030 6207 13082
rect 6259 13030 9653 13082
rect 9705 13030 9717 13082
rect 9769 13030 9781 13082
rect 9833 13030 9845 13082
rect 9897 13030 9909 13082
rect 9961 13030 13355 13082
rect 13407 13030 13419 13082
rect 13471 13030 13483 13082
rect 13535 13030 13547 13082
rect 13599 13030 13611 13082
rect 13663 13030 15364 13082
rect 552 13008 15364 13030
rect 6454 12928 6460 12980
rect 6512 12968 6518 12980
rect 6733 12971 6791 12977
rect 6733 12968 6745 12971
rect 6512 12940 6745 12968
rect 6512 12928 6518 12940
rect 6733 12937 6745 12940
rect 6779 12937 6791 12971
rect 6733 12931 6791 12937
rect 7101 12971 7159 12977
rect 7101 12937 7113 12971
rect 7147 12968 7159 12971
rect 7282 12968 7288 12980
rect 7147 12940 7288 12968
rect 7147 12937 7159 12940
rect 7101 12931 7159 12937
rect 7282 12928 7288 12940
rect 7340 12928 7346 12980
rect 7558 12928 7564 12980
rect 7616 12928 7622 12980
rect 7650 12928 7656 12980
rect 7708 12968 7714 12980
rect 7745 12971 7803 12977
rect 7745 12968 7757 12971
rect 7708 12940 7757 12968
rect 7708 12928 7714 12940
rect 7745 12937 7757 12940
rect 7791 12937 7803 12971
rect 7745 12931 7803 12937
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 9033 12971 9091 12977
rect 9033 12968 9045 12971
rect 8720 12940 9045 12968
rect 8720 12928 8726 12940
rect 9033 12937 9045 12940
rect 9079 12937 9091 12971
rect 9033 12931 9091 12937
rect 9306 12928 9312 12980
rect 9364 12968 9370 12980
rect 9953 12971 10011 12977
rect 9953 12968 9965 12971
rect 9364 12940 9965 12968
rect 9364 12928 9370 12940
rect 9953 12937 9965 12940
rect 9999 12937 10011 12971
rect 9953 12931 10011 12937
rect 10686 12928 10692 12980
rect 10744 12968 10750 12980
rect 10873 12971 10931 12977
rect 10873 12968 10885 12971
rect 10744 12940 10885 12968
rect 10744 12928 10750 12940
rect 10873 12937 10885 12940
rect 10919 12968 10931 12971
rect 11054 12968 11060 12980
rect 10919 12940 11060 12968
rect 10919 12937 10931 12940
rect 10873 12931 10931 12937
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 11790 12928 11796 12980
rect 11848 12968 11854 12980
rect 11848 12940 12940 12968
rect 11848 12928 11854 12940
rect 7576 12900 7604 12928
rect 10704 12900 10732 12928
rect 7024 12872 7972 12900
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 5258 12832 5264 12844
rect 4663 12804 5264 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 7024 12841 7052 12872
rect 7009 12835 7067 12841
rect 7009 12801 7021 12835
rect 7055 12801 7067 12835
rect 7009 12795 7067 12801
rect 7116 12804 7328 12832
rect 4361 12767 4419 12773
rect 4361 12733 4373 12767
rect 4407 12764 4419 12767
rect 4522 12764 4528 12776
rect 4407 12736 4528 12764
rect 4407 12733 4419 12736
rect 4361 12727 4419 12733
rect 4522 12724 4528 12736
rect 4580 12724 4586 12776
rect 5528 12767 5586 12773
rect 5528 12733 5540 12767
rect 5574 12764 5586 12767
rect 5810 12764 5816 12776
rect 5574 12736 5816 12764
rect 5574 12733 5586 12736
rect 5528 12727 5586 12733
rect 5810 12724 5816 12736
rect 5868 12724 5874 12776
rect 7116 12773 7144 12804
rect 7095 12767 7153 12773
rect 7095 12733 7107 12767
rect 7141 12733 7153 12767
rect 7095 12727 7153 12733
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12733 7251 12767
rect 7300 12764 7328 12804
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 7944 12841 7972 12872
rect 8680 12872 10732 12900
rect 7929 12835 7987 12841
rect 7432 12804 7696 12832
rect 7432 12792 7438 12804
rect 7668 12773 7696 12804
rect 7929 12801 7941 12835
rect 7975 12801 7987 12835
rect 7929 12795 7987 12801
rect 7653 12767 7711 12773
rect 7300 12736 7604 12764
rect 7193 12727 7251 12733
rect 7208 12696 7236 12727
rect 6932 12668 7236 12696
rect 7576 12696 7604 12736
rect 7653 12733 7665 12767
rect 7699 12733 7711 12767
rect 7653 12727 7711 12733
rect 8680 12696 8708 12872
rect 8754 12792 8760 12844
rect 8812 12832 8818 12844
rect 10226 12832 10232 12844
rect 8812 12804 10232 12832
rect 8812 12792 8818 12804
rect 10226 12792 10232 12804
rect 10284 12792 10290 12844
rect 10428 12804 11054 12832
rect 8849 12767 8907 12773
rect 8849 12733 8861 12767
rect 8895 12764 8907 12767
rect 9030 12764 9036 12776
rect 8895 12736 9036 12764
rect 8895 12733 8907 12736
rect 8849 12727 8907 12733
rect 9030 12724 9036 12736
rect 9088 12724 9094 12776
rect 10137 12767 10195 12773
rect 10137 12733 10149 12767
rect 10183 12733 10195 12767
rect 10137 12727 10195 12733
rect 7576 12668 8708 12696
rect 6932 12640 6960 12668
rect 3234 12588 3240 12640
rect 3292 12588 3298 12640
rect 6641 12631 6699 12637
rect 6641 12597 6653 12631
rect 6687 12628 6699 12631
rect 6914 12628 6920 12640
rect 6687 12600 6920 12628
rect 6687 12597 6699 12600
rect 6641 12591 6699 12597
rect 6914 12588 6920 12600
rect 6972 12588 6978 12640
rect 7282 12588 7288 12640
rect 7340 12588 7346 12640
rect 8205 12631 8263 12637
rect 8205 12597 8217 12631
rect 8251 12628 8263 12631
rect 8389 12631 8447 12637
rect 8389 12628 8401 12631
rect 8251 12600 8401 12628
rect 8251 12597 8263 12600
rect 8205 12591 8263 12597
rect 8389 12597 8401 12600
rect 8435 12597 8447 12631
rect 10152 12628 10180 12727
rect 10244 12696 10272 12792
rect 10428 12776 10456 12804
rect 10410 12724 10416 12776
rect 10468 12724 10474 12776
rect 10873 12767 10931 12773
rect 10873 12733 10885 12767
rect 10919 12733 10931 12767
rect 11026 12764 11054 12804
rect 11241 12767 11299 12773
rect 11241 12764 11253 12767
rect 11026 12736 11253 12764
rect 10873 12727 10931 12733
rect 11241 12733 11253 12736
rect 11287 12733 11299 12767
rect 11241 12727 11299 12733
rect 11333 12767 11391 12773
rect 11333 12733 11345 12767
rect 11379 12733 11391 12767
rect 11333 12727 11391 12733
rect 10888 12696 10916 12727
rect 10244 12668 10916 12696
rect 10502 12628 10508 12640
rect 10152 12600 10508 12628
rect 8389 12591 8447 12597
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 10597 12631 10655 12637
rect 10597 12597 10609 12631
rect 10643 12628 10655 12631
rect 10689 12631 10747 12637
rect 10689 12628 10701 12631
rect 10643 12600 10701 12628
rect 10643 12597 10655 12600
rect 10597 12591 10655 12597
rect 10689 12597 10701 12600
rect 10735 12597 10747 12631
rect 10689 12591 10747 12597
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 11348 12628 11376 12727
rect 11422 12724 11428 12776
rect 11480 12764 11486 12776
rect 11808 12773 11836 12928
rect 12912 12912 12940 12940
rect 12618 12900 12624 12912
rect 11992 12872 12624 12900
rect 11882 12792 11888 12844
rect 11940 12832 11946 12844
rect 11992 12832 12020 12872
rect 12618 12860 12624 12872
rect 12676 12860 12682 12912
rect 12713 12903 12771 12909
rect 12713 12869 12725 12903
rect 12759 12869 12771 12903
rect 12713 12863 12771 12869
rect 11940 12804 12020 12832
rect 11940 12792 11946 12804
rect 11992 12773 12020 12804
rect 12342 12792 12348 12844
rect 12400 12792 12406 12844
rect 12728 12832 12756 12863
rect 12894 12860 12900 12912
rect 12952 12860 12958 12912
rect 12728 12804 14044 12832
rect 11517 12767 11575 12773
rect 11517 12764 11529 12767
rect 11480 12736 11529 12764
rect 11480 12724 11486 12736
rect 11517 12733 11529 12736
rect 11563 12733 11575 12767
rect 11517 12727 11575 12733
rect 11793 12767 11851 12773
rect 11793 12733 11805 12767
rect 11839 12733 11851 12767
rect 11793 12727 11851 12733
rect 11977 12767 12035 12773
rect 11977 12733 11989 12767
rect 12023 12733 12035 12767
rect 11977 12727 12035 12733
rect 12069 12767 12127 12773
rect 12069 12733 12081 12767
rect 12115 12733 12127 12767
rect 12069 12727 12127 12733
rect 12161 12767 12219 12773
rect 12161 12733 12173 12767
rect 12207 12764 12219 12767
rect 12360 12764 12388 12792
rect 12207 12736 12388 12764
rect 12437 12767 12495 12773
rect 12207 12733 12219 12736
rect 12161 12727 12219 12733
rect 12437 12733 12449 12767
rect 12483 12733 12495 12767
rect 12437 12727 12495 12733
rect 12529 12767 12587 12773
rect 12529 12733 12541 12767
rect 12575 12764 12587 12767
rect 13173 12767 13231 12773
rect 13173 12764 13185 12767
rect 12575 12736 13185 12764
rect 12575 12733 12587 12736
rect 12529 12727 12587 12733
rect 13173 12733 13185 12736
rect 13219 12733 13231 12767
rect 13173 12727 13231 12733
rect 13817 12767 13875 12773
rect 13817 12733 13829 12767
rect 13863 12733 13875 12767
rect 13817 12727 13875 12733
rect 11701 12699 11759 12705
rect 11701 12665 11713 12699
rect 11747 12696 11759 12699
rect 12084 12696 12112 12727
rect 11747 12668 12112 12696
rect 11747 12665 11759 12668
rect 11701 12659 11759 12665
rect 12250 12656 12256 12708
rect 12308 12696 12314 12708
rect 12345 12699 12403 12705
rect 12345 12696 12357 12699
rect 12308 12668 12357 12696
rect 12308 12656 12314 12668
rect 12345 12665 12357 12668
rect 12391 12665 12403 12699
rect 12452 12696 12480 12727
rect 12452 12668 12572 12696
rect 12345 12659 12403 12665
rect 11296 12600 11376 12628
rect 11885 12631 11943 12637
rect 11296 12588 11302 12600
rect 11885 12597 11897 12631
rect 11931 12628 11943 12631
rect 11974 12628 11980 12640
rect 11931 12600 11980 12628
rect 11931 12597 11943 12600
rect 11885 12591 11943 12597
rect 11974 12588 11980 12600
rect 12032 12628 12038 12640
rect 12544 12628 12572 12668
rect 12618 12656 12624 12708
rect 12676 12696 12682 12708
rect 12805 12699 12863 12705
rect 12805 12696 12817 12699
rect 12676 12668 12817 12696
rect 12676 12656 12682 12668
rect 12805 12665 12817 12668
rect 12851 12665 12863 12699
rect 12805 12659 12863 12665
rect 12894 12656 12900 12708
rect 12952 12696 12958 12708
rect 12989 12699 13047 12705
rect 12989 12696 13001 12699
rect 12952 12668 13001 12696
rect 12952 12656 12958 12668
rect 12989 12665 13001 12668
rect 13035 12696 13047 12699
rect 13832 12696 13860 12727
rect 13906 12724 13912 12776
rect 13964 12724 13970 12776
rect 14016 12773 14044 12804
rect 14001 12767 14059 12773
rect 14001 12733 14013 12767
rect 14047 12733 14059 12767
rect 14001 12727 14059 12733
rect 14182 12724 14188 12776
rect 14240 12764 14246 12776
rect 14642 12764 14648 12776
rect 14240 12736 14648 12764
rect 14240 12724 14246 12736
rect 14642 12724 14648 12736
rect 14700 12724 14706 12776
rect 15102 12724 15108 12776
rect 15160 12724 15166 12776
rect 15120 12696 15148 12724
rect 13035 12668 15148 12696
rect 13035 12665 13047 12668
rect 12989 12659 13047 12665
rect 12032 12600 12572 12628
rect 13541 12631 13599 12637
rect 12032 12588 12038 12600
rect 13541 12597 13553 12631
rect 13587 12628 13599 12631
rect 13630 12628 13636 12640
rect 13587 12600 13636 12628
rect 13587 12597 13599 12600
rect 13541 12591 13599 12597
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 552 12538 15520 12560
rect 552 12486 4100 12538
rect 4152 12486 4164 12538
rect 4216 12486 4228 12538
rect 4280 12486 4292 12538
rect 4344 12486 4356 12538
rect 4408 12486 7802 12538
rect 7854 12486 7866 12538
rect 7918 12486 7930 12538
rect 7982 12486 7994 12538
rect 8046 12486 8058 12538
rect 8110 12486 11504 12538
rect 11556 12486 11568 12538
rect 11620 12486 11632 12538
rect 11684 12486 11696 12538
rect 11748 12486 11760 12538
rect 11812 12486 15206 12538
rect 15258 12486 15270 12538
rect 15322 12486 15334 12538
rect 15386 12486 15398 12538
rect 15450 12486 15462 12538
rect 15514 12486 15520 12538
rect 552 12464 15520 12486
rect 4249 12427 4307 12433
rect 4249 12393 4261 12427
rect 4295 12424 4307 12427
rect 4430 12424 4436 12436
rect 4295 12396 4436 12424
rect 4295 12393 4307 12396
rect 4249 12387 4307 12393
rect 4430 12384 4436 12396
rect 4488 12384 4494 12436
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 11882 12424 11888 12436
rect 8904 12396 11888 12424
rect 8904 12384 8910 12396
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 11974 12384 11980 12436
rect 12032 12384 12038 12436
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 12621 12427 12679 12433
rect 12621 12424 12633 12427
rect 12584 12396 12633 12424
rect 12584 12384 12590 12396
rect 12621 12393 12633 12396
rect 12667 12393 12679 12427
rect 12621 12387 12679 12393
rect 5350 12356 5356 12368
rect 4540 12328 5356 12356
rect 4540 12297 4568 12328
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 4525 12291 4583 12297
rect 4525 12257 4537 12291
rect 4571 12257 4583 12291
rect 4525 12251 4583 12257
rect 4801 12291 4859 12297
rect 4801 12257 4813 12291
rect 4847 12257 4859 12291
rect 4801 12251 4859 12257
rect 4816 12220 4844 12251
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 7837 12291 7895 12297
rect 7837 12288 7849 12291
rect 7064 12260 7849 12288
rect 7064 12248 7070 12260
rect 7837 12257 7849 12260
rect 7883 12257 7895 12291
rect 7837 12251 7895 12257
rect 8110 12248 8116 12300
rect 8168 12248 8174 12300
rect 8202 12248 8208 12300
rect 8260 12248 8266 12300
rect 11992 12288 12020 12384
rect 15013 12359 15071 12365
rect 15013 12325 15025 12359
rect 15059 12356 15071 12359
rect 15102 12356 15108 12368
rect 15059 12328 15108 12356
rect 15059 12325 15071 12328
rect 15013 12319 15071 12325
rect 15102 12316 15108 12328
rect 15160 12316 15166 12368
rect 12437 12291 12495 12297
rect 12437 12288 12449 12291
rect 11992 12260 12449 12288
rect 12437 12257 12449 12260
rect 12483 12257 12495 12291
rect 12437 12251 12495 12257
rect 13262 12248 13268 12300
rect 13320 12288 13326 12300
rect 13357 12291 13415 12297
rect 13357 12288 13369 12291
rect 13320 12260 13369 12288
rect 13320 12248 13326 12260
rect 13357 12257 13369 12260
rect 13403 12257 13415 12291
rect 13357 12251 13415 12257
rect 13630 12248 13636 12300
rect 13688 12248 13694 12300
rect 3896 12192 4844 12220
rect 3896 12096 3924 12192
rect 7374 12180 7380 12232
rect 7432 12220 7438 12232
rect 7929 12223 7987 12229
rect 7929 12220 7941 12223
rect 7432 12192 7941 12220
rect 7432 12180 7438 12192
rect 7929 12189 7941 12192
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12220 8539 12223
rect 8570 12220 8576 12232
rect 8527 12192 8576 12220
rect 8527 12189 8539 12192
rect 8481 12183 8539 12189
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 8846 12180 8852 12232
rect 8904 12220 8910 12232
rect 9493 12223 9551 12229
rect 9493 12220 9505 12223
rect 8904 12192 9505 12220
rect 8904 12180 8910 12192
rect 9493 12189 9505 12192
rect 9539 12189 9551 12223
rect 9493 12183 9551 12189
rect 11422 12180 11428 12232
rect 11480 12220 11486 12232
rect 12250 12220 12256 12232
rect 11480 12192 12256 12220
rect 11480 12180 11486 12192
rect 12250 12180 12256 12192
rect 12308 12180 12314 12232
rect 8662 12152 8668 12164
rect 3988 12124 8668 12152
rect 3988 12096 4016 12124
rect 8662 12112 8668 12124
rect 8720 12112 8726 12164
rect 8754 12112 8760 12164
rect 8812 12152 8818 12164
rect 9122 12152 9128 12164
rect 8812 12124 9128 12152
rect 8812 12112 8818 12124
rect 9122 12112 9128 12124
rect 9180 12112 9186 12164
rect 9861 12155 9919 12161
rect 9861 12121 9873 12155
rect 9907 12152 9919 12155
rect 10410 12152 10416 12164
rect 9907 12124 10416 12152
rect 9907 12121 9919 12124
rect 9861 12115 9919 12121
rect 10410 12112 10416 12124
rect 10468 12112 10474 12164
rect 3878 12044 3884 12096
rect 3936 12044 3942 12096
rect 3970 12044 3976 12096
rect 4028 12044 4034 12096
rect 4709 12087 4767 12093
rect 4709 12053 4721 12087
rect 4755 12084 4767 12087
rect 4890 12084 4896 12096
rect 4755 12056 4896 12084
rect 4755 12053 4767 12056
rect 4709 12047 4767 12053
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 8386 12044 8392 12096
rect 8444 12044 8450 12096
rect 8941 12087 8999 12093
rect 8941 12053 8953 12087
rect 8987 12084 8999 12087
rect 9214 12084 9220 12096
rect 8987 12056 9220 12084
rect 8987 12053 8999 12056
rect 8941 12047 8999 12053
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 9398 12044 9404 12096
rect 9456 12084 9462 12096
rect 9953 12087 10011 12093
rect 9953 12084 9965 12087
rect 9456 12056 9965 12084
rect 9456 12044 9462 12056
rect 9953 12053 9965 12056
rect 9999 12053 10011 12087
rect 9953 12047 10011 12053
rect 552 11994 15364 12016
rect 552 11942 2249 11994
rect 2301 11942 2313 11994
rect 2365 11942 2377 11994
rect 2429 11942 2441 11994
rect 2493 11942 2505 11994
rect 2557 11942 5951 11994
rect 6003 11942 6015 11994
rect 6067 11942 6079 11994
rect 6131 11942 6143 11994
rect 6195 11942 6207 11994
rect 6259 11942 9653 11994
rect 9705 11942 9717 11994
rect 9769 11942 9781 11994
rect 9833 11942 9845 11994
rect 9897 11942 9909 11994
rect 9961 11942 13355 11994
rect 13407 11942 13419 11994
rect 13471 11942 13483 11994
rect 13535 11942 13547 11994
rect 13599 11942 13611 11994
rect 13663 11942 15364 11994
rect 552 11920 15364 11942
rect 7374 11880 7380 11892
rect 7116 11852 7380 11880
rect 6641 11815 6699 11821
rect 6641 11781 6653 11815
rect 6687 11812 6699 11815
rect 6914 11812 6920 11824
rect 6687 11784 6920 11812
rect 6687 11781 6699 11784
rect 6641 11775 6699 11781
rect 6914 11772 6920 11784
rect 6972 11772 6978 11824
rect 3234 11704 3240 11756
rect 3292 11744 3298 11756
rect 3878 11744 3884 11756
rect 3292 11716 3884 11744
rect 3292 11704 3298 11716
rect 3878 11704 3884 11716
rect 3936 11704 3942 11756
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11744 4399 11747
rect 4982 11744 4988 11756
rect 4387 11716 4988 11744
rect 4387 11713 4399 11716
rect 4341 11707 4399 11713
rect 4982 11704 4988 11716
rect 5040 11744 5046 11756
rect 5040 11716 5488 11744
rect 5040 11704 5046 11716
rect 3970 11636 3976 11688
rect 4028 11636 4034 11688
rect 4614 11636 4620 11688
rect 4672 11676 4678 11688
rect 5077 11679 5135 11685
rect 5077 11676 5089 11679
rect 4672 11648 5089 11676
rect 4672 11636 4678 11648
rect 5077 11645 5089 11648
rect 5123 11645 5135 11679
rect 5077 11639 5135 11645
rect 5261 11679 5319 11685
rect 5261 11645 5273 11679
rect 5307 11645 5319 11679
rect 5261 11639 5319 11645
rect 5276 11608 5304 11639
rect 5350 11636 5356 11688
rect 5408 11636 5414 11688
rect 5460 11685 5488 11716
rect 7006 11685 7012 11688
rect 5445 11679 5503 11685
rect 5445 11645 5457 11679
rect 5491 11645 5503 11679
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 5445 11639 5503 11645
rect 6748 11648 6837 11676
rect 5626 11608 5632 11620
rect 5276 11580 5632 11608
rect 5626 11568 5632 11580
rect 5684 11568 5690 11620
rect 6270 11568 6276 11620
rect 6328 11568 6334 11620
rect 5718 11500 5724 11552
rect 5776 11500 5782 11552
rect 5994 11500 6000 11552
rect 6052 11540 6058 11552
rect 6748 11549 6776 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 6973 11679 7012 11685
rect 6973 11645 6985 11679
rect 6973 11639 7012 11645
rect 7006 11636 7012 11639
rect 7064 11636 7070 11688
rect 7116 11685 7144 11852
rect 7374 11840 7380 11852
rect 7432 11840 7438 11892
rect 8202 11840 8208 11892
rect 8260 11840 8266 11892
rect 8662 11840 8668 11892
rect 8720 11880 8726 11892
rect 9306 11880 9312 11892
rect 8720 11852 9312 11880
rect 8720 11840 8726 11852
rect 9306 11840 9312 11852
rect 9364 11880 9370 11892
rect 9364 11852 11192 11880
rect 9364 11840 9370 11852
rect 7282 11772 7288 11824
rect 7340 11812 7346 11824
rect 8220 11812 8248 11840
rect 7340 11784 8156 11812
rect 8220 11784 8524 11812
rect 7340 11772 7346 11784
rect 8128 11753 8156 11784
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 8294 11704 8300 11756
rect 8352 11704 8358 11756
rect 7101 11679 7159 11685
rect 7101 11645 7113 11679
rect 7147 11645 7159 11679
rect 7101 11639 7159 11645
rect 7331 11679 7389 11685
rect 7331 11645 7343 11679
rect 7377 11676 7389 11679
rect 7466 11676 7472 11688
rect 7377 11648 7472 11676
rect 7377 11645 7389 11648
rect 7331 11639 7389 11645
rect 7466 11636 7472 11648
rect 7524 11676 7530 11688
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 7524 11648 7757 11676
rect 7524 11636 7530 11648
rect 7745 11645 7757 11648
rect 7791 11645 7803 11679
rect 7745 11639 7803 11645
rect 7837 11679 7895 11685
rect 7837 11645 7849 11679
rect 7883 11645 7895 11679
rect 7837 11639 7895 11645
rect 7193 11611 7251 11617
rect 7193 11577 7205 11611
rect 7239 11608 7251 11611
rect 7852 11608 7880 11639
rect 7239 11580 7880 11608
rect 7239 11577 7251 11580
rect 7193 11571 7251 11577
rect 7668 11552 7696 11580
rect 8110 11568 8116 11620
rect 8168 11568 8174 11620
rect 8205 11611 8263 11617
rect 8205 11577 8217 11611
rect 8251 11608 8263 11611
rect 8312 11608 8340 11704
rect 8496 11676 8524 11784
rect 9140 11716 9444 11744
rect 9140 11685 9168 11716
rect 9416 11688 9444 11716
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 9677 11747 9735 11753
rect 9677 11744 9689 11747
rect 9548 11716 9689 11744
rect 9548 11704 9554 11716
rect 9677 11713 9689 11716
rect 9723 11713 9735 11747
rect 9677 11707 9735 11713
rect 11164 11744 11192 11852
rect 12618 11840 12624 11892
rect 12676 11880 12682 11892
rect 12713 11883 12771 11889
rect 12713 11880 12725 11883
rect 12676 11852 12725 11880
rect 12676 11840 12682 11852
rect 12713 11849 12725 11852
rect 12759 11849 12771 11883
rect 12713 11843 12771 11849
rect 12894 11840 12900 11892
rect 12952 11840 12958 11892
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11164 11716 11713 11744
rect 8711 11679 8769 11685
rect 8711 11676 8723 11679
rect 8496 11648 8723 11676
rect 8711 11645 8723 11648
rect 8757 11645 8769 11679
rect 8711 11639 8769 11645
rect 9124 11679 9182 11685
rect 9124 11645 9136 11679
rect 9170 11645 9182 11679
rect 9124 11639 9182 11645
rect 9214 11636 9220 11688
rect 9272 11636 9278 11688
rect 9398 11636 9404 11688
rect 9456 11636 9462 11688
rect 8849 11611 8907 11617
rect 8849 11608 8861 11611
rect 8251 11580 8340 11608
rect 8404 11580 8861 11608
rect 8251 11577 8263 11580
rect 8205 11571 8263 11577
rect 6733 11543 6791 11549
rect 6733 11540 6745 11543
rect 6052 11512 6745 11540
rect 6052 11500 6058 11512
rect 6733 11509 6745 11512
rect 6779 11509 6791 11543
rect 6733 11503 6791 11509
rect 7466 11500 7472 11552
rect 7524 11500 7530 11552
rect 7558 11500 7564 11552
rect 7616 11500 7622 11552
rect 7650 11500 7656 11552
rect 7708 11500 7714 11552
rect 8128 11540 8156 11568
rect 8404 11540 8432 11580
rect 8849 11577 8861 11580
rect 8895 11577 8907 11611
rect 8849 11571 8907 11577
rect 8938 11568 8944 11620
rect 8996 11568 9002 11620
rect 9674 11568 9680 11620
rect 9732 11608 9738 11620
rect 9922 11611 9980 11617
rect 9922 11608 9934 11611
rect 9732 11580 9934 11608
rect 9732 11568 9738 11580
rect 9922 11577 9934 11580
rect 9968 11577 9980 11611
rect 11164 11608 11192 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11238 11636 11244 11688
rect 11296 11676 11302 11688
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 11296 11648 12081 11676
rect 11296 11636 11302 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11676 12311 11679
rect 12636 11676 12664 11840
rect 12299 11648 12664 11676
rect 13817 11679 13875 11685
rect 12299 11645 12311 11648
rect 12253 11639 12311 11645
rect 13817 11645 13829 11679
rect 13863 11645 13875 11679
rect 13817 11639 13875 11645
rect 9922 11571 9980 11577
rect 11072 11580 11192 11608
rect 8128 11512 8432 11540
rect 8570 11500 8576 11552
rect 8628 11500 8634 11552
rect 11072 11549 11100 11580
rect 13078 11568 13084 11620
rect 13136 11608 13142 11620
rect 13832 11608 13860 11639
rect 13906 11636 13912 11688
rect 13964 11636 13970 11688
rect 13998 11636 14004 11688
rect 14056 11636 14062 11688
rect 14182 11636 14188 11688
rect 14240 11636 14246 11688
rect 13136 11580 13860 11608
rect 13136 11568 13142 11580
rect 11057 11543 11115 11549
rect 11057 11509 11069 11543
rect 11103 11509 11115 11543
rect 11057 11503 11115 11509
rect 11146 11500 11152 11552
rect 11204 11500 11210 11552
rect 12161 11543 12219 11549
rect 12161 11509 12173 11543
rect 12207 11540 12219 11543
rect 12434 11540 12440 11552
rect 12207 11512 12440 11540
rect 12207 11509 12219 11512
rect 12161 11503 12219 11509
rect 12434 11500 12440 11512
rect 12492 11500 12498 11552
rect 12894 11549 12900 11552
rect 12881 11543 12900 11549
rect 12881 11509 12893 11543
rect 12881 11503 12900 11509
rect 12894 11500 12900 11503
rect 12952 11500 12958 11552
rect 13541 11543 13599 11549
rect 13541 11509 13553 11543
rect 13587 11540 13599 11543
rect 13630 11540 13636 11552
rect 13587 11512 13636 11540
rect 13587 11509 13599 11512
rect 13541 11503 13599 11509
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 552 11450 15520 11472
rect 552 11398 4100 11450
rect 4152 11398 4164 11450
rect 4216 11398 4228 11450
rect 4280 11398 4292 11450
rect 4344 11398 4356 11450
rect 4408 11398 7802 11450
rect 7854 11398 7866 11450
rect 7918 11398 7930 11450
rect 7982 11398 7994 11450
rect 8046 11398 8058 11450
rect 8110 11398 11504 11450
rect 11556 11398 11568 11450
rect 11620 11398 11632 11450
rect 11684 11398 11696 11450
rect 11748 11398 11760 11450
rect 11812 11398 15206 11450
rect 15258 11398 15270 11450
rect 15322 11398 15334 11450
rect 15386 11398 15398 11450
rect 15450 11398 15462 11450
rect 15514 11398 15520 11450
rect 552 11376 15520 11398
rect 3970 11296 3976 11348
rect 4028 11296 4034 11348
rect 4249 11339 4307 11345
rect 4249 11305 4261 11339
rect 4295 11336 4307 11339
rect 4614 11336 4620 11348
rect 4295 11308 4620 11336
rect 4295 11305 4307 11308
rect 4249 11299 4307 11305
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 4801 11339 4859 11345
rect 4801 11305 4813 11339
rect 4847 11336 4859 11339
rect 5350 11336 5356 11348
rect 4847 11308 5356 11336
rect 4847 11305 4859 11308
rect 4801 11299 4859 11305
rect 3789 11203 3847 11209
rect 3789 11169 3801 11203
rect 3835 11200 3847 11203
rect 3988 11200 4016 11296
rect 3835 11172 4016 11200
rect 3835 11169 3847 11172
rect 3789 11163 3847 11169
rect 4338 11160 4344 11212
rect 4396 11160 4402 11212
rect 4908 11209 4936 11308
rect 5350 11296 5356 11308
rect 5408 11296 5414 11348
rect 7374 11336 7380 11348
rect 6656 11308 7380 11336
rect 4893 11203 4951 11209
rect 4893 11169 4905 11203
rect 4939 11169 4951 11203
rect 4893 11163 4951 11169
rect 5718 11160 5724 11212
rect 5776 11200 5782 11212
rect 5905 11203 5963 11209
rect 5905 11200 5917 11203
rect 5776 11172 5917 11200
rect 5776 11160 5782 11172
rect 5905 11169 5917 11172
rect 5951 11169 5963 11203
rect 5905 11163 5963 11169
rect 5994 11160 6000 11212
rect 6052 11160 6058 11212
rect 6656 11209 6684 11308
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 7745 11339 7803 11345
rect 7745 11305 7757 11339
rect 7791 11336 7803 11339
rect 8570 11336 8576 11348
rect 7791 11308 8576 11336
rect 7791 11305 7803 11308
rect 7745 11299 7803 11305
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 8938 11296 8944 11348
rect 8996 11296 9002 11348
rect 9674 11296 9680 11348
rect 9732 11296 9738 11348
rect 11882 11296 11888 11348
rect 11940 11296 11946 11348
rect 12989 11339 13047 11345
rect 12989 11305 13001 11339
rect 13035 11336 13047 11339
rect 13998 11336 14004 11348
rect 13035 11308 14004 11336
rect 13035 11305 13047 11308
rect 12989 11299 13047 11305
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 6748 11240 7696 11268
rect 6748 11209 6776 11240
rect 7668 11212 7696 11240
rect 8662 11228 8668 11280
rect 8720 11228 8726 11280
rect 10505 11271 10563 11277
rect 10505 11268 10517 11271
rect 9876 11240 10517 11268
rect 6181 11203 6239 11209
rect 6181 11169 6193 11203
rect 6227 11169 6239 11203
rect 6181 11163 6239 11169
rect 6641 11203 6699 11209
rect 6641 11169 6653 11203
rect 6687 11169 6699 11203
rect 6641 11163 6699 11169
rect 6733 11203 6791 11209
rect 6733 11169 6745 11203
rect 6779 11169 6791 11203
rect 6733 11163 6791 11169
rect 5166 11092 5172 11144
rect 5224 11092 5230 11144
rect 6196 11132 6224 11163
rect 7006 11160 7012 11212
rect 7064 11160 7070 11212
rect 7377 11203 7435 11209
rect 7377 11169 7389 11203
rect 7423 11200 7435 11203
rect 7466 11200 7472 11212
rect 7423 11172 7472 11200
rect 7423 11169 7435 11172
rect 7377 11163 7435 11169
rect 7466 11160 7472 11172
rect 7524 11160 7530 11212
rect 7558 11160 7564 11212
rect 7616 11160 7622 11212
rect 7650 11160 7656 11212
rect 7708 11160 7714 11212
rect 7837 11203 7895 11209
rect 7837 11169 7849 11203
rect 7883 11200 7895 11203
rect 8386 11200 8392 11212
rect 7883 11172 8392 11200
rect 7883 11169 7895 11172
rect 7837 11163 7895 11169
rect 8386 11160 8392 11172
rect 8444 11160 8450 11212
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11200 8539 11203
rect 8680 11200 8708 11228
rect 9876 11209 9904 11240
rect 10505 11237 10517 11240
rect 10551 11237 10563 11271
rect 10505 11231 10563 11237
rect 12084 11240 12848 11268
rect 12084 11212 12112 11240
rect 8527 11172 8708 11200
rect 9861 11203 9919 11209
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 9861 11169 9873 11203
rect 9907 11169 9919 11203
rect 9861 11163 9919 11169
rect 5460 11104 7328 11132
rect 5460 11073 5488 11104
rect 5445 11067 5503 11073
rect 5445 11033 5457 11067
rect 5491 11033 5503 11067
rect 5445 11027 5503 11033
rect 6089 11067 6147 11073
rect 6089 11033 6101 11067
rect 6135 11064 6147 11067
rect 6457 11067 6515 11073
rect 6457 11064 6469 11067
rect 6135 11036 6469 11064
rect 6135 11033 6147 11036
rect 6089 11027 6147 11033
rect 6457 11033 6469 11036
rect 6503 11033 6515 11067
rect 6457 11027 6515 11033
rect 6914 11024 6920 11076
rect 6972 11024 6978 11076
rect 3878 10956 3884 11008
rect 3936 10956 3942 11008
rect 4617 10999 4675 11005
rect 4617 10965 4629 10999
rect 4663 10996 4675 10999
rect 4798 10996 4804 11008
rect 4663 10968 4804 10996
rect 4663 10965 4675 10968
rect 4617 10959 4675 10965
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 4982 10956 4988 11008
rect 5040 10956 5046 11008
rect 6362 10956 6368 11008
rect 6420 10956 6426 11008
rect 7101 10999 7159 11005
rect 7101 10965 7113 10999
rect 7147 10996 7159 10999
rect 7190 10996 7196 11008
rect 7147 10968 7196 10996
rect 7147 10965 7159 10968
rect 7101 10959 7159 10965
rect 7190 10956 7196 10968
rect 7248 10956 7254 11008
rect 7300 10996 7328 11104
rect 7469 11067 7527 11073
rect 7469 11033 7481 11067
rect 7515 11064 7527 11067
rect 7576 11064 7604 11160
rect 7515 11036 7604 11064
rect 7515 11033 7527 11036
rect 7469 11027 7527 11033
rect 8386 11024 8392 11076
rect 8444 11064 8450 11076
rect 8496 11064 8524 11163
rect 10134 11160 10140 11212
rect 10192 11160 10198 11212
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11169 10379 11203
rect 10321 11163 10379 11169
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11200 10655 11203
rect 11146 11200 11152 11212
rect 10643 11172 11152 11200
rect 10643 11169 10655 11172
rect 10597 11163 10655 11169
rect 8444 11036 8524 11064
rect 8444 11024 8450 11036
rect 9490 11024 9496 11076
rect 9548 11064 9554 11076
rect 9953 11067 10011 11073
rect 9953 11064 9965 11067
rect 9548 11036 9965 11064
rect 9548 11024 9554 11036
rect 9953 11033 9965 11036
rect 9999 11033 10011 11067
rect 9953 11027 10011 11033
rect 10042 11024 10048 11076
rect 10100 11024 10106 11076
rect 10336 11008 10364 11163
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 12066 11160 12072 11212
rect 12124 11160 12130 11212
rect 12342 11160 12348 11212
rect 12400 11160 12406 11212
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 12492 11172 12537 11200
rect 12492 11160 12498 11172
rect 12618 11160 12624 11212
rect 12676 11160 12682 11212
rect 12710 11160 12716 11212
rect 12768 11160 12774 11212
rect 12820 11209 12848 11240
rect 12810 11203 12868 11209
rect 12810 11169 12822 11203
rect 12856 11169 12868 11203
rect 12810 11163 12868 11169
rect 13262 11160 13268 11212
rect 13320 11200 13326 11212
rect 13357 11203 13415 11209
rect 13357 11200 13369 11203
rect 13320 11172 13369 11200
rect 13320 11160 13326 11172
rect 13357 11169 13369 11172
rect 13403 11169 13415 11203
rect 13357 11163 13415 11169
rect 13630 11160 13636 11212
rect 13688 11160 13694 11212
rect 11422 11092 11428 11144
rect 11480 11132 11486 11144
rect 11609 11135 11667 11141
rect 11609 11132 11621 11135
rect 11480 11104 11621 11132
rect 11480 11092 11486 11104
rect 11609 11101 11621 11104
rect 11655 11101 11667 11135
rect 11609 11095 11667 11101
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11132 11851 11135
rect 13170 11132 13176 11144
rect 11839 11104 13176 11132
rect 11839 11101 11851 11104
rect 11793 11095 11851 11101
rect 13170 11092 13176 11104
rect 13228 11092 13234 11144
rect 15102 11132 15108 11144
rect 13280 11104 15108 11132
rect 13078 11024 13084 11076
rect 13136 11064 13142 11076
rect 13280 11064 13308 11104
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 13136 11036 13308 11064
rect 13136 11024 13142 11036
rect 7561 10999 7619 11005
rect 7561 10996 7573 10999
rect 7300 10968 7573 10996
rect 7561 10965 7573 10968
rect 7607 10965 7619 10999
rect 7561 10959 7619 10965
rect 8754 10956 8760 11008
rect 8812 10956 8818 11008
rect 9398 10956 9404 11008
rect 9456 10996 9462 11008
rect 10318 10996 10324 11008
rect 9456 10968 10324 10996
rect 9456 10956 9462 10968
rect 10318 10956 10324 10968
rect 10376 10956 10382 11008
rect 12253 10999 12311 11005
rect 12253 10965 12265 10999
rect 12299 10996 12311 10999
rect 12434 10996 12440 11008
rect 12299 10968 12440 10996
rect 12299 10965 12311 10968
rect 12253 10959 12311 10965
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 14921 10999 14979 11005
rect 14921 10965 14933 10999
rect 14967 10996 14979 10999
rect 15102 10996 15108 11008
rect 14967 10968 15108 10996
rect 14967 10965 14979 10968
rect 14921 10959 14979 10965
rect 15102 10956 15108 10968
rect 15160 10956 15166 11008
rect 552 10906 15364 10928
rect 552 10854 2249 10906
rect 2301 10854 2313 10906
rect 2365 10854 2377 10906
rect 2429 10854 2441 10906
rect 2493 10854 2505 10906
rect 2557 10854 5951 10906
rect 6003 10854 6015 10906
rect 6067 10854 6079 10906
rect 6131 10854 6143 10906
rect 6195 10854 6207 10906
rect 6259 10854 9653 10906
rect 9705 10854 9717 10906
rect 9769 10854 9781 10906
rect 9833 10854 9845 10906
rect 9897 10854 9909 10906
rect 9961 10854 13355 10906
rect 13407 10854 13419 10906
rect 13471 10854 13483 10906
rect 13535 10854 13547 10906
rect 13599 10854 13611 10906
rect 13663 10854 15364 10906
rect 552 10832 15364 10854
rect 4985 10795 5043 10801
rect 4985 10761 4997 10795
rect 5031 10792 5043 10795
rect 5166 10792 5172 10804
rect 5031 10764 5172 10792
rect 5031 10761 5043 10764
rect 4985 10755 5043 10761
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5258 10752 5264 10804
rect 5316 10792 5322 10804
rect 5537 10795 5595 10801
rect 5537 10792 5549 10795
rect 5316 10764 5549 10792
rect 5316 10752 5322 10764
rect 5537 10761 5549 10764
rect 5583 10761 5595 10795
rect 5537 10755 5595 10761
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10321 10795 10379 10801
rect 10321 10792 10333 10795
rect 10192 10764 10333 10792
rect 10192 10752 10198 10764
rect 10321 10761 10333 10764
rect 10367 10761 10379 10795
rect 10321 10755 10379 10761
rect 12618 10752 12624 10804
rect 12676 10752 12682 10804
rect 13078 10792 13084 10804
rect 12728 10764 13084 10792
rect 4798 10684 4804 10736
rect 4856 10684 4862 10736
rect 8570 10684 8576 10736
rect 8628 10724 8634 10736
rect 8628 10696 10088 10724
rect 8628 10684 8634 10696
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 4525 10659 4583 10665
rect 4525 10656 4537 10659
rect 4396 10628 4537 10656
rect 4396 10616 4402 10628
rect 4525 10625 4537 10628
rect 4571 10656 4583 10659
rect 8662 10656 8668 10668
rect 4571 10628 8668 10656
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 8662 10616 8668 10628
rect 8720 10656 8726 10668
rect 10060 10665 10088 10696
rect 9953 10659 10011 10665
rect 9953 10656 9965 10659
rect 8720 10628 9965 10656
rect 8720 10616 8726 10628
rect 9953 10625 9965 10628
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10656 10103 10659
rect 12342 10656 12348 10668
rect 10091 10628 12348 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 12342 10616 12348 10628
rect 12400 10616 12406 10668
rect 9306 10548 9312 10600
rect 9364 10588 9370 10600
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9364 10560 9873 10588
rect 9364 10548 9370 10560
rect 9861 10557 9873 10560
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 10134 10548 10140 10600
rect 10192 10548 10198 10600
rect 12728 10588 12756 10764
rect 13078 10752 13084 10764
rect 13136 10752 13142 10804
rect 13170 10752 13176 10804
rect 13228 10792 13234 10804
rect 13265 10795 13323 10801
rect 13265 10792 13277 10795
rect 13228 10764 13277 10792
rect 13228 10752 13234 10764
rect 13265 10761 13277 10764
rect 13311 10761 13323 10795
rect 13265 10755 13323 10761
rect 12802 10684 12808 10736
rect 12860 10684 12866 10736
rect 12820 10656 12848 10684
rect 12820 10628 13216 10656
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12728 10560 12817 10588
rect 12805 10557 12817 10560
rect 12851 10557 12863 10591
rect 12805 10551 12863 10557
rect 12894 10548 12900 10600
rect 12952 10588 12958 10600
rect 13078 10588 13084 10600
rect 12952 10560 13084 10588
rect 12952 10548 12958 10560
rect 13078 10548 13084 10560
rect 13136 10548 13142 10600
rect 13188 10597 13216 10628
rect 13173 10591 13231 10597
rect 13173 10557 13185 10591
rect 13219 10557 13231 10591
rect 13173 10551 13231 10557
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10557 13415 10591
rect 13357 10551 13415 10557
rect 7009 10523 7067 10529
rect 7009 10489 7021 10523
rect 7055 10520 7067 10523
rect 8938 10520 8944 10532
rect 7055 10492 8944 10520
rect 7055 10489 7067 10492
rect 7009 10483 7067 10489
rect 8938 10480 8944 10492
rect 8996 10520 9002 10532
rect 10413 10523 10471 10529
rect 10413 10520 10425 10523
rect 8996 10492 10425 10520
rect 8996 10480 9002 10492
rect 10413 10489 10425 10492
rect 10459 10489 10471 10523
rect 10413 10483 10471 10489
rect 12066 10480 12072 10532
rect 12124 10520 12130 10532
rect 12161 10523 12219 10529
rect 12161 10520 12173 10523
rect 12124 10492 12173 10520
rect 12124 10480 12130 10492
rect 12161 10489 12173 10492
rect 12207 10520 12219 10523
rect 13262 10520 13268 10532
rect 12207 10492 13268 10520
rect 12207 10489 12219 10492
rect 12161 10483 12219 10489
rect 13262 10480 13268 10492
rect 13320 10480 13326 10532
rect 6546 10412 6552 10464
rect 6604 10452 6610 10464
rect 10226 10452 10232 10464
rect 6604 10424 10232 10452
rect 6604 10412 6610 10424
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 12894 10412 12900 10464
rect 12952 10452 12958 10464
rect 12989 10455 13047 10461
rect 12989 10452 13001 10455
rect 12952 10424 13001 10452
rect 12952 10412 12958 10424
rect 12989 10421 13001 10424
rect 13035 10421 13047 10455
rect 12989 10415 13047 10421
rect 13078 10412 13084 10464
rect 13136 10452 13142 10464
rect 13372 10452 13400 10551
rect 13136 10424 13400 10452
rect 13136 10412 13142 10424
rect 552 10362 15520 10384
rect 552 10310 4100 10362
rect 4152 10310 4164 10362
rect 4216 10310 4228 10362
rect 4280 10310 4292 10362
rect 4344 10310 4356 10362
rect 4408 10310 7802 10362
rect 7854 10310 7866 10362
rect 7918 10310 7930 10362
rect 7982 10310 7994 10362
rect 8046 10310 8058 10362
rect 8110 10310 11504 10362
rect 11556 10310 11568 10362
rect 11620 10310 11632 10362
rect 11684 10310 11696 10362
rect 11748 10310 11760 10362
rect 11812 10310 15206 10362
rect 15258 10310 15270 10362
rect 15322 10310 15334 10362
rect 15386 10310 15398 10362
rect 15450 10310 15462 10362
rect 15514 10310 15520 10362
rect 552 10288 15520 10310
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 6546 10248 6552 10260
rect 5592 10220 6552 10248
rect 5592 10208 5598 10220
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7374 10248 7380 10260
rect 7064 10220 7380 10248
rect 7064 10208 7070 10220
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 7650 10208 7656 10260
rect 7708 10208 7714 10260
rect 8570 10208 8576 10260
rect 8628 10208 8634 10260
rect 8662 10208 8668 10260
rect 8720 10248 8726 10260
rect 9861 10251 9919 10257
rect 9861 10248 9873 10251
rect 8720 10220 9873 10248
rect 8720 10208 8726 10220
rect 9861 10217 9873 10220
rect 9907 10217 9919 10251
rect 9861 10211 9919 10217
rect 10870 10208 10876 10260
rect 10928 10248 10934 10260
rect 11425 10251 11483 10257
rect 11425 10248 11437 10251
rect 10928 10220 11437 10248
rect 10928 10208 10934 10220
rect 11425 10217 11437 10220
rect 11471 10217 11483 10251
rect 14090 10248 14096 10260
rect 11425 10211 11483 10217
rect 12360 10220 14096 10248
rect 5626 10140 5632 10192
rect 5684 10180 5690 10192
rect 5905 10183 5963 10189
rect 5905 10180 5917 10183
rect 5684 10152 5917 10180
rect 5684 10140 5690 10152
rect 5905 10149 5917 10152
rect 5951 10180 5963 10183
rect 6457 10183 6515 10189
rect 6457 10180 6469 10183
rect 5951 10152 6469 10180
rect 5951 10149 5963 10152
rect 5905 10143 5963 10149
rect 6457 10149 6469 10152
rect 6503 10149 6515 10183
rect 6457 10143 6515 10149
rect 5169 10115 5227 10121
rect 5169 10081 5181 10115
rect 5215 10081 5227 10115
rect 5169 10075 5227 10081
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10112 5411 10115
rect 5810 10112 5816 10124
rect 5399 10084 5816 10112
rect 5399 10081 5411 10084
rect 5353 10075 5411 10081
rect 5184 10044 5212 10075
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 6270 10072 6276 10124
rect 6328 10072 6334 10124
rect 6564 10121 6592 10208
rect 7558 10140 7564 10192
rect 7616 10180 7622 10192
rect 10134 10180 10140 10192
rect 7616 10152 10140 10180
rect 7616 10140 7622 10152
rect 6549 10115 6607 10121
rect 6549 10081 6561 10115
rect 6595 10081 6607 10115
rect 6549 10075 6607 10081
rect 7469 10115 7527 10121
rect 7469 10081 7481 10115
rect 7515 10081 7527 10115
rect 7469 10075 7527 10081
rect 5442 10044 5448 10056
rect 5184 10016 5448 10044
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 6288 10044 6316 10072
rect 6914 10044 6920 10056
rect 6288 10016 6920 10044
rect 6914 10004 6920 10016
rect 6972 10044 6978 10056
rect 7484 10044 7512 10075
rect 7742 10072 7748 10124
rect 7800 10072 7806 10124
rect 8478 10072 8484 10124
rect 8536 10072 8542 10124
rect 8662 10072 8668 10124
rect 8720 10112 8726 10124
rect 8757 10115 8815 10121
rect 8757 10112 8769 10115
rect 8720 10084 8769 10112
rect 8720 10072 8726 10084
rect 8757 10081 8769 10084
rect 8803 10081 8815 10115
rect 9033 10115 9091 10121
rect 9033 10112 9045 10115
rect 8757 10075 8815 10081
rect 8864 10084 9045 10112
rect 6972 10016 7512 10044
rect 6972 10004 6978 10016
rect 8864 9976 8892 10084
rect 9033 10081 9045 10084
rect 9079 10081 9091 10115
rect 9033 10075 9091 10081
rect 9217 10115 9275 10121
rect 9217 10081 9229 10115
rect 9263 10081 9275 10115
rect 9217 10075 9275 10081
rect 9309 10115 9367 10121
rect 9309 10081 9321 10115
rect 9355 10081 9367 10115
rect 9309 10075 9367 10081
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10044 8999 10047
rect 9232 10044 9260 10075
rect 8987 10016 9260 10044
rect 9324 10044 9352 10075
rect 9398 10072 9404 10124
rect 9456 10072 9462 10124
rect 9784 10121 9812 10152
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 10226 10140 10232 10192
rect 10284 10180 10290 10192
rect 11146 10180 11152 10192
rect 10284 10152 11152 10180
rect 10284 10140 10290 10152
rect 11146 10140 11152 10152
rect 11204 10180 11210 10192
rect 11333 10183 11391 10189
rect 11333 10180 11345 10183
rect 11204 10152 11345 10180
rect 11204 10140 11210 10152
rect 11333 10149 11345 10152
rect 11379 10180 11391 10183
rect 12158 10180 12164 10192
rect 11379 10152 12164 10180
rect 11379 10149 11391 10152
rect 11333 10143 11391 10149
rect 12158 10140 12164 10152
rect 12216 10140 12222 10192
rect 9769 10115 9827 10121
rect 9769 10081 9781 10115
rect 9815 10081 9827 10115
rect 9769 10075 9827 10081
rect 10045 10115 10103 10121
rect 10045 10081 10057 10115
rect 10091 10081 10103 10115
rect 10045 10075 10103 10081
rect 10060 10044 10088 10075
rect 10318 10072 10324 10124
rect 10376 10112 10382 10124
rect 12253 10115 12311 10121
rect 12253 10112 12265 10115
rect 10376 10084 12265 10112
rect 10376 10072 10382 10084
rect 12253 10081 12265 10084
rect 12299 10112 12311 10115
rect 12360 10112 12388 10220
rect 14090 10208 14096 10220
rect 14148 10208 14154 10260
rect 12544 10152 12940 10180
rect 12299 10084 12388 10112
rect 12299 10081 12311 10084
rect 12253 10075 12311 10081
rect 12434 10072 12440 10124
rect 12492 10072 12498 10124
rect 11054 10044 11060 10056
rect 9324 10016 9444 10044
rect 10060 10016 11060 10044
rect 8987 10013 8999 10016
rect 8941 10007 8999 10013
rect 9306 9976 9312 9988
rect 8864 9948 9312 9976
rect 9306 9936 9312 9948
rect 9364 9936 9370 9988
rect 5166 9868 5172 9920
rect 5224 9908 5230 9920
rect 5353 9911 5411 9917
rect 5353 9908 5365 9911
rect 5224 9880 5365 9908
rect 5224 9868 5230 9880
rect 5353 9877 5365 9880
rect 5399 9877 5411 9911
rect 5353 9871 5411 9877
rect 6181 9911 6239 9917
rect 6181 9877 6193 9911
rect 6227 9908 6239 9911
rect 6638 9908 6644 9920
rect 6227 9880 6644 9908
rect 6227 9877 6239 9880
rect 6181 9871 6239 9877
rect 6638 9868 6644 9880
rect 6696 9868 6702 9920
rect 9416 9908 9444 10016
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 12544 10053 12572 10152
rect 12802 10072 12808 10124
rect 12860 10072 12866 10124
rect 12912 10110 12940 10152
rect 13069 10118 13127 10121
rect 13004 10115 13127 10118
rect 13004 10110 13081 10115
rect 12912 10090 13081 10110
rect 12912 10082 13032 10090
rect 13069 10081 13081 10090
rect 13115 10081 13127 10115
rect 13069 10075 13127 10081
rect 13173 10115 13231 10121
rect 13173 10081 13185 10115
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 13265 10115 13323 10121
rect 13265 10081 13277 10115
rect 13311 10081 13323 10115
rect 13265 10075 13323 10081
rect 12529 10047 12587 10053
rect 12529 10044 12541 10047
rect 12452 10016 12541 10044
rect 9677 9979 9735 9985
rect 9677 9945 9689 9979
rect 9723 9976 9735 9979
rect 10134 9976 10140 9988
rect 9723 9948 10140 9976
rect 9723 9945 9735 9948
rect 9677 9939 9735 9945
rect 10134 9936 10140 9948
rect 10192 9936 10198 9988
rect 12452 9920 12480 10016
rect 12529 10013 12541 10016
rect 12575 10013 12587 10047
rect 12529 10007 12587 10013
rect 12621 10047 12679 10053
rect 12621 10013 12633 10047
rect 12667 10044 12679 10047
rect 13188 10044 13216 10075
rect 12667 10016 13216 10044
rect 12667 10013 12679 10016
rect 12621 10007 12679 10013
rect 12802 9936 12808 9988
rect 12860 9976 12866 9988
rect 12989 9979 13047 9985
rect 12860 9948 12940 9976
rect 12860 9936 12866 9948
rect 10042 9908 10048 9920
rect 9416 9880 10048 9908
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 12434 9868 12440 9920
rect 12492 9868 12498 9920
rect 12912 9908 12940 9948
rect 12989 9945 13001 9979
rect 13035 9945 13047 9979
rect 12989 9939 13047 9945
rect 13004 9908 13032 9939
rect 13170 9936 13176 9988
rect 13228 9976 13234 9988
rect 13280 9976 13308 10075
rect 13446 10072 13452 10124
rect 13504 10072 13510 10124
rect 13354 10004 13360 10056
rect 13412 10004 13418 10056
rect 13464 10044 13492 10072
rect 13633 10047 13691 10053
rect 13633 10044 13645 10047
rect 13464 10016 13645 10044
rect 13633 10013 13645 10016
rect 13679 10013 13691 10047
rect 13633 10007 13691 10013
rect 13228 9948 13308 9976
rect 13228 9936 13234 9948
rect 12912 9880 13032 9908
rect 14921 9911 14979 9917
rect 14921 9877 14933 9911
rect 14967 9908 14979 9911
rect 15102 9908 15108 9920
rect 14967 9880 15108 9908
rect 14967 9877 14979 9880
rect 14921 9871 14979 9877
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 552 9818 15364 9840
rect 552 9766 2249 9818
rect 2301 9766 2313 9818
rect 2365 9766 2377 9818
rect 2429 9766 2441 9818
rect 2493 9766 2505 9818
rect 2557 9766 5951 9818
rect 6003 9766 6015 9818
rect 6067 9766 6079 9818
rect 6131 9766 6143 9818
rect 6195 9766 6207 9818
rect 6259 9766 9653 9818
rect 9705 9766 9717 9818
rect 9769 9766 9781 9818
rect 9833 9766 9845 9818
rect 9897 9766 9909 9818
rect 9961 9766 13355 9818
rect 13407 9766 13419 9818
rect 13471 9766 13483 9818
rect 13535 9766 13547 9818
rect 13599 9766 13611 9818
rect 13663 9766 15364 9818
rect 552 9744 15364 9766
rect 5258 9704 5264 9716
rect 4908 9676 5264 9704
rect 4908 9577 4936 9676
rect 5258 9664 5264 9676
rect 5316 9664 5322 9716
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 6733 9707 6791 9713
rect 6733 9704 6745 9707
rect 5868 9676 6745 9704
rect 5868 9664 5874 9676
rect 6733 9673 6745 9676
rect 6779 9673 6791 9707
rect 6733 9667 6791 9673
rect 7558 9664 7564 9716
rect 7616 9664 7622 9716
rect 7742 9664 7748 9716
rect 7800 9664 7806 9716
rect 8478 9664 8484 9716
rect 8536 9664 8542 9716
rect 8570 9664 8576 9716
rect 8628 9664 8634 9716
rect 8662 9664 8668 9716
rect 8720 9704 8726 9716
rect 9309 9707 9367 9713
rect 9309 9704 9321 9707
rect 8720 9676 9321 9704
rect 8720 9664 8726 9676
rect 9309 9673 9321 9676
rect 9355 9673 9367 9707
rect 9309 9667 9367 9673
rect 11238 9664 11244 9716
rect 11296 9704 11302 9716
rect 11333 9707 11391 9713
rect 11333 9704 11345 9707
rect 11296 9676 11345 9704
rect 11296 9664 11302 9676
rect 11333 9673 11345 9676
rect 11379 9673 11391 9707
rect 13170 9704 13176 9716
rect 11333 9667 11391 9673
rect 12728 9676 13176 9704
rect 6270 9596 6276 9648
rect 6328 9596 6334 9648
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 7101 9571 7159 9577
rect 7101 9537 7113 9571
rect 7147 9568 7159 9571
rect 7576 9568 7604 9664
rect 7147 9540 7604 9568
rect 7760 9568 7788 9664
rect 8496 9636 8524 9664
rect 8757 9639 8815 9645
rect 8757 9636 8769 9639
rect 8496 9608 8769 9636
rect 8757 9605 8769 9608
rect 8803 9605 8815 9639
rect 8757 9599 8815 9605
rect 10870 9596 10876 9648
rect 10928 9636 10934 9648
rect 12618 9636 12624 9648
rect 10928 9608 12624 9636
rect 10928 9596 10934 9608
rect 12618 9596 12624 9608
rect 12676 9596 12682 9648
rect 8570 9568 8576 9580
rect 7760 9540 8576 9568
rect 7147 9537 7159 9540
rect 7101 9531 7159 9537
rect 8570 9528 8576 9540
rect 8628 9528 8634 9580
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9568 10747 9571
rect 12066 9568 12072 9580
rect 10735 9540 12072 9568
rect 10735 9537 10747 9540
rect 10689 9531 10747 9537
rect 12066 9528 12072 9540
rect 12124 9528 12130 9580
rect 5166 9509 5172 9512
rect 5160 9500 5172 9509
rect 5127 9472 5172 9500
rect 5160 9463 5172 9472
rect 5166 9460 5172 9463
rect 5224 9460 5230 9512
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 6472 9472 6929 9500
rect 6472 9376 6500 9472
rect 6917 9469 6929 9472
rect 6963 9469 6975 9503
rect 6917 9463 6975 9469
rect 7006 9460 7012 9512
rect 7064 9460 7070 9512
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9500 7251 9503
rect 7282 9500 7288 9512
rect 7239 9472 7288 9500
rect 7239 9469 7251 9472
rect 7193 9463 7251 9469
rect 7282 9460 7288 9472
rect 7340 9460 7346 9512
rect 7374 9460 7380 9512
rect 7432 9460 7438 9512
rect 10134 9460 10140 9512
rect 10192 9500 10198 9512
rect 10422 9503 10480 9509
rect 10422 9500 10434 9503
rect 10192 9472 10434 9500
rect 10192 9460 10198 9472
rect 10422 9469 10434 9472
rect 10468 9469 10480 9503
rect 10422 9463 10480 9469
rect 10778 9460 10784 9512
rect 10836 9460 10842 9512
rect 10870 9460 10876 9512
rect 10928 9500 10934 9512
rect 10965 9503 11023 9509
rect 10965 9500 10977 9503
rect 10928 9472 10977 9500
rect 10928 9460 10934 9472
rect 10965 9469 10977 9472
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 11146 9460 11152 9512
rect 11204 9460 11210 9512
rect 12434 9460 12440 9512
rect 12492 9460 12498 9512
rect 12618 9509 12624 9512
rect 12585 9503 12624 9509
rect 12585 9469 12597 9503
rect 12585 9463 12624 9469
rect 12618 9460 12624 9463
rect 12676 9460 12682 9512
rect 12728 9509 12756 9676
rect 13170 9664 13176 9676
rect 13228 9704 13234 9716
rect 13357 9707 13415 9713
rect 13357 9704 13369 9707
rect 13228 9676 13369 9704
rect 13228 9664 13234 9676
rect 13357 9673 13369 9676
rect 13403 9673 13415 9707
rect 13357 9667 13415 9673
rect 13081 9639 13139 9645
rect 13081 9605 13093 9639
rect 13127 9636 13139 9639
rect 13127 9608 14044 9636
rect 13127 9605 13139 9608
rect 13081 9599 13139 9605
rect 12713 9503 12771 9509
rect 12713 9469 12725 9503
rect 12759 9469 12771 9503
rect 12713 9463 12771 9469
rect 12802 9460 12808 9512
rect 12860 9460 12866 9512
rect 12902 9503 12960 9509
rect 12902 9469 12914 9503
rect 12948 9469 12960 9503
rect 12902 9463 12960 9469
rect 7929 9435 7987 9441
rect 7929 9432 7941 9435
rect 6932 9404 7941 9432
rect 6932 9376 6960 9404
rect 7929 9401 7941 9404
rect 7975 9432 7987 9435
rect 8294 9432 8300 9444
rect 7975 9404 8300 9432
rect 7975 9401 7987 9404
rect 7929 9395 7987 9401
rect 8294 9392 8300 9404
rect 8352 9432 8358 9444
rect 8389 9435 8447 9441
rect 8389 9432 8401 9435
rect 8352 9404 8401 9432
rect 8352 9392 8358 9404
rect 8389 9401 8401 9404
rect 8435 9401 8447 9435
rect 8389 9395 8447 9401
rect 9030 9392 9036 9444
rect 9088 9432 9094 9444
rect 9088 9404 12664 9432
rect 9088 9392 9094 9404
rect 6454 9324 6460 9376
rect 6512 9324 6518 9376
rect 6914 9324 6920 9376
rect 6972 9324 6978 9376
rect 7466 9324 7472 9376
rect 7524 9364 7530 9376
rect 7719 9367 7777 9373
rect 7719 9364 7731 9367
rect 7524 9336 7731 9364
rect 7524 9324 7530 9336
rect 7719 9333 7731 9336
rect 7765 9333 7777 9367
rect 7719 9327 7777 9333
rect 8599 9367 8657 9373
rect 8599 9333 8611 9367
rect 8645 9364 8657 9367
rect 9122 9364 9128 9376
rect 8645 9336 9128 9364
rect 8645 9333 8657 9336
rect 8599 9327 8657 9333
rect 9122 9324 9128 9336
rect 9180 9324 9186 9376
rect 9398 9324 9404 9376
rect 9456 9364 9462 9376
rect 10870 9364 10876 9376
rect 9456 9336 10876 9364
rect 9456 9324 9462 9336
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 10962 9324 10968 9376
rect 11020 9324 11026 9376
rect 12636 9364 12664 9404
rect 12912 9364 12940 9463
rect 13170 9460 13176 9512
rect 13228 9460 13234 9512
rect 13357 9503 13415 9509
rect 13357 9469 13369 9503
rect 13403 9469 13415 9503
rect 13357 9463 13415 9469
rect 13817 9503 13875 9509
rect 13817 9469 13829 9503
rect 13863 9469 13875 9503
rect 13817 9463 13875 9469
rect 13372 9432 13400 9463
rect 13188 9404 13400 9432
rect 13832 9432 13860 9463
rect 13906 9460 13912 9512
rect 13964 9460 13970 9512
rect 14016 9509 14044 9608
rect 14001 9503 14059 9509
rect 14001 9469 14013 9503
rect 14047 9469 14059 9503
rect 14001 9463 14059 9469
rect 14090 9460 14096 9512
rect 14148 9500 14154 9512
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 14148 9472 14197 9500
rect 14148 9460 14154 9472
rect 14185 9469 14197 9472
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 14918 9460 14924 9512
rect 14976 9460 14982 9512
rect 14936 9432 14964 9460
rect 13832 9404 14964 9432
rect 13188 9376 13216 9404
rect 12636 9336 12940 9364
rect 13170 9324 13176 9376
rect 13228 9324 13234 9376
rect 13541 9367 13599 9373
rect 13541 9333 13553 9367
rect 13587 9364 13599 9367
rect 13630 9364 13636 9376
rect 13587 9336 13636 9364
rect 13587 9333 13599 9336
rect 13541 9327 13599 9333
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 552 9274 15520 9296
rect 552 9222 4100 9274
rect 4152 9222 4164 9274
rect 4216 9222 4228 9274
rect 4280 9222 4292 9274
rect 4344 9222 4356 9274
rect 4408 9222 7802 9274
rect 7854 9222 7866 9274
rect 7918 9222 7930 9274
rect 7982 9222 7994 9274
rect 8046 9222 8058 9274
rect 8110 9222 11504 9274
rect 11556 9222 11568 9274
rect 11620 9222 11632 9274
rect 11684 9222 11696 9274
rect 11748 9222 11760 9274
rect 11812 9222 15206 9274
rect 15258 9222 15270 9274
rect 15322 9222 15334 9274
rect 15386 9222 15398 9274
rect 15450 9222 15462 9274
rect 15514 9222 15520 9274
rect 552 9200 15520 9222
rect 5258 9120 5264 9172
rect 5316 9120 5322 9172
rect 5442 9120 5448 9172
rect 5500 9120 5506 9172
rect 6825 9163 6883 9169
rect 6825 9129 6837 9163
rect 6871 9160 6883 9163
rect 7098 9160 7104 9172
rect 6871 9132 7104 9160
rect 6871 9129 6883 9132
rect 6825 9123 6883 9129
rect 5276 9092 5304 9120
rect 5460 9092 5488 9120
rect 6454 9092 6460 9104
rect 5184 9064 5304 9092
rect 5368 9064 5488 9092
rect 6196 9064 6460 9092
rect 5184 9033 5212 9064
rect 4913 9027 4971 9033
rect 4913 8993 4925 9027
rect 4959 9024 4971 9027
rect 5169 9027 5227 9033
rect 4959 8996 5120 9024
rect 4959 8993 4971 8996
rect 4913 8987 4971 8993
rect 5092 8956 5120 8996
rect 5169 8993 5181 9027
rect 5215 8993 5227 9027
rect 5169 8987 5227 8993
rect 5261 9027 5319 9033
rect 5261 8993 5273 9027
rect 5307 9024 5319 9027
rect 5368 9024 5396 9064
rect 6196 9033 6224 9064
rect 6454 9052 6460 9064
rect 6512 9052 6518 9104
rect 6840 9092 6868 9123
rect 7098 9120 7104 9132
rect 7156 9120 7162 9172
rect 7653 9163 7711 9169
rect 7653 9129 7665 9163
rect 7699 9160 7711 9163
rect 8202 9160 8208 9172
rect 7699 9132 8208 9160
rect 7699 9129 7711 9132
rect 7653 9123 7711 9129
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 11514 9160 11520 9172
rect 10244 9132 11520 9160
rect 6656 9064 6868 9092
rect 5307 8996 5396 9024
rect 5445 9027 5503 9033
rect 5307 8993 5319 8996
rect 5261 8987 5319 8993
rect 5445 8993 5457 9027
rect 5491 9024 5503 9027
rect 6181 9027 6239 9033
rect 5491 8996 5580 9024
rect 5491 8993 5503 8996
rect 5445 8987 5503 8993
rect 5353 8959 5411 8965
rect 5353 8956 5365 8959
rect 5092 8928 5365 8956
rect 5353 8925 5365 8928
rect 5399 8925 5411 8959
rect 5552 8956 5580 8996
rect 6181 8993 6193 9027
rect 6227 8993 6239 9027
rect 6181 8987 6239 8993
rect 6365 9027 6423 9033
rect 6365 8993 6377 9027
rect 6411 9024 6423 9027
rect 6546 9024 6552 9036
rect 6411 8996 6552 9024
rect 6411 8993 6423 8996
rect 6365 8987 6423 8993
rect 6546 8984 6552 8996
rect 6604 8984 6610 9036
rect 6656 9033 6684 9064
rect 6914 9052 6920 9104
rect 6972 9052 6978 9104
rect 10244 9101 10272 9132
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 11609 9163 11667 9169
rect 11609 9129 11621 9163
rect 11655 9129 11667 9163
rect 11609 9123 11667 9129
rect 7285 9095 7343 9101
rect 7285 9061 7297 9095
rect 7331 9092 7343 9095
rect 10229 9095 10287 9101
rect 7331 9064 8616 9092
rect 7331 9061 7343 9064
rect 7285 9055 7343 9061
rect 6641 9027 6699 9033
rect 6641 8993 6653 9027
rect 6687 8993 6699 9027
rect 6641 8987 6699 8993
rect 6733 9027 6791 9033
rect 6733 8993 6745 9027
rect 6779 8993 6791 9027
rect 6932 9024 6960 9052
rect 8588 9036 8616 9064
rect 10229 9061 10241 9095
rect 10275 9061 10287 9095
rect 10229 9055 10287 9061
rect 7101 9027 7159 9033
rect 7101 9024 7113 9027
rect 6932 8996 7113 9024
rect 6733 8987 6791 8993
rect 7101 8993 7113 8996
rect 7147 8993 7159 9027
rect 7101 8987 7159 8993
rect 7377 9027 7435 9033
rect 7377 8993 7389 9027
rect 7423 9024 7435 9027
rect 7466 9024 7472 9036
rect 7423 8996 7472 9024
rect 7423 8993 7435 8996
rect 7377 8987 7435 8993
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5552 8928 6009 8956
rect 5353 8919 5411 8925
rect 5997 8925 6009 8928
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 6270 8848 6276 8900
rect 6328 8848 6334 8900
rect 6472 8888 6500 8919
rect 6638 8888 6644 8900
rect 6472 8860 6644 8888
rect 6638 8848 6644 8860
rect 6696 8848 6702 8900
rect 6748 8832 6776 8987
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 7558 8984 7564 9036
rect 7616 8984 7622 9036
rect 8570 8984 8576 9036
rect 8628 8984 8634 9036
rect 10962 8984 10968 9036
rect 11020 9024 11026 9036
rect 11240 9027 11298 9033
rect 11240 9024 11252 9027
rect 11020 8996 11252 9024
rect 11020 8984 11026 8996
rect 11240 8993 11252 8996
rect 11286 8993 11298 9027
rect 11240 8987 11298 8993
rect 11333 9027 11391 9033
rect 11333 8993 11345 9027
rect 11379 9024 11391 9027
rect 11624 9024 11652 9123
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 15010 9160 15016 9172
rect 11756 9132 15016 9160
rect 11756 9120 11762 9132
rect 15010 9120 15016 9132
rect 15068 9120 15074 9172
rect 12158 9092 12164 9104
rect 11900 9064 12164 9092
rect 11900 9033 11928 9064
rect 12158 9052 12164 9064
rect 12216 9052 12222 9104
rect 12618 9052 12624 9104
rect 12676 9092 12682 9104
rect 12713 9095 12771 9101
rect 12713 9092 12725 9095
rect 12676 9064 12725 9092
rect 12676 9052 12682 9064
rect 12713 9061 12725 9064
rect 12759 9061 12771 9095
rect 12713 9055 12771 9061
rect 13262 9052 13268 9104
rect 13320 9092 13326 9104
rect 13320 9064 13400 9092
rect 13320 9052 13326 9064
rect 11379 8996 11652 9024
rect 11885 9027 11943 9033
rect 11379 8993 11391 8996
rect 11333 8987 11391 8993
rect 11885 8993 11897 9027
rect 11931 8993 11943 9027
rect 11885 8987 11943 8993
rect 11974 8984 11980 9036
rect 12032 9024 12038 9036
rect 12345 9027 12403 9033
rect 12345 9024 12357 9027
rect 12032 8996 12357 9024
rect 12032 8984 12038 8996
rect 12345 8993 12357 8996
rect 12391 8993 12403 9027
rect 12345 8987 12403 8993
rect 12526 8984 12532 9036
rect 12584 8984 12590 9036
rect 13372 9033 13400 9064
rect 13357 9027 13415 9033
rect 13357 8993 13369 9027
rect 13403 8993 13415 9027
rect 13357 8987 13415 8993
rect 13630 8984 13636 9036
rect 13688 8984 13694 9036
rect 13906 8984 13912 9036
rect 13964 8984 13970 9036
rect 7006 8916 7012 8968
rect 7064 8916 7070 8968
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 11057 8959 11115 8965
rect 11057 8956 11069 8959
rect 10744 8928 11069 8956
rect 10744 8916 10750 8928
rect 11057 8925 11069 8928
rect 11103 8925 11115 8959
rect 11057 8919 11115 8925
rect 11146 8916 11152 8968
rect 11204 8916 11210 8968
rect 11514 8916 11520 8968
rect 11572 8916 11578 8968
rect 11698 8916 11704 8968
rect 11756 8956 11762 8968
rect 13924 8956 13952 8984
rect 11756 8928 13952 8956
rect 11756 8916 11762 8928
rect 7024 8888 7052 8916
rect 7101 8891 7159 8897
rect 7101 8888 7113 8891
rect 7024 8860 7113 8888
rect 7101 8857 7113 8860
rect 7147 8857 7159 8891
rect 11164 8888 11192 8916
rect 11532 8888 11560 8916
rect 11164 8860 11560 8888
rect 7101 8851 7159 8857
rect 3789 8823 3847 8829
rect 3789 8789 3801 8823
rect 3835 8820 3847 8823
rect 5810 8820 5816 8832
rect 3835 8792 5816 8820
rect 3835 8789 3847 8792
rect 3789 8783 3847 8789
rect 5810 8780 5816 8792
rect 5868 8820 5874 8832
rect 6730 8820 6736 8832
rect 5868 8792 6736 8820
rect 5868 8780 5874 8792
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 8938 8780 8944 8832
rect 8996 8780 9002 8832
rect 11517 8823 11575 8829
rect 11517 8789 11529 8823
rect 11563 8820 11575 8823
rect 11698 8820 11704 8832
rect 11563 8792 11704 8820
rect 11563 8789 11575 8792
rect 11517 8783 11575 8789
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 11790 8780 11796 8832
rect 11848 8780 11854 8832
rect 14921 8823 14979 8829
rect 14921 8789 14933 8823
rect 14967 8820 14979 8823
rect 15010 8820 15016 8832
rect 14967 8792 15016 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15010 8780 15016 8792
rect 15068 8780 15074 8832
rect 552 8730 15364 8752
rect 552 8678 2249 8730
rect 2301 8678 2313 8730
rect 2365 8678 2377 8730
rect 2429 8678 2441 8730
rect 2493 8678 2505 8730
rect 2557 8678 5951 8730
rect 6003 8678 6015 8730
rect 6067 8678 6079 8730
rect 6131 8678 6143 8730
rect 6195 8678 6207 8730
rect 6259 8678 9653 8730
rect 9705 8678 9717 8730
rect 9769 8678 9781 8730
rect 9833 8678 9845 8730
rect 9897 8678 9909 8730
rect 9961 8678 13355 8730
rect 13407 8678 13419 8730
rect 13471 8678 13483 8730
rect 13535 8678 13547 8730
rect 13599 8678 13611 8730
rect 13663 8678 15364 8730
rect 552 8656 15364 8678
rect 6181 8619 6239 8625
rect 6181 8585 6193 8619
rect 6227 8616 6239 8619
rect 6270 8616 6276 8628
rect 6227 8588 6276 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6546 8576 6552 8628
rect 6604 8616 6610 8628
rect 7466 8616 7472 8628
rect 6604 8588 7472 8616
rect 6604 8576 6610 8588
rect 7466 8576 7472 8588
rect 7524 8576 7530 8628
rect 7576 8588 10916 8616
rect 6638 8508 6644 8560
rect 6696 8548 6702 8560
rect 7282 8548 7288 8560
rect 6696 8520 7288 8548
rect 6696 8508 6702 8520
rect 7282 8508 7288 8520
rect 7340 8548 7346 8560
rect 7576 8548 7604 8588
rect 10888 8560 10916 8588
rect 11790 8576 11796 8628
rect 11848 8576 11854 8628
rect 11974 8576 11980 8628
rect 12032 8576 12038 8628
rect 12161 8619 12219 8625
rect 12161 8585 12173 8619
rect 12207 8616 12219 8619
rect 12802 8616 12808 8628
rect 12207 8588 12808 8616
rect 12207 8585 12219 8588
rect 12161 8579 12219 8585
rect 7340 8520 7604 8548
rect 9401 8551 9459 8557
rect 7340 8508 7346 8520
rect 9401 8517 9413 8551
rect 9447 8517 9459 8551
rect 9401 8511 9459 8517
rect 7745 8483 7803 8489
rect 5828 8452 6224 8480
rect 5828 8424 5856 8452
rect 4522 8372 4528 8424
rect 4580 8372 4586 8424
rect 5810 8372 5816 8424
rect 5868 8372 5874 8424
rect 6196 8421 6224 8452
rect 7745 8449 7757 8483
rect 7791 8480 7803 8483
rect 8662 8480 8668 8492
rect 7791 8452 8668 8480
rect 7791 8449 7803 8452
rect 7745 8443 7803 8449
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 9416 8480 9444 8511
rect 10870 8508 10876 8560
rect 10928 8548 10934 8560
rect 11422 8548 11428 8560
rect 10928 8520 11428 8548
rect 10928 8508 10934 8520
rect 11422 8508 11428 8520
rect 11480 8508 11486 8560
rect 12176 8480 12204 8579
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 13170 8576 13176 8628
rect 13228 8616 13234 8628
rect 13265 8619 13323 8625
rect 13265 8616 13277 8619
rect 13228 8588 13277 8616
rect 13228 8576 13234 8588
rect 13265 8585 13277 8588
rect 13311 8585 13323 8619
rect 13265 8579 13323 8585
rect 8772 8452 9444 8480
rect 5905 8415 5963 8421
rect 5905 8381 5917 8415
rect 5951 8381 5963 8415
rect 5905 8375 5963 8381
rect 6181 8415 6239 8421
rect 6181 8381 6193 8415
rect 6227 8381 6239 8415
rect 6181 8375 6239 8381
rect 5920 8288 5948 8375
rect 6362 8372 6368 8424
rect 6420 8412 6426 8424
rect 7101 8415 7159 8421
rect 7101 8412 7113 8415
rect 6420 8384 7113 8412
rect 6420 8372 6426 8384
rect 7101 8381 7113 8384
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 7116 8344 7144 8375
rect 7190 8372 7196 8424
rect 7248 8412 7254 8424
rect 7285 8415 7343 8421
rect 7285 8412 7297 8415
rect 7248 8384 7297 8412
rect 7248 8372 7254 8384
rect 7285 8381 7297 8384
rect 7331 8412 7343 8415
rect 7377 8415 7435 8421
rect 7377 8412 7389 8415
rect 7331 8384 7389 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 7377 8381 7389 8384
rect 7423 8381 7435 8415
rect 7377 8375 7435 8381
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8381 7619 8415
rect 7561 8375 7619 8381
rect 7576 8344 7604 8375
rect 8294 8372 8300 8424
rect 8352 8412 8358 8424
rect 8570 8421 8576 8424
rect 8389 8415 8447 8421
rect 8389 8412 8401 8415
rect 8352 8384 8401 8412
rect 8352 8372 8358 8384
rect 8389 8381 8401 8384
rect 8435 8381 8447 8415
rect 8389 8375 8447 8381
rect 8547 8415 8576 8421
rect 8547 8381 8559 8415
rect 8628 8412 8634 8424
rect 8772 8412 8800 8452
rect 8628 8384 8800 8412
rect 8849 8415 8907 8421
rect 8547 8375 8576 8381
rect 8570 8372 8576 8375
rect 8628 8372 8634 8384
rect 8849 8381 8861 8415
rect 8895 8381 8907 8415
rect 8849 8375 8907 8381
rect 7116 8316 7604 8344
rect 7837 8347 7895 8353
rect 7837 8313 7849 8347
rect 7883 8313 7895 8347
rect 7837 8307 7895 8313
rect 8021 8347 8079 8353
rect 8021 8313 8033 8347
rect 8067 8344 8079 8347
rect 8588 8344 8616 8372
rect 8067 8316 8616 8344
rect 8067 8313 8079 8316
rect 8021 8307 8079 8313
rect 5169 8279 5227 8285
rect 5169 8245 5181 8279
rect 5215 8276 5227 8279
rect 5350 8276 5356 8288
rect 5215 8248 5356 8276
rect 5215 8245 5227 8248
rect 5169 8239 5227 8245
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 5902 8236 5908 8288
rect 5960 8236 5966 8288
rect 5997 8279 6055 8285
rect 5997 8245 6009 8279
rect 6043 8276 6055 8279
rect 6086 8276 6092 8288
rect 6043 8248 6092 8276
rect 6043 8245 6055 8248
rect 5997 8239 6055 8245
rect 6086 8236 6092 8248
rect 6144 8236 6150 8288
rect 7285 8279 7343 8285
rect 7285 8245 7297 8279
rect 7331 8276 7343 8279
rect 7374 8276 7380 8288
rect 7331 8248 7380 8276
rect 7331 8245 7343 8248
rect 7285 8239 7343 8245
rect 7374 8236 7380 8248
rect 7432 8236 7438 8288
rect 7466 8236 7472 8288
rect 7524 8276 7530 8288
rect 7852 8276 7880 8307
rect 8662 8304 8668 8356
rect 8720 8304 8726 8356
rect 8757 8347 8815 8353
rect 8757 8313 8769 8347
rect 8803 8313 8815 8347
rect 8864 8344 8892 8375
rect 9122 8372 9128 8424
rect 9180 8372 9186 8424
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8412 9367 8415
rect 9416 8412 9444 8452
rect 11624 8452 12204 8480
rect 9355 8384 9444 8412
rect 9355 8381 9367 8384
rect 9309 8375 9367 8381
rect 10778 8372 10784 8424
rect 10836 8372 10842 8424
rect 11624 8421 11652 8452
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 12713 8483 12771 8489
rect 12713 8480 12725 8483
rect 12584 8452 12725 8480
rect 12584 8440 12590 8452
rect 12713 8449 12725 8452
rect 12759 8480 12771 8483
rect 15010 8480 15016 8492
rect 12759 8452 15016 8480
rect 12759 8449 12771 8452
rect 12713 8443 12771 8449
rect 15010 8440 15016 8452
rect 15068 8440 15074 8492
rect 11517 8415 11575 8421
rect 11517 8381 11529 8415
rect 11563 8381 11575 8415
rect 11517 8375 11575 8381
rect 11609 8415 11667 8421
rect 11609 8381 11621 8415
rect 11655 8381 11667 8415
rect 11609 8375 11667 8381
rect 9217 8347 9275 8353
rect 9217 8344 9229 8347
rect 8864 8316 9229 8344
rect 8757 8307 8815 8313
rect 9217 8313 9229 8316
rect 9263 8313 9275 8347
rect 9217 8307 9275 8313
rect 7524 8248 7880 8276
rect 8205 8279 8263 8285
rect 7524 8236 7530 8248
rect 8205 8245 8217 8279
rect 8251 8276 8263 8279
rect 8772 8276 8800 8307
rect 9674 8304 9680 8356
rect 9732 8344 9738 8356
rect 10514 8347 10572 8353
rect 10514 8344 10526 8347
rect 9732 8316 10526 8344
rect 9732 8304 9738 8316
rect 10514 8313 10526 8316
rect 10560 8313 10572 8347
rect 10514 8307 10572 8313
rect 8251 8248 8800 8276
rect 8251 8245 8263 8248
rect 8205 8239 8263 8245
rect 9030 8236 9036 8288
rect 9088 8236 9094 8288
rect 11422 8236 11428 8288
rect 11480 8276 11486 8288
rect 11532 8276 11560 8375
rect 11698 8372 11704 8424
rect 11756 8412 11762 8424
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 11756 8384 13737 8412
rect 11756 8372 11762 8384
rect 13725 8381 13737 8384
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 13906 8372 13912 8424
rect 13964 8412 13970 8424
rect 14001 8415 14059 8421
rect 14001 8412 14013 8415
rect 13964 8384 14013 8412
rect 13964 8372 13970 8384
rect 14001 8381 14013 8384
rect 14047 8381 14059 8415
rect 14001 8375 14059 8381
rect 14185 8415 14243 8421
rect 14185 8381 14197 8415
rect 14231 8412 14243 8415
rect 14369 8415 14427 8421
rect 14369 8412 14381 8415
rect 14231 8384 14381 8412
rect 14231 8381 14243 8384
rect 14185 8375 14243 8381
rect 14369 8381 14381 8384
rect 14415 8381 14427 8415
rect 14369 8375 14427 8381
rect 14921 8415 14979 8421
rect 14921 8381 14933 8415
rect 14967 8412 14979 8415
rect 15102 8412 15108 8424
rect 14967 8384 15108 8412
rect 14967 8381 14979 8384
rect 14921 8375 14979 8381
rect 11793 8347 11851 8353
rect 11793 8313 11805 8347
rect 11839 8344 11851 8347
rect 12345 8347 12403 8353
rect 12345 8344 12357 8347
rect 11839 8316 12357 8344
rect 11839 8313 11851 8316
rect 11793 8307 11851 8313
rect 12345 8313 12357 8316
rect 12391 8344 12403 8347
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 12391 8316 12909 8344
rect 12391 8313 12403 8316
rect 12345 8307 12403 8313
rect 12897 8313 12909 8316
rect 12943 8344 12955 8347
rect 14936 8344 14964 8375
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 12943 8316 14964 8344
rect 12943 8313 12955 8316
rect 12897 8307 12955 8313
rect 12145 8279 12203 8285
rect 12145 8276 12157 8279
rect 11480 8248 12157 8276
rect 11480 8236 11486 8248
rect 12145 8245 12157 8248
rect 12191 8276 12203 8279
rect 12618 8276 12624 8288
rect 12191 8248 12624 8276
rect 12191 8245 12203 8248
rect 12145 8239 12203 8245
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 12802 8236 12808 8288
rect 12860 8276 12866 8288
rect 12989 8279 13047 8285
rect 12989 8276 13001 8279
rect 12860 8248 13001 8276
rect 12860 8236 12866 8248
rect 12989 8245 13001 8248
rect 13035 8245 13047 8279
rect 12989 8239 13047 8245
rect 13081 8279 13139 8285
rect 13081 8245 13093 8279
rect 13127 8276 13139 8279
rect 13170 8276 13176 8288
rect 13127 8248 13176 8276
rect 13127 8245 13139 8248
rect 13081 8239 13139 8245
rect 13170 8236 13176 8248
rect 13228 8236 13234 8288
rect 13541 8279 13599 8285
rect 13541 8245 13553 8279
rect 13587 8276 13599 8279
rect 13630 8276 13636 8288
rect 13587 8248 13636 8276
rect 13587 8245 13599 8248
rect 13541 8239 13599 8245
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 552 8186 15520 8208
rect 552 8134 4100 8186
rect 4152 8134 4164 8186
rect 4216 8134 4228 8186
rect 4280 8134 4292 8186
rect 4344 8134 4356 8186
rect 4408 8134 7802 8186
rect 7854 8134 7866 8186
rect 7918 8134 7930 8186
rect 7982 8134 7994 8186
rect 8046 8134 8058 8186
rect 8110 8134 11504 8186
rect 11556 8134 11568 8186
rect 11620 8134 11632 8186
rect 11684 8134 11696 8186
rect 11748 8134 11760 8186
rect 11812 8134 15206 8186
rect 15258 8134 15270 8186
rect 15322 8134 15334 8186
rect 15386 8134 15398 8186
rect 15450 8134 15462 8186
rect 15514 8134 15520 8186
rect 552 8112 15520 8134
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 4522 8072 4528 8084
rect 3559 8044 4528 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 4522 8032 4528 8044
rect 4580 8072 4586 8084
rect 6917 8075 6975 8081
rect 4580 8044 5856 8072
rect 4580 8032 4586 8044
rect 4648 8007 4706 8013
rect 4648 7973 4660 8007
rect 4694 8004 4706 8007
rect 5169 8007 5227 8013
rect 4694 7976 5120 8004
rect 4694 7973 4706 7976
rect 4648 7967 4706 7973
rect 4982 7896 4988 7948
rect 5040 7896 5046 7948
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7837 4951 7871
rect 5092 7868 5120 7976
rect 5169 7973 5181 8007
rect 5215 8004 5227 8007
rect 5445 8007 5503 8013
rect 5445 8004 5457 8007
rect 5215 7976 5457 8004
rect 5215 7973 5227 7976
rect 5169 7967 5227 7973
rect 5445 7973 5457 7976
rect 5491 7973 5503 8007
rect 5445 7967 5503 7973
rect 5261 7939 5319 7945
rect 5261 7905 5273 7939
rect 5307 7905 5319 7939
rect 5261 7899 5319 7905
rect 4893 7831 4951 7837
rect 5000 7840 5120 7868
rect 5276 7868 5304 7899
rect 5350 7896 5356 7948
rect 5408 7896 5414 7948
rect 5537 7939 5595 7945
rect 5537 7905 5549 7939
rect 5583 7936 5595 7939
rect 5718 7936 5724 7948
rect 5583 7908 5724 7936
rect 5583 7905 5595 7908
rect 5537 7899 5595 7905
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 5828 7936 5856 8044
rect 6917 8041 6929 8075
rect 6963 8072 6975 8075
rect 7558 8072 7564 8084
rect 6963 8044 7564 8072
rect 6963 8041 6975 8044
rect 6917 8035 6975 8041
rect 5902 7964 5908 8016
rect 5960 8004 5966 8016
rect 5960 7976 6500 8004
rect 5960 7964 5966 7976
rect 6012 7945 6040 7976
rect 6472 7948 6500 7976
rect 6730 7964 6736 8016
rect 6788 7964 6794 8016
rect 5997 7939 6055 7945
rect 5828 7908 5948 7936
rect 5813 7871 5871 7877
rect 5813 7868 5825 7871
rect 5276 7840 5825 7868
rect 4522 7692 4528 7744
rect 4580 7732 4586 7744
rect 4908 7732 4936 7831
rect 5000 7809 5028 7840
rect 5813 7837 5825 7840
rect 5859 7837 5871 7871
rect 5920 7868 5948 7908
rect 5997 7905 6009 7939
rect 6043 7905 6055 7939
rect 5997 7899 6055 7905
rect 6086 7896 6092 7948
rect 6144 7936 6150 7948
rect 6273 7939 6331 7945
rect 6144 7908 6224 7936
rect 6144 7896 6150 7908
rect 6196 7868 6224 7908
rect 6273 7905 6285 7939
rect 6319 7905 6331 7939
rect 6273 7899 6331 7905
rect 5920 7840 6224 7868
rect 6288 7868 6316 7899
rect 6362 7896 6368 7948
rect 6420 7896 6426 7948
rect 6454 7896 6460 7948
rect 6512 7896 6518 7948
rect 6641 7939 6699 7945
rect 6641 7905 6653 7939
rect 6687 7936 6699 7939
rect 6932 7936 6960 8035
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 8386 8032 8392 8084
rect 8444 8032 8450 8084
rect 9030 8032 9036 8084
rect 9088 8032 9094 8084
rect 9674 8032 9680 8084
rect 9732 8032 9738 8084
rect 11532 8044 12296 8072
rect 7006 7964 7012 8016
rect 7064 8004 7070 8016
rect 8404 8004 8432 8032
rect 7064 7976 8432 8004
rect 7064 7964 7070 7976
rect 6687 7908 6960 7936
rect 7101 7939 7159 7945
rect 6687 7905 6699 7908
rect 6641 7899 6699 7905
rect 7101 7905 7113 7939
rect 7147 7936 7159 7939
rect 8846 7936 8852 7948
rect 7147 7908 8852 7936
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 6549 7871 6607 7877
rect 6549 7868 6561 7871
rect 6288 7840 6561 7868
rect 5813 7831 5871 7837
rect 4985 7803 5043 7809
rect 4985 7769 4997 7803
rect 5031 7769 5043 7803
rect 4985 7763 5043 7769
rect 5718 7760 5724 7812
rect 5776 7760 5782 7812
rect 6196 7800 6224 7840
rect 6549 7837 6561 7840
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 6656 7800 6684 7899
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 9048 7936 9076 8032
rect 11238 8004 11244 8016
rect 10428 7976 11244 8004
rect 10428 7948 10456 7976
rect 11238 7964 11244 7976
rect 11296 8004 11302 8016
rect 11532 8004 11560 8044
rect 11296 7976 11560 8004
rect 11296 7964 11302 7976
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 9048 7908 9229 7936
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 9217 7899 9275 7905
rect 9401 7939 9459 7945
rect 9401 7905 9413 7939
rect 9447 7936 9459 7939
rect 9493 7939 9551 7945
rect 9493 7936 9505 7939
rect 9447 7908 9505 7936
rect 9447 7905 9459 7908
rect 9401 7899 9459 7905
rect 9493 7905 9505 7908
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 10410 7896 10416 7948
rect 10468 7896 10474 7948
rect 11422 7896 11428 7948
rect 11480 7896 11486 7948
rect 11532 7936 11560 7976
rect 11609 8007 11667 8013
rect 11609 7973 11621 8007
rect 11655 8004 11667 8007
rect 12161 8007 12219 8013
rect 12161 8004 12173 8007
rect 11655 7976 12173 8004
rect 11655 7973 11667 7976
rect 11609 7967 11667 7973
rect 12161 7973 12173 7976
rect 12207 7973 12219 8007
rect 12161 7967 12219 7973
rect 12268 7948 12296 8044
rect 11701 7939 11759 7945
rect 11701 7936 11713 7939
rect 11532 7908 11713 7936
rect 11701 7905 11713 7908
rect 11747 7905 11759 7939
rect 11701 7899 11759 7905
rect 11793 7939 11851 7945
rect 11793 7905 11805 7939
rect 11839 7905 11851 7939
rect 11793 7899 11851 7905
rect 12069 7939 12127 7945
rect 12069 7905 12081 7939
rect 12115 7905 12127 7939
rect 12069 7899 12127 7905
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9306 7868 9312 7880
rect 9088 7840 9312 7868
rect 9088 7828 9094 7840
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 11330 7828 11336 7880
rect 11388 7868 11394 7880
rect 11808 7868 11836 7899
rect 11388 7840 11836 7868
rect 12084 7868 12112 7899
rect 12250 7896 12256 7948
rect 12308 7896 12314 7948
rect 12802 7896 12808 7948
rect 12860 7896 12866 7948
rect 13630 7896 13636 7948
rect 13688 7896 13694 7948
rect 12820 7868 12848 7896
rect 12084 7840 12848 7868
rect 11388 7828 11394 7840
rect 13262 7828 13268 7880
rect 13320 7868 13326 7880
rect 13357 7871 13415 7877
rect 13357 7868 13369 7871
rect 13320 7840 13369 7868
rect 13320 7828 13326 7840
rect 13357 7837 13369 7840
rect 13403 7837 13415 7871
rect 13357 7831 13415 7837
rect 9398 7800 9404 7812
rect 6196 7772 6684 7800
rect 7208 7772 9404 7800
rect 4580 7704 4936 7732
rect 5736 7732 5764 7760
rect 7208 7732 7236 7772
rect 9398 7760 9404 7772
rect 9456 7760 9462 7812
rect 5736 7704 7236 7732
rect 4580 7692 4586 7704
rect 7282 7692 7288 7744
rect 7340 7692 7346 7744
rect 11977 7735 12035 7741
rect 11977 7701 11989 7735
rect 12023 7732 12035 7735
rect 12158 7732 12164 7744
rect 12023 7704 12164 7732
rect 12023 7701 12035 7704
rect 11977 7695 12035 7701
rect 12158 7692 12164 7704
rect 12216 7692 12222 7744
rect 14921 7735 14979 7741
rect 14921 7701 14933 7735
rect 14967 7732 14979 7735
rect 15102 7732 15108 7744
rect 14967 7704 15108 7732
rect 14967 7701 14979 7704
rect 14921 7695 14979 7701
rect 15102 7692 15108 7704
rect 15160 7692 15166 7744
rect 552 7642 15364 7664
rect 552 7590 2249 7642
rect 2301 7590 2313 7642
rect 2365 7590 2377 7642
rect 2429 7590 2441 7642
rect 2493 7590 2505 7642
rect 2557 7590 5951 7642
rect 6003 7590 6015 7642
rect 6067 7590 6079 7642
rect 6131 7590 6143 7642
rect 6195 7590 6207 7642
rect 6259 7590 9653 7642
rect 9705 7590 9717 7642
rect 9769 7590 9781 7642
rect 9833 7590 9845 7642
rect 9897 7590 9909 7642
rect 9961 7590 13355 7642
rect 13407 7590 13419 7642
rect 13471 7590 13483 7642
rect 13535 7590 13547 7642
rect 13599 7590 13611 7642
rect 13663 7590 15364 7642
rect 552 7568 15364 7590
rect 7929 7531 7987 7537
rect 7929 7497 7941 7531
rect 7975 7528 7987 7531
rect 9122 7528 9128 7540
rect 7975 7500 9128 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 12437 7463 12495 7469
rect 12437 7429 12449 7463
rect 12483 7460 12495 7463
rect 13078 7460 13084 7472
rect 12483 7432 13084 7460
rect 12483 7429 12495 7432
rect 12437 7423 12495 7429
rect 13078 7420 13084 7432
rect 13136 7420 13142 7472
rect 7282 7352 7288 7404
rect 7340 7392 7346 7404
rect 7340 7364 7788 7392
rect 7340 7352 7346 7364
rect 7650 7284 7656 7336
rect 7708 7284 7714 7336
rect 7760 7333 7788 7364
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 9033 7395 9091 7401
rect 9033 7392 9045 7395
rect 8352 7364 9045 7392
rect 8352 7352 8358 7364
rect 9033 7361 9045 7364
rect 9079 7392 9091 7395
rect 10410 7392 10416 7404
rect 9079 7364 10416 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 10502 7352 10508 7404
rect 10560 7392 10566 7404
rect 10560 7364 12204 7392
rect 10560 7352 10566 7364
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7293 7803 7327
rect 7745 7287 7803 7293
rect 8202 7284 8208 7336
rect 8260 7324 8266 7336
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 8260 7296 8585 7324
rect 8260 7284 8266 7296
rect 8573 7293 8585 7296
rect 8619 7293 8631 7327
rect 8573 7287 8631 7293
rect 8846 7284 8852 7336
rect 8904 7333 8910 7336
rect 8904 7327 8933 7333
rect 8921 7293 8933 7327
rect 8904 7287 8933 7293
rect 11977 7327 12035 7333
rect 11977 7293 11989 7327
rect 12023 7324 12035 7327
rect 12066 7324 12072 7336
rect 12023 7296 12072 7324
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 8904 7284 8910 7287
rect 12066 7284 12072 7296
rect 12124 7284 12130 7336
rect 12176 7333 12204 7364
rect 12618 7352 12624 7404
rect 12676 7392 12682 7404
rect 12676 7364 13216 7392
rect 12676 7352 12682 7364
rect 12161 7327 12219 7333
rect 12161 7293 12173 7327
rect 12207 7293 12219 7327
rect 12161 7287 12219 7293
rect 12250 7284 12256 7336
rect 12308 7284 12314 7336
rect 12535 7327 12593 7333
rect 12535 7293 12547 7327
rect 12581 7324 12593 7327
rect 12636 7324 12664 7352
rect 13188 7336 13216 7364
rect 12581 7296 12664 7324
rect 12713 7327 12771 7333
rect 12581 7293 12593 7296
rect 12535 7287 12593 7293
rect 12713 7293 12725 7327
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 8294 7216 8300 7268
rect 8352 7256 8358 7268
rect 8665 7259 8723 7265
rect 8665 7256 8677 7259
rect 8352 7228 8677 7256
rect 8352 7216 8358 7228
rect 8665 7225 8677 7228
rect 8711 7225 8723 7259
rect 8665 7219 8723 7225
rect 8754 7216 8760 7268
rect 8812 7256 8818 7268
rect 9217 7259 9275 7265
rect 9217 7256 9229 7259
rect 8812 7228 9229 7256
rect 8812 7216 8818 7228
rect 9217 7225 9229 7228
rect 9263 7225 9275 7259
rect 9217 7219 9275 7225
rect 9585 7259 9643 7265
rect 9585 7225 9597 7259
rect 9631 7256 9643 7259
rect 10226 7256 10232 7268
rect 9631 7228 10232 7256
rect 9631 7225 9643 7228
rect 9585 7219 9643 7225
rect 10226 7216 10232 7228
rect 10284 7216 10290 7268
rect 6270 7148 6276 7200
rect 6328 7188 6334 7200
rect 6638 7188 6644 7200
rect 6328 7160 6644 7188
rect 6328 7148 6334 7160
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 8386 7148 8392 7200
rect 8444 7148 8450 7200
rect 10502 7148 10508 7200
rect 10560 7188 10566 7200
rect 11333 7191 11391 7197
rect 11333 7188 11345 7191
rect 10560 7160 11345 7188
rect 10560 7148 10566 7160
rect 11333 7157 11345 7160
rect 11379 7157 11391 7191
rect 12268 7188 12296 7284
rect 12437 7259 12495 7265
rect 12437 7225 12449 7259
rect 12483 7256 12495 7259
rect 12618 7256 12624 7268
rect 12483 7228 12624 7256
rect 12483 7225 12495 7228
rect 12437 7219 12495 7225
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 12728 7188 12756 7287
rect 13170 7284 13176 7336
rect 13228 7324 13234 7336
rect 14918 7324 14924 7336
rect 13228 7296 14924 7324
rect 13228 7284 13234 7296
rect 14918 7284 14924 7296
rect 14976 7284 14982 7336
rect 12268 7160 12756 7188
rect 11333 7151 11391 7157
rect 552 7098 15520 7120
rect 552 7046 4100 7098
rect 4152 7046 4164 7098
rect 4216 7046 4228 7098
rect 4280 7046 4292 7098
rect 4344 7046 4356 7098
rect 4408 7046 7802 7098
rect 7854 7046 7866 7098
rect 7918 7046 7930 7098
rect 7982 7046 7994 7098
rect 8046 7046 8058 7098
rect 8110 7046 11504 7098
rect 11556 7046 11568 7098
rect 11620 7046 11632 7098
rect 11684 7046 11696 7098
rect 11748 7046 11760 7098
rect 11812 7046 15206 7098
rect 15258 7046 15270 7098
rect 15322 7046 15334 7098
rect 15386 7046 15398 7098
rect 15450 7046 15462 7098
rect 15514 7046 15520 7098
rect 552 7024 15520 7046
rect 6454 6944 6460 6996
rect 6512 6984 6518 6996
rect 6549 6987 6607 6993
rect 6549 6984 6561 6987
rect 6512 6956 6561 6984
rect 6512 6944 6518 6956
rect 6549 6953 6561 6956
rect 6595 6953 6607 6987
rect 6549 6947 6607 6953
rect 6717 6987 6775 6993
rect 6717 6953 6729 6987
rect 6763 6984 6775 6987
rect 7650 6984 7656 6996
rect 6763 6956 7656 6984
rect 6763 6953 6775 6956
rect 6717 6947 6775 6953
rect 6564 6916 6592 6947
rect 7650 6944 7656 6956
rect 7708 6944 7714 6996
rect 8113 6987 8171 6993
rect 8113 6953 8125 6987
rect 8159 6984 8171 6987
rect 8294 6984 8300 6996
rect 8159 6956 8300 6984
rect 8159 6953 8171 6956
rect 8113 6947 8171 6953
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 8386 6944 8392 6996
rect 8444 6944 8450 6996
rect 8665 6987 8723 6993
rect 8665 6953 8677 6987
rect 8711 6984 8723 6987
rect 8846 6984 8852 6996
rect 8711 6956 8852 6984
rect 8711 6953 8723 6956
rect 8665 6947 8723 6953
rect 6196 6888 6592 6916
rect 6917 6919 6975 6925
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6817 4675 6851
rect 4617 6811 4675 6817
rect 4801 6851 4859 6857
rect 4801 6817 4813 6851
rect 4847 6848 4859 6851
rect 5442 6848 5448 6860
rect 4847 6820 5448 6848
rect 4847 6817 4859 6820
rect 4801 6811 4859 6817
rect 4632 6780 4660 6811
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 6196 6857 6224 6888
rect 6917 6885 6929 6919
rect 6963 6916 6975 6919
rect 7006 6916 7012 6928
rect 6963 6888 7012 6916
rect 6963 6885 6975 6888
rect 6917 6879 6975 6885
rect 7006 6876 7012 6888
rect 7064 6876 7070 6928
rect 7561 6919 7619 6925
rect 7561 6916 7573 6919
rect 7208 6888 7573 6916
rect 5997 6851 6055 6857
rect 5997 6817 6009 6851
rect 6043 6817 6055 6851
rect 5997 6811 6055 6817
rect 6181 6851 6239 6857
rect 6181 6817 6193 6851
rect 6227 6817 6239 6851
rect 6181 6811 6239 6817
rect 5813 6783 5871 6789
rect 5813 6780 5825 6783
rect 4632 6752 5825 6780
rect 5813 6749 5825 6752
rect 5859 6749 5871 6783
rect 6012 6780 6040 6811
rect 6270 6808 6276 6860
rect 6328 6808 6334 6860
rect 6454 6808 6460 6860
rect 6512 6848 6518 6860
rect 7208 6857 7236 6888
rect 7561 6885 7573 6888
rect 7607 6916 7619 6919
rect 8202 6916 8208 6928
rect 7607 6888 8208 6916
rect 7607 6885 7619 6888
rect 7561 6879 7619 6885
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 7193 6851 7251 6857
rect 6512 6846 6592 6848
rect 6512 6820 6684 6846
rect 6512 6808 6518 6820
rect 6564 6818 6684 6820
rect 6362 6780 6368 6792
rect 6012 6752 6368 6780
rect 5813 6743 5871 6749
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 6656 6780 6684 6818
rect 7193 6817 7205 6851
rect 7239 6817 7251 6851
rect 7193 6811 7251 6817
rect 7469 6851 7527 6857
rect 7469 6817 7481 6851
rect 7515 6817 7527 6851
rect 7469 6811 7527 6817
rect 7377 6783 7435 6789
rect 7377 6780 7389 6783
rect 6656 6752 7389 6780
rect 7377 6749 7389 6752
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 7484 6780 7512 6811
rect 7650 6808 7656 6860
rect 7708 6848 7714 6860
rect 8404 6857 8432 6944
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 7708 6820 7757 6848
rect 7708 6808 7714 6820
rect 7745 6817 7757 6820
rect 7791 6817 7803 6851
rect 7745 6811 7803 6817
rect 7929 6851 7987 6857
rect 7929 6817 7941 6851
rect 7975 6848 7987 6851
rect 8389 6851 8447 6857
rect 7975 6820 8340 6848
rect 7975 6817 7987 6820
rect 7929 6811 7987 6817
rect 7944 6780 7972 6811
rect 7484 6752 7972 6780
rect 8205 6783 8263 6789
rect 6089 6715 6147 6721
rect 6089 6681 6101 6715
rect 6135 6712 6147 6715
rect 7009 6715 7067 6721
rect 7009 6712 7021 6715
rect 6135 6684 6408 6712
rect 6135 6681 6147 6684
rect 6089 6675 6147 6681
rect 4430 6604 4436 6656
rect 4488 6644 4494 6656
rect 4617 6647 4675 6653
rect 4617 6644 4629 6647
rect 4488 6616 4629 6644
rect 4488 6604 4494 6616
rect 4617 6613 4629 6616
rect 4663 6613 4675 6647
rect 6380 6644 6408 6684
rect 6564 6684 7021 6712
rect 6564 6644 6592 6684
rect 7009 6681 7021 6684
rect 7055 6681 7067 6715
rect 7009 6675 7067 6681
rect 6380 6616 6592 6644
rect 6733 6647 6791 6653
rect 4617 6607 4675 6613
rect 6733 6613 6745 6647
rect 6779 6644 6791 6647
rect 7484 6644 7512 6752
rect 8205 6749 8217 6783
rect 8251 6749 8263 6783
rect 8312 6780 8340 6820
rect 8389 6817 8401 6851
rect 8435 6817 8447 6851
rect 8389 6811 8447 6817
rect 8680 6780 8708 6947
rect 8846 6944 8852 6956
rect 8904 6944 8910 6996
rect 10781 6987 10839 6993
rect 10781 6953 10793 6987
rect 10827 6984 10839 6987
rect 10827 6956 11008 6984
rect 10827 6953 10839 6956
rect 10781 6947 10839 6953
rect 10980 6916 11008 6956
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 12066 6984 12072 6996
rect 11756 6956 12072 6984
rect 11756 6944 11762 6956
rect 12066 6944 12072 6956
rect 12124 6984 12130 6996
rect 12345 6987 12403 6993
rect 12345 6984 12357 6987
rect 12124 6956 12357 6984
rect 12124 6944 12130 6956
rect 12345 6953 12357 6956
rect 12391 6953 12403 6987
rect 13906 6984 13912 6996
rect 12345 6947 12403 6953
rect 13004 6956 13912 6984
rect 11210 6919 11268 6925
rect 11210 6916 11222 6919
rect 10060 6888 10824 6916
rect 10980 6888 11222 6916
rect 9490 6808 9496 6860
rect 9548 6848 9554 6860
rect 10060 6857 10088 6888
rect 10796 6860 10824 6888
rect 11210 6885 11222 6888
rect 11256 6885 11268 6919
rect 11210 6879 11268 6885
rect 12434 6876 12440 6928
rect 12492 6916 12498 6928
rect 12492 6888 12756 6916
rect 12492 6876 12498 6888
rect 9778 6851 9836 6857
rect 9778 6848 9790 6851
rect 9548 6820 9790 6848
rect 9548 6808 9554 6820
rect 9778 6817 9790 6820
rect 9824 6817 9836 6851
rect 9778 6811 9836 6817
rect 10045 6851 10103 6857
rect 10045 6817 10057 6851
rect 10091 6817 10103 6851
rect 10045 6811 10103 6817
rect 10226 6808 10232 6860
rect 10284 6808 10290 6860
rect 10321 6851 10379 6857
rect 10321 6817 10333 6851
rect 10367 6848 10379 6851
rect 10502 6848 10508 6860
rect 10367 6820 10508 6848
rect 10367 6817 10379 6820
rect 10321 6811 10379 6817
rect 10502 6808 10508 6820
rect 10560 6808 10566 6860
rect 10594 6808 10600 6860
rect 10652 6808 10658 6860
rect 10778 6808 10784 6860
rect 10836 6848 10842 6860
rect 10965 6851 11023 6857
rect 10965 6848 10977 6851
rect 10836 6820 10977 6848
rect 10836 6808 10842 6820
rect 10965 6817 10977 6820
rect 11011 6817 11023 6851
rect 12544 6848 12572 6888
rect 10965 6811 11023 6817
rect 11072 6820 12572 6848
rect 8312 6752 8708 6780
rect 10244 6780 10272 6808
rect 10413 6783 10471 6789
rect 10413 6780 10425 6783
rect 10244 6752 10425 6780
rect 8205 6743 8263 6749
rect 10413 6749 10425 6752
rect 10459 6780 10471 6783
rect 11072 6780 11100 6820
rect 12618 6808 12624 6860
rect 12676 6808 12682 6860
rect 12728 6857 12756 6888
rect 13004 6857 13032 6956
rect 13906 6944 13912 6956
rect 13964 6944 13970 6996
rect 13262 6876 13268 6928
rect 13320 6876 13326 6928
rect 12713 6851 12771 6857
rect 12713 6817 12725 6851
rect 12759 6817 12771 6851
rect 12713 6811 12771 6817
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6817 13047 6851
rect 12989 6811 13047 6817
rect 13078 6808 13084 6860
rect 13136 6808 13142 6860
rect 13280 6848 13308 6876
rect 13357 6851 13415 6857
rect 13357 6848 13369 6851
rect 13280 6820 13369 6848
rect 13357 6817 13369 6820
rect 13403 6817 13415 6851
rect 14090 6848 14096 6860
rect 13357 6811 13415 6817
rect 13556 6820 14096 6848
rect 10459 6752 11100 6780
rect 12437 6783 12495 6789
rect 10459 6749 10471 6752
rect 10413 6743 10471 6749
rect 12437 6749 12449 6783
rect 12483 6749 12495 6783
rect 12437 6743 12495 6749
rect 13265 6783 13323 6789
rect 13265 6749 13277 6783
rect 13311 6780 13323 6783
rect 13556 6780 13584 6820
rect 14090 6808 14096 6820
rect 14148 6808 14154 6860
rect 13311 6752 13584 6780
rect 13633 6783 13691 6789
rect 13311 6749 13323 6752
rect 13265 6743 13323 6749
rect 13633 6749 13645 6783
rect 13679 6780 13691 6783
rect 13722 6780 13728 6792
rect 13679 6752 13728 6780
rect 13679 6749 13691 6752
rect 13633 6743 13691 6749
rect 8220 6712 8248 6743
rect 9030 6712 9036 6724
rect 8220 6684 9036 6712
rect 9030 6672 9036 6684
rect 9088 6672 9094 6724
rect 12452 6712 12480 6743
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 12802 6712 12808 6724
rect 12452 6684 12808 6712
rect 12802 6672 12808 6684
rect 12860 6712 12866 6724
rect 12860 6684 13308 6712
rect 12860 6672 12866 6684
rect 6779 6616 7512 6644
rect 6779 6613 6791 6616
rect 6733 6607 6791 6613
rect 8570 6604 8576 6656
rect 8628 6604 8634 6656
rect 12526 6604 12532 6656
rect 12584 6604 12590 6656
rect 13170 6604 13176 6656
rect 13228 6604 13234 6656
rect 13280 6644 13308 6684
rect 14458 6672 14464 6724
rect 14516 6672 14522 6724
rect 14476 6644 14504 6672
rect 13280 6616 14504 6644
rect 14921 6647 14979 6653
rect 14921 6613 14933 6647
rect 14967 6644 14979 6647
rect 15010 6644 15016 6656
rect 14967 6616 15016 6644
rect 14967 6613 14979 6616
rect 14921 6607 14979 6613
rect 15010 6604 15016 6616
rect 15068 6604 15074 6656
rect 552 6554 15364 6576
rect 552 6502 2249 6554
rect 2301 6502 2313 6554
rect 2365 6502 2377 6554
rect 2429 6502 2441 6554
rect 2493 6502 2505 6554
rect 2557 6502 5951 6554
rect 6003 6502 6015 6554
rect 6067 6502 6079 6554
rect 6131 6502 6143 6554
rect 6195 6502 6207 6554
rect 6259 6502 9653 6554
rect 9705 6502 9717 6554
rect 9769 6502 9781 6554
rect 9833 6502 9845 6554
rect 9897 6502 9909 6554
rect 9961 6502 13355 6554
rect 13407 6502 13419 6554
rect 13471 6502 13483 6554
rect 13535 6502 13547 6554
rect 13599 6502 13611 6554
rect 13663 6502 15364 6554
rect 552 6480 15364 6502
rect 6365 6443 6423 6449
rect 6365 6409 6377 6443
rect 6411 6440 6423 6443
rect 6454 6440 6460 6452
rect 6411 6412 6460 6440
rect 6411 6409 6423 6412
rect 6365 6403 6423 6409
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 7377 6443 7435 6449
rect 7377 6409 7389 6443
rect 7423 6440 7435 6443
rect 9125 6443 9183 6449
rect 7423 6412 7604 6440
rect 7423 6409 7435 6412
rect 7377 6403 7435 6409
rect 7576 6384 7604 6412
rect 9125 6409 9137 6443
rect 9171 6440 9183 6443
rect 9490 6440 9496 6452
rect 9171 6412 9496 6440
rect 9171 6409 9183 6412
rect 9125 6403 9183 6409
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 10594 6400 10600 6452
rect 10652 6400 10658 6452
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6409 12311 6443
rect 12253 6403 12311 6409
rect 13541 6443 13599 6449
rect 13541 6409 13553 6443
rect 13587 6440 13599 6443
rect 13722 6440 13728 6452
rect 13587 6412 13728 6440
rect 13587 6409 13599 6412
rect 13541 6403 13599 6409
rect 5537 6375 5595 6381
rect 5537 6341 5549 6375
rect 5583 6372 5595 6375
rect 7193 6375 7251 6381
rect 5583 6344 6316 6372
rect 5583 6341 5595 6344
rect 5537 6335 5595 6341
rect 6288 6245 6316 6344
rect 7193 6341 7205 6375
rect 7239 6372 7251 6375
rect 7466 6372 7472 6384
rect 7239 6344 7472 6372
rect 7239 6341 7251 6344
rect 7193 6335 7251 6341
rect 7466 6332 7472 6344
rect 7524 6332 7530 6384
rect 7558 6332 7564 6384
rect 7616 6372 7622 6384
rect 12268 6372 12296 6403
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 12713 6375 12771 6381
rect 7616 6344 7788 6372
rect 12268 6344 12480 6372
rect 7616 6332 7622 6344
rect 7208 6276 7512 6304
rect 4157 6239 4215 6245
rect 4157 6205 4169 6239
rect 4203 6236 4215 6239
rect 6273 6239 6331 6245
rect 4203 6208 4568 6236
rect 4203 6205 4215 6208
rect 4157 6199 4215 6205
rect 4430 6177 4436 6180
rect 4424 6168 4436 6177
rect 4391 6140 4436 6168
rect 4424 6131 4436 6140
rect 4430 6128 4436 6131
rect 4488 6128 4494 6180
rect 4540 6112 4568 6208
rect 6273 6205 6285 6239
rect 6319 6236 6331 6239
rect 7006 6236 7012 6248
rect 6319 6208 7012 6236
rect 6319 6205 6331 6208
rect 6273 6199 6331 6205
rect 7006 6196 7012 6208
rect 7064 6196 7070 6248
rect 6914 6128 6920 6180
rect 6972 6168 6978 6180
rect 7208 6168 7236 6276
rect 6972 6140 7236 6168
rect 7331 6205 7389 6211
rect 7331 6171 7343 6205
rect 7377 6171 7389 6205
rect 7331 6168 7389 6171
rect 7484 6168 7512 6276
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6238 7711 6239
rect 7760 6238 7788 6344
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6304 8815 6307
rect 11882 6304 11888 6316
rect 8803 6276 11888 6304
rect 8803 6273 8815 6276
rect 8757 6267 8815 6273
rect 11882 6264 11888 6276
rect 11940 6264 11946 6316
rect 7699 6210 7788 6238
rect 7837 6239 7895 6245
rect 7699 6205 7711 6210
rect 7653 6199 7711 6205
rect 7837 6205 7849 6239
rect 7883 6205 7895 6239
rect 7837 6199 7895 6205
rect 7561 6171 7619 6177
rect 7561 6168 7573 6171
rect 7331 6165 7420 6168
rect 7360 6140 7420 6165
rect 7484 6140 7573 6168
rect 6972 6128 6978 6140
rect 4522 6060 4528 6112
rect 4580 6060 4586 6112
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 7392 6100 7420 6140
rect 7561 6137 7573 6140
rect 7607 6168 7619 6171
rect 7852 6168 7880 6199
rect 8570 6196 8576 6248
rect 8628 6236 8634 6248
rect 12158 6245 12164 6248
rect 8941 6239 8999 6245
rect 8941 6236 8953 6239
rect 8628 6208 8953 6236
rect 8628 6196 8634 6208
rect 8941 6205 8953 6208
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 10873 6239 10931 6245
rect 10873 6205 10885 6239
rect 10919 6205 10931 6239
rect 12151 6239 12164 6245
rect 12151 6236 12163 6239
rect 12119 6208 12163 6236
rect 10873 6199 10931 6205
rect 12151 6205 12163 6208
rect 12151 6199 12164 6205
rect 7607 6140 7880 6168
rect 7607 6137 7619 6140
rect 7561 6131 7619 6137
rect 8202 6128 8208 6180
rect 8260 6168 8266 6180
rect 8481 6171 8539 6177
rect 8481 6168 8493 6171
rect 8260 6140 8493 6168
rect 8260 6128 8266 6140
rect 8481 6137 8493 6140
rect 8527 6137 8539 6171
rect 8481 6131 8539 6137
rect 10502 6128 10508 6180
rect 10560 6168 10566 6180
rect 10597 6171 10655 6177
rect 10597 6168 10609 6171
rect 10560 6140 10609 6168
rect 10560 6128 10566 6140
rect 10597 6137 10609 6140
rect 10643 6168 10655 6171
rect 10686 6168 10692 6180
rect 10643 6140 10692 6168
rect 10643 6137 10655 6140
rect 10597 6131 10655 6137
rect 10686 6128 10692 6140
rect 10744 6128 10750 6180
rect 10888 6168 10916 6199
rect 12158 6196 12164 6199
rect 12216 6196 12222 6248
rect 12452 6245 12480 6344
rect 12713 6341 12725 6375
rect 12759 6372 12771 6375
rect 12986 6372 12992 6384
rect 12759 6344 12992 6372
rect 12759 6341 12771 6344
rect 12713 6335 12771 6341
rect 12986 6332 12992 6344
rect 13044 6332 13050 6384
rect 12345 6239 12403 6245
rect 12345 6205 12357 6239
rect 12391 6205 12403 6239
rect 12345 6199 12403 6205
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6205 12495 6239
rect 12437 6199 12495 6205
rect 11330 6168 11336 6180
rect 10888 6140 11336 6168
rect 11330 6128 11336 6140
rect 11388 6168 11394 6180
rect 11698 6168 11704 6180
rect 11388 6140 11704 6168
rect 11388 6128 11394 6140
rect 11698 6128 11704 6140
rect 11756 6128 11762 6180
rect 7340 6072 7420 6100
rect 7340 6060 7346 6072
rect 7742 6060 7748 6112
rect 7800 6060 7806 6112
rect 10781 6103 10839 6109
rect 10781 6069 10793 6103
rect 10827 6100 10839 6103
rect 10870 6100 10876 6112
rect 10827 6072 10876 6100
rect 10827 6069 10839 6072
rect 10781 6063 10839 6069
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 11882 6060 11888 6112
rect 11940 6100 11946 6112
rect 12360 6100 12388 6199
rect 12526 6196 12532 6248
rect 12584 6196 12590 6248
rect 12713 6239 12771 6245
rect 12713 6205 12725 6239
rect 12759 6236 12771 6239
rect 12894 6236 12900 6248
rect 12759 6208 12900 6236
rect 12759 6205 12771 6208
rect 12713 6199 12771 6205
rect 12894 6196 12900 6208
rect 12952 6196 12958 6248
rect 13078 6196 13084 6248
rect 13136 6196 13142 6248
rect 13170 6196 13176 6248
rect 13228 6236 13234 6248
rect 13541 6239 13599 6245
rect 13541 6236 13553 6239
rect 13228 6208 13553 6236
rect 13228 6196 13234 6208
rect 13541 6205 13553 6208
rect 13587 6205 13599 6239
rect 13541 6199 13599 6205
rect 13817 6239 13875 6245
rect 13817 6205 13829 6239
rect 13863 6205 13875 6239
rect 13817 6199 13875 6205
rect 13096 6168 13124 6196
rect 13832 6168 13860 6199
rect 13906 6196 13912 6248
rect 13964 6196 13970 6248
rect 13096 6140 13860 6168
rect 13725 6103 13783 6109
rect 13725 6100 13737 6103
rect 11940 6072 13737 6100
rect 11940 6060 11946 6072
rect 13725 6069 13737 6072
rect 13771 6100 13783 6103
rect 13924 6100 13952 6196
rect 13771 6072 13952 6100
rect 13771 6069 13783 6072
rect 13725 6063 13783 6069
rect 552 6010 15520 6032
rect 552 5958 4100 6010
rect 4152 5958 4164 6010
rect 4216 5958 4228 6010
rect 4280 5958 4292 6010
rect 4344 5958 4356 6010
rect 4408 5958 7802 6010
rect 7854 5958 7866 6010
rect 7918 5958 7930 6010
rect 7982 5958 7994 6010
rect 8046 5958 8058 6010
rect 8110 5958 11504 6010
rect 11556 5958 11568 6010
rect 11620 5958 11632 6010
rect 11684 5958 11696 6010
rect 11748 5958 11760 6010
rect 11812 5958 15206 6010
rect 15258 5958 15270 6010
rect 15322 5958 15334 6010
rect 15386 5958 15398 6010
rect 15450 5958 15462 6010
rect 15514 5958 15520 6010
rect 552 5936 15520 5958
rect 10778 5856 10784 5908
rect 10836 5896 10842 5908
rect 11974 5896 11980 5908
rect 10836 5868 11980 5896
rect 10836 5856 10842 5868
rect 11974 5856 11980 5868
rect 12032 5896 12038 5908
rect 12032 5868 12756 5896
rect 12032 5856 12038 5868
rect 7561 5831 7619 5837
rect 7561 5797 7573 5831
rect 7607 5828 7619 5831
rect 8938 5828 8944 5840
rect 7607 5800 8944 5828
rect 7607 5797 7619 5800
rect 7561 5791 7619 5797
rect 8938 5788 8944 5800
rect 8996 5828 9002 5840
rect 10965 5831 11023 5837
rect 10965 5828 10977 5831
rect 8996 5800 10977 5828
rect 8996 5788 9002 5800
rect 10965 5797 10977 5800
rect 11011 5797 11023 5831
rect 10965 5791 11023 5797
rect 4516 5763 4574 5769
rect 4516 5729 4528 5763
rect 4562 5760 4574 5763
rect 5534 5760 5540 5772
rect 4562 5732 5540 5760
rect 4562 5729 4574 5732
rect 4516 5723 4574 5729
rect 5534 5720 5540 5732
rect 5592 5720 5598 5772
rect 7374 5720 7380 5772
rect 7432 5760 7438 5772
rect 7837 5763 7895 5769
rect 7837 5760 7849 5763
rect 7432 5732 7849 5760
rect 7432 5720 7438 5732
rect 7837 5729 7849 5732
rect 7883 5760 7895 5763
rect 8202 5760 8208 5772
rect 7883 5732 8208 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 12728 5769 12756 5868
rect 12713 5763 12771 5769
rect 12713 5729 12725 5763
rect 12759 5760 12771 5763
rect 12805 5763 12863 5769
rect 12805 5760 12817 5763
rect 12759 5732 12817 5760
rect 12759 5729 12771 5732
rect 12713 5723 12771 5729
rect 12805 5729 12817 5732
rect 12851 5760 12863 5763
rect 12851 5732 13308 5760
rect 12851 5729 12863 5732
rect 12805 5723 12863 5729
rect 13280 5704 13308 5732
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5661 4307 5695
rect 8018 5692 8024 5704
rect 4249 5655 4307 5661
rect 6288 5664 8024 5692
rect 4264 5556 4292 5655
rect 6288 5633 6316 5664
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 12986 5652 12992 5704
rect 13044 5692 13050 5704
rect 13081 5695 13139 5701
rect 13081 5692 13093 5695
rect 13044 5664 13093 5692
rect 13044 5652 13050 5664
rect 13081 5661 13093 5664
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 13262 5652 13268 5704
rect 13320 5652 13326 5704
rect 6273 5627 6331 5633
rect 6273 5624 6285 5627
rect 5506 5596 6285 5624
rect 4522 5556 4528 5568
rect 4264 5528 4528 5556
rect 4522 5516 4528 5528
rect 4580 5556 4586 5568
rect 5506 5556 5534 5596
rect 6273 5593 6285 5596
rect 6319 5593 6331 5627
rect 6273 5587 6331 5593
rect 6362 5584 6368 5636
rect 6420 5624 6426 5636
rect 6420 5596 8064 5624
rect 6420 5584 6426 5596
rect 4580 5528 5534 5556
rect 5629 5559 5687 5565
rect 4580 5516 4586 5528
rect 5629 5525 5641 5559
rect 5675 5556 5687 5559
rect 6914 5556 6920 5568
rect 5675 5528 6920 5556
rect 5675 5525 5687 5528
rect 5629 5519 5687 5525
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 8036 5565 8064 5596
rect 8021 5559 8079 5565
rect 8021 5525 8033 5559
rect 8067 5556 8079 5559
rect 8202 5556 8208 5568
rect 8067 5528 8208 5556
rect 8067 5525 8079 5528
rect 8021 5519 8079 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 10870 5516 10876 5568
rect 10928 5556 10934 5568
rect 12066 5556 12072 5568
rect 10928 5528 12072 5556
rect 10928 5516 10934 5528
rect 12066 5516 12072 5528
rect 12124 5516 12130 5568
rect 14369 5559 14427 5565
rect 14369 5525 14381 5559
rect 14415 5556 14427 5559
rect 14458 5556 14464 5568
rect 14415 5528 14464 5556
rect 14415 5525 14427 5528
rect 14369 5519 14427 5525
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 552 5466 15364 5488
rect 552 5414 2249 5466
rect 2301 5414 2313 5466
rect 2365 5414 2377 5466
rect 2429 5414 2441 5466
rect 2493 5414 2505 5466
rect 2557 5414 5951 5466
rect 6003 5414 6015 5466
rect 6067 5414 6079 5466
rect 6131 5414 6143 5466
rect 6195 5414 6207 5466
rect 6259 5414 9653 5466
rect 9705 5414 9717 5466
rect 9769 5414 9781 5466
rect 9833 5414 9845 5466
rect 9897 5414 9909 5466
rect 9961 5414 13355 5466
rect 13407 5414 13419 5466
rect 13471 5414 13483 5466
rect 13535 5414 13547 5466
rect 13599 5414 13611 5466
rect 13663 5414 15364 5466
rect 552 5392 15364 5414
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 5997 5355 6055 5361
rect 5997 5352 6009 5355
rect 5592 5324 6009 5352
rect 5592 5312 5598 5324
rect 5997 5321 6009 5324
rect 6043 5321 6055 5355
rect 5997 5315 6055 5321
rect 8220 5324 10364 5352
rect 8220 5296 8248 5324
rect 8202 5244 8208 5296
rect 8260 5244 8266 5296
rect 10336 5284 10364 5324
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 12434 5352 12440 5364
rect 11388 5324 12440 5352
rect 11388 5312 11394 5324
rect 12434 5312 12440 5324
rect 12492 5312 12498 5364
rect 13357 5287 13415 5293
rect 13357 5284 13369 5287
rect 10336 5256 11008 5284
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7285 5219 7343 5225
rect 7285 5216 7297 5219
rect 6972 5188 7297 5216
rect 6972 5176 6978 5188
rect 7285 5185 7297 5188
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 8018 5176 8024 5228
rect 8076 5216 8082 5228
rect 8665 5219 8723 5225
rect 8665 5216 8677 5219
rect 8076 5188 8677 5216
rect 8076 5176 8082 5188
rect 8665 5185 8677 5188
rect 8711 5185 8723 5219
rect 8665 5179 8723 5185
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5185 10195 5219
rect 10137 5179 10195 5185
rect 5626 5108 5632 5160
rect 5684 5148 5690 5160
rect 5810 5148 5816 5160
rect 5684 5120 5816 5148
rect 5684 5108 5690 5120
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 5994 5108 6000 5160
rect 6052 5108 6058 5160
rect 6273 5151 6331 5157
rect 6273 5117 6285 5151
rect 6319 5148 6331 5151
rect 6365 5151 6423 5157
rect 6365 5148 6377 5151
rect 6319 5120 6377 5148
rect 6319 5117 6331 5120
rect 6273 5111 6331 5117
rect 6365 5117 6377 5120
rect 6411 5117 6423 5151
rect 6365 5111 6423 5117
rect 7469 5151 7527 5157
rect 7469 5117 7481 5151
rect 7515 5148 7527 5151
rect 8294 5148 8300 5160
rect 7515 5120 8300 5148
rect 7515 5117 7527 5120
rect 7469 5111 7527 5117
rect 8294 5108 8300 5120
rect 8352 5108 8358 5160
rect 8389 5151 8447 5157
rect 8389 5117 8401 5151
rect 8435 5117 8447 5151
rect 8389 5111 8447 5117
rect 8573 5151 8631 5157
rect 8573 5117 8585 5151
rect 8619 5148 8631 5151
rect 10152 5148 10180 5179
rect 10336 5157 10364 5256
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 8619 5120 10180 5148
rect 10321 5151 10379 5157
rect 8619 5117 8631 5120
rect 8573 5111 8631 5117
rect 10321 5117 10333 5151
rect 10367 5117 10379 5151
rect 10321 5111 10379 5117
rect 7742 5080 7748 5092
rect 7300 5052 7748 5080
rect 7300 5024 7328 5052
rect 7742 5040 7748 5052
rect 7800 5080 7806 5092
rect 7837 5083 7895 5089
rect 7837 5080 7849 5083
rect 7800 5052 7849 5080
rect 7800 5040 7806 5052
rect 7837 5049 7849 5052
rect 7883 5049 7895 5083
rect 7837 5043 7895 5049
rect 6181 5015 6239 5021
rect 6181 4981 6193 5015
rect 6227 5012 6239 5015
rect 6546 5012 6552 5024
rect 6227 4984 6552 5012
rect 6227 4981 6239 4984
rect 6181 4975 6239 4981
rect 6546 4972 6552 4984
rect 6604 4972 6610 5024
rect 7282 4972 7288 5024
rect 7340 4972 7346 5024
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 7561 5015 7619 5021
rect 7561 5012 7573 5015
rect 7524 4984 7573 5012
rect 7524 4972 7530 4984
rect 7561 4981 7573 4984
rect 7607 4981 7619 5015
rect 7561 4975 7619 4981
rect 7650 4972 7656 5024
rect 7708 4972 7714 5024
rect 8404 5012 8432 5111
rect 10410 5108 10416 5160
rect 10468 5108 10474 5160
rect 10520 5148 10548 5179
rect 10594 5176 10600 5228
rect 10652 5176 10658 5228
rect 10686 5148 10692 5160
rect 10520 5120 10692 5148
rect 10686 5108 10692 5120
rect 10744 5108 10750 5160
rect 10778 5108 10784 5160
rect 10836 5108 10842 5160
rect 10873 5151 10931 5157
rect 10873 5117 10885 5151
rect 10919 5117 10931 5151
rect 10980 5148 11008 5256
rect 11992 5256 13369 5284
rect 11992 5225 12020 5256
rect 13357 5253 13369 5256
rect 13403 5253 13415 5287
rect 13357 5247 13415 5253
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5185 12035 5219
rect 11977 5179 12035 5185
rect 12066 5176 12072 5228
rect 12124 5176 12130 5228
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5216 13047 5219
rect 13035 5188 13584 5216
rect 13035 5185 13047 5188
rect 12989 5179 13047 5185
rect 11793 5151 11851 5157
rect 11793 5148 11805 5151
rect 10980 5120 11805 5148
rect 10873 5111 10931 5117
rect 11793 5117 11805 5120
rect 11839 5117 11851 5151
rect 11793 5111 11851 5117
rect 8481 5083 8539 5089
rect 8481 5049 8493 5083
rect 8527 5080 8539 5083
rect 8910 5083 8968 5089
rect 8910 5080 8922 5083
rect 8527 5052 8922 5080
rect 8527 5049 8539 5052
rect 8481 5043 8539 5049
rect 8910 5049 8922 5052
rect 8956 5049 8968 5083
rect 10888 5080 10916 5111
rect 11882 5108 11888 5160
rect 11940 5108 11946 5160
rect 12253 5151 12311 5157
rect 12253 5117 12265 5151
rect 12299 5117 12311 5151
rect 12253 5111 12311 5117
rect 8910 5043 8968 5049
rect 10060 5052 10916 5080
rect 10060 5024 10088 5052
rect 11238 5040 11244 5092
rect 11296 5080 11302 5092
rect 12268 5080 12296 5111
rect 12342 5108 12348 5160
rect 12400 5108 12406 5160
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 13556 5157 13584 5188
rect 13081 5151 13139 5157
rect 13081 5148 13093 5151
rect 12492 5120 13093 5148
rect 12492 5108 12498 5120
rect 13081 5117 13093 5120
rect 13127 5117 13139 5151
rect 13081 5111 13139 5117
rect 13541 5151 13599 5157
rect 13541 5117 13553 5151
rect 13587 5117 13599 5151
rect 13541 5111 13599 5117
rect 11296 5052 12020 5080
rect 12268 5052 13308 5080
rect 11296 5040 11302 5052
rect 9950 5012 9956 5024
rect 8404 4984 9956 5012
rect 9950 4972 9956 4984
rect 10008 4972 10014 5024
rect 10042 4972 10048 5024
rect 10100 4972 10106 5024
rect 11422 4972 11428 5024
rect 11480 5012 11486 5024
rect 11517 5015 11575 5021
rect 11517 5012 11529 5015
rect 11480 4984 11529 5012
rect 11480 4972 11486 4984
rect 11517 4981 11529 4984
rect 11563 4981 11575 5015
rect 11517 4975 11575 4981
rect 11609 5015 11667 5021
rect 11609 4981 11621 5015
rect 11655 5012 11667 5015
rect 11882 5012 11888 5024
rect 11655 4984 11888 5012
rect 11655 4981 11667 4984
rect 11609 4975 11667 4981
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 11992 5012 12020 5052
rect 13173 5015 13231 5021
rect 13173 5012 13185 5015
rect 11992 4984 13185 5012
rect 13173 4981 13185 4984
rect 13219 4981 13231 5015
rect 13280 5012 13308 5052
rect 13354 5040 13360 5092
rect 13412 5040 13418 5092
rect 13633 5015 13691 5021
rect 13633 5012 13645 5015
rect 13280 4984 13645 5012
rect 13173 4975 13231 4981
rect 13633 4981 13645 4984
rect 13679 4981 13691 5015
rect 13633 4975 13691 4981
rect 552 4922 15520 4944
rect 552 4870 4100 4922
rect 4152 4870 4164 4922
rect 4216 4870 4228 4922
rect 4280 4870 4292 4922
rect 4344 4870 4356 4922
rect 4408 4870 7802 4922
rect 7854 4870 7866 4922
rect 7918 4870 7930 4922
rect 7982 4870 7994 4922
rect 8046 4870 8058 4922
rect 8110 4870 11504 4922
rect 11556 4870 11568 4922
rect 11620 4870 11632 4922
rect 11684 4870 11696 4922
rect 11748 4870 11760 4922
rect 11812 4870 15206 4922
rect 15258 4870 15270 4922
rect 15322 4870 15334 4922
rect 15386 4870 15398 4922
rect 15450 4870 15462 4922
rect 15514 4870 15520 4922
rect 552 4848 15520 4870
rect 5994 4768 6000 4820
rect 6052 4808 6058 4820
rect 6181 4811 6239 4817
rect 6181 4808 6193 4811
rect 6052 4780 6193 4808
rect 6052 4768 6058 4780
rect 6181 4777 6193 4780
rect 6227 4777 6239 4811
rect 6181 4771 6239 4777
rect 6546 4768 6552 4820
rect 6604 4768 6610 4820
rect 7558 4768 7564 4820
rect 7616 4768 7622 4820
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 8205 4811 8263 4817
rect 8205 4808 8217 4811
rect 7708 4780 8217 4808
rect 7708 4768 7714 4780
rect 8205 4777 8217 4780
rect 8251 4777 8263 4811
rect 8205 4771 8263 4777
rect 8294 4768 8300 4820
rect 8352 4768 8358 4820
rect 10413 4811 10471 4817
rect 10413 4777 10425 4811
rect 10459 4808 10471 4811
rect 10870 4808 10876 4820
rect 10459 4780 10876 4808
rect 10459 4777 10471 4780
rect 10413 4771 10471 4777
rect 5445 4743 5503 4749
rect 5445 4709 5457 4743
rect 5491 4740 5503 4743
rect 6270 4740 6276 4752
rect 5491 4712 6276 4740
rect 5491 4709 5503 4712
rect 5445 4703 5503 4709
rect 6270 4700 6276 4712
rect 6328 4700 6334 4752
rect 6564 4740 6592 4768
rect 7576 4740 7604 4768
rect 6564 4712 6868 4740
rect 4982 4632 4988 4684
rect 5040 4672 5046 4684
rect 5261 4675 5319 4681
rect 5261 4672 5273 4675
rect 5040 4644 5273 4672
rect 5040 4632 5046 4644
rect 5261 4641 5273 4644
rect 5307 4672 5319 4675
rect 5350 4672 5356 4684
rect 5307 4644 5356 4672
rect 5307 4641 5319 4644
rect 5261 4635 5319 4641
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 5537 4675 5595 4681
rect 5537 4641 5549 4675
rect 5583 4641 5595 4675
rect 5537 4635 5595 4641
rect 5258 4428 5264 4480
rect 5316 4428 5322 4480
rect 5552 4468 5580 4635
rect 6362 4632 6368 4684
rect 6420 4632 6426 4684
rect 6638 4632 6644 4684
rect 6696 4632 6702 4684
rect 6840 4681 6868 4712
rect 7208 4712 7604 4740
rect 7208 4681 7236 4712
rect 7834 4700 7840 4752
rect 7892 4740 7898 4752
rect 8312 4740 8340 4768
rect 7892 4712 8340 4740
rect 7892 4700 7898 4712
rect 6825 4675 6883 4681
rect 6825 4641 6837 4675
rect 6871 4641 6883 4675
rect 6825 4635 6883 4641
rect 7193 4675 7251 4681
rect 7193 4641 7205 4675
rect 7239 4641 7251 4675
rect 7193 4635 7251 4641
rect 7374 4632 7380 4684
rect 7432 4632 7438 4684
rect 7469 4675 7527 4681
rect 7469 4641 7481 4675
rect 7515 4641 7527 4675
rect 7469 4635 7527 4641
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4604 6607 4607
rect 7282 4604 7288 4616
rect 6595 4576 7288 4604
rect 6595 4573 6607 4576
rect 6549 4567 6607 4573
rect 7282 4564 7288 4576
rect 7340 4564 7346 4616
rect 6457 4539 6515 4545
rect 6457 4505 6469 4539
rect 6503 4536 6515 4539
rect 7392 4536 7420 4632
rect 7484 4548 7512 4635
rect 7558 4632 7564 4684
rect 7616 4672 7622 4684
rect 7745 4675 7803 4681
rect 7745 4672 7757 4675
rect 7616 4644 7757 4672
rect 7616 4632 7622 4644
rect 7745 4641 7757 4644
rect 7791 4641 7803 4675
rect 7745 4635 7803 4641
rect 6503 4508 7420 4536
rect 6503 4505 6515 4508
rect 6457 4499 6515 4505
rect 7466 4496 7472 4548
rect 7524 4496 7530 4548
rect 6917 4471 6975 4477
rect 6917 4468 6929 4471
rect 5552 4440 6929 4468
rect 6917 4437 6929 4440
rect 6963 4437 6975 4471
rect 6917 4431 6975 4437
rect 7190 4428 7196 4480
rect 7248 4428 7254 4480
rect 7760 4468 7788 4635
rect 7926 4632 7932 4684
rect 7984 4672 7990 4684
rect 8389 4675 8447 4681
rect 8389 4672 8401 4675
rect 7984 4644 8401 4672
rect 7984 4632 7990 4644
rect 8389 4641 8401 4644
rect 8435 4641 8447 4675
rect 8389 4635 8447 4641
rect 10042 4632 10048 4684
rect 10100 4672 10106 4684
rect 10137 4675 10195 4681
rect 10137 4672 10149 4675
rect 10100 4644 10149 4672
rect 10100 4632 10106 4644
rect 10137 4641 10149 4644
rect 10183 4641 10195 4675
rect 10137 4635 10195 4641
rect 10321 4675 10379 4681
rect 10321 4641 10333 4675
rect 10367 4672 10379 4675
rect 10428 4672 10456 4771
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 11238 4768 11244 4820
rect 11296 4768 11302 4820
rect 11330 4768 11336 4820
rect 11388 4768 11394 4820
rect 12342 4808 12348 4820
rect 11716 4780 12348 4808
rect 10581 4743 10639 4749
rect 10581 4709 10593 4743
rect 10627 4740 10639 4743
rect 10781 4743 10839 4749
rect 10627 4712 10732 4740
rect 10627 4709 10639 4712
rect 10581 4703 10639 4709
rect 10367 4644 10456 4672
rect 10704 4672 10732 4712
rect 10781 4709 10793 4743
rect 10827 4740 10839 4743
rect 11149 4743 11207 4749
rect 11149 4740 11161 4743
rect 10827 4712 11161 4740
rect 10827 4709 10839 4712
rect 10781 4703 10839 4709
rect 11149 4709 11161 4712
rect 11195 4740 11207 4743
rect 11716 4740 11744 4780
rect 12342 4768 12348 4780
rect 12400 4808 12406 4820
rect 13354 4808 13360 4820
rect 12400 4780 13360 4808
rect 12400 4768 12406 4780
rect 13354 4768 13360 4780
rect 13412 4768 13418 4820
rect 11195 4712 11744 4740
rect 11195 4709 11207 4712
rect 11149 4703 11207 4709
rect 11790 4700 11796 4752
rect 11848 4740 11854 4752
rect 12222 4743 12280 4749
rect 12222 4740 12234 4743
rect 11848 4712 12234 4740
rect 11848 4700 11854 4712
rect 12222 4709 12234 4712
rect 12268 4709 12280 4743
rect 12222 4703 12280 4709
rect 11330 4672 11336 4684
rect 10704 4644 11336 4672
rect 10367 4641 10379 4644
rect 10321 4635 10379 4641
rect 8110 4564 8116 4616
rect 8168 4604 8174 4616
rect 8573 4607 8631 4613
rect 8573 4604 8585 4607
rect 8168 4576 8585 4604
rect 8168 4564 8174 4576
rect 8573 4573 8585 4576
rect 8619 4573 8631 4607
rect 10152 4604 10180 4635
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 11422 4632 11428 4684
rect 11480 4672 11486 4684
rect 11701 4675 11759 4681
rect 11701 4672 11713 4675
rect 11480 4644 11713 4672
rect 11480 4632 11486 4644
rect 11701 4641 11713 4644
rect 11747 4641 11759 4675
rect 11701 4635 11759 4641
rect 11974 4632 11980 4684
rect 12032 4632 12038 4684
rect 10965 4607 11023 4613
rect 10965 4604 10977 4607
rect 10152 4576 10977 4604
rect 8573 4567 8631 4573
rect 10965 4573 10977 4576
rect 11011 4573 11023 4607
rect 10965 4567 11023 4573
rect 11440 4576 11836 4604
rect 10321 4539 10379 4545
rect 10321 4505 10333 4539
rect 10367 4536 10379 4539
rect 10686 4536 10692 4548
rect 10367 4508 10692 4536
rect 10367 4505 10379 4508
rect 10321 4499 10379 4505
rect 10686 4496 10692 4508
rect 10744 4496 10750 4548
rect 10778 4496 10784 4548
rect 10836 4536 10842 4548
rect 11440 4536 11468 4576
rect 10836 4508 11468 4536
rect 10836 4496 10842 4508
rect 11514 4496 11520 4548
rect 11572 4496 11578 4548
rect 11808 4545 11836 4576
rect 11793 4539 11851 4545
rect 11793 4505 11805 4539
rect 11839 4505 11851 4539
rect 11793 4499 11851 4505
rect 9490 4468 9496 4480
rect 7760 4440 9496 4468
rect 9490 4428 9496 4440
rect 9548 4428 9554 4480
rect 10597 4471 10655 4477
rect 10597 4437 10609 4471
rect 10643 4468 10655 4471
rect 11238 4468 11244 4480
rect 10643 4440 11244 4468
rect 10643 4437 10655 4440
rect 10597 4431 10655 4437
rect 11238 4428 11244 4440
rect 11296 4428 11302 4480
rect 552 4378 15364 4400
rect 552 4326 2249 4378
rect 2301 4326 2313 4378
rect 2365 4326 2377 4378
rect 2429 4326 2441 4378
rect 2493 4326 2505 4378
rect 2557 4326 5951 4378
rect 6003 4326 6015 4378
rect 6067 4326 6079 4378
rect 6131 4326 6143 4378
rect 6195 4326 6207 4378
rect 6259 4326 9653 4378
rect 9705 4326 9717 4378
rect 9769 4326 9781 4378
rect 9833 4326 9845 4378
rect 9897 4326 9909 4378
rect 9961 4326 13355 4378
rect 13407 4326 13419 4378
rect 13471 4326 13483 4378
rect 13535 4326 13547 4378
rect 13599 4326 13611 4378
rect 13663 4326 15364 4378
rect 552 4304 15364 4326
rect 5350 4224 5356 4276
rect 5408 4264 5414 4276
rect 5408 4236 6224 4264
rect 5408 4224 5414 4236
rect 5629 4199 5687 4205
rect 5629 4165 5641 4199
rect 5675 4165 5687 4199
rect 6196 4196 6224 4236
rect 6270 4224 6276 4276
rect 6328 4264 6334 4276
rect 6641 4267 6699 4273
rect 6641 4264 6653 4267
rect 6328 4236 6653 4264
rect 6328 4224 6334 4236
rect 6641 4233 6653 4236
rect 6687 4233 6699 4267
rect 6641 4227 6699 4233
rect 6917 4267 6975 4273
rect 6917 4233 6929 4267
rect 6963 4264 6975 4267
rect 7466 4264 7472 4276
rect 6963 4236 7472 4264
rect 6963 4233 6975 4236
rect 6917 4227 6975 4233
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 11330 4224 11336 4276
rect 11388 4224 11394 4276
rect 11701 4267 11759 4273
rect 11701 4233 11713 4267
rect 11747 4264 11759 4267
rect 11790 4264 11796 4276
rect 11747 4236 11796 4264
rect 11747 4233 11759 4236
rect 11701 4227 11759 4233
rect 11790 4224 11796 4236
rect 11848 4224 11854 4276
rect 11882 4224 11888 4276
rect 11940 4224 11946 4276
rect 8754 4196 8760 4208
rect 6196 4168 8760 4196
rect 5629 4159 5687 4165
rect 5644 4128 5672 4159
rect 8754 4156 8760 4168
rect 8812 4156 8818 4208
rect 8938 4156 8944 4208
rect 8996 4156 9002 4208
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5644 4100 5917 4128
rect 5905 4097 5917 4100
rect 5951 4128 5963 4131
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 5951 4100 7389 4128
rect 5951 4097 5963 4100
rect 5905 4091 5963 4097
rect 7377 4097 7389 4100
rect 7423 4128 7435 4131
rect 8110 4128 8116 4140
rect 7423 4100 8116 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 11057 4131 11115 4137
rect 8312 4100 9352 4128
rect 4249 4063 4307 4069
rect 4249 4029 4261 4063
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 4516 4063 4574 4069
rect 4516 4029 4528 4063
rect 4562 4060 4574 4063
rect 5258 4060 5264 4072
rect 4562 4032 5264 4060
rect 4562 4029 4574 4032
rect 4516 4023 4574 4029
rect 4264 3992 4292 4023
rect 5258 4020 5264 4032
rect 5316 4020 5322 4072
rect 5718 4020 5724 4072
rect 5776 4020 5782 4072
rect 6457 4063 6515 4069
rect 6457 4029 6469 4063
rect 6503 4060 6515 4063
rect 6549 4063 6607 4069
rect 6549 4060 6561 4063
rect 6503 4032 6561 4060
rect 6503 4029 6515 4032
rect 6457 4023 6515 4029
rect 6549 4029 6561 4032
rect 6595 4029 6607 4063
rect 6724 4063 6782 4069
rect 6724 4060 6736 4063
rect 6549 4023 6607 4029
rect 6656 4032 6736 4060
rect 5736 3992 5764 4020
rect 6656 4004 6684 4032
rect 6724 4029 6736 4032
rect 6770 4029 6782 4063
rect 6724 4023 6782 4029
rect 7101 4063 7159 4069
rect 7101 4029 7113 4063
rect 7147 4029 7159 4063
rect 7101 4023 7159 4029
rect 7193 4063 7251 4069
rect 7193 4029 7205 4063
rect 7239 4029 7251 4063
rect 7193 4023 7251 4029
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4060 7343 4063
rect 7926 4060 7932 4072
rect 7331 4032 7932 4060
rect 7331 4029 7343 4032
rect 7285 4023 7343 4029
rect 6638 3992 6644 4004
rect 4264 3964 4568 3992
rect 5736 3964 6644 3992
rect 4540 3936 4568 3964
rect 6638 3952 6644 3964
rect 6696 3952 6702 4004
rect 4522 3884 4528 3936
rect 4580 3884 4586 3936
rect 7116 3924 7144 4023
rect 7208 3992 7236 4023
rect 7926 4020 7932 4032
rect 7984 4060 7990 4072
rect 8202 4060 8208 4072
rect 7984 4032 8208 4060
rect 7984 4020 7990 4032
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 7650 3992 7656 4004
rect 7208 3964 7656 3992
rect 7650 3952 7656 3964
rect 7708 3992 7714 4004
rect 7834 3992 7840 4004
rect 7708 3964 7840 3992
rect 7708 3952 7714 3964
rect 7834 3952 7840 3964
rect 7892 3992 7898 4004
rect 8312 3992 8340 4100
rect 9214 4020 9220 4072
rect 9272 4020 9278 4072
rect 9324 4069 9352 4100
rect 11057 4097 11069 4131
rect 11103 4128 11115 4131
rect 11348 4128 11376 4224
rect 11900 4128 11928 4224
rect 11103 4100 11376 4128
rect 11716 4100 11928 4128
rect 11103 4097 11115 4100
rect 11057 4091 11115 4097
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4029 9367 4063
rect 9309 4023 9367 4029
rect 9490 4020 9496 4072
rect 9548 4060 9554 4072
rect 10410 4060 10416 4072
rect 9548 4032 10416 4060
rect 9548 4020 9554 4032
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 10502 4020 10508 4072
rect 10560 4020 10566 4072
rect 10965 4063 11023 4069
rect 10965 4029 10977 4063
rect 11011 4060 11023 4063
rect 11238 4060 11244 4072
rect 11011 4032 11244 4060
rect 11011 4029 11023 4032
rect 10965 4023 11023 4029
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 11716 4069 11744 4100
rect 11701 4063 11759 4069
rect 11701 4029 11713 4063
rect 11747 4029 11759 4063
rect 11701 4023 11759 4029
rect 11882 4020 11888 4072
rect 11940 4060 11946 4072
rect 12894 4060 12900 4072
rect 11940 4032 12900 4060
rect 11940 4020 11946 4032
rect 12894 4020 12900 4032
rect 12952 4020 12958 4072
rect 7892 3964 8340 3992
rect 7892 3952 7898 3964
rect 8754 3952 8760 4004
rect 8812 3992 8818 4004
rect 8941 3995 8999 4001
rect 8941 3992 8953 3995
rect 8812 3964 8953 3992
rect 8812 3952 8818 3964
rect 8941 3961 8953 3964
rect 8987 3992 8999 3995
rect 10520 3992 10548 4020
rect 8987 3964 10548 3992
rect 8987 3961 8999 3964
rect 8941 3955 8999 3961
rect 7558 3924 7564 3936
rect 7116 3896 7564 3924
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 9122 3884 9128 3936
rect 9180 3884 9186 3936
rect 9398 3884 9404 3936
rect 9456 3884 9462 3936
rect 11330 3884 11336 3936
rect 11388 3884 11394 3936
rect 552 3834 15520 3856
rect 552 3782 4100 3834
rect 4152 3782 4164 3834
rect 4216 3782 4228 3834
rect 4280 3782 4292 3834
rect 4344 3782 4356 3834
rect 4408 3782 7802 3834
rect 7854 3782 7866 3834
rect 7918 3782 7930 3834
rect 7982 3782 7994 3834
rect 8046 3782 8058 3834
rect 8110 3782 11504 3834
rect 11556 3782 11568 3834
rect 11620 3782 11632 3834
rect 11684 3782 11696 3834
rect 11748 3782 11760 3834
rect 11812 3782 15206 3834
rect 15258 3782 15270 3834
rect 15322 3782 15334 3834
rect 15386 3782 15398 3834
rect 15450 3782 15462 3834
rect 15514 3782 15520 3834
rect 552 3760 15520 3782
rect 7558 3680 7564 3732
rect 7616 3680 7622 3732
rect 8113 3723 8171 3729
rect 8113 3689 8125 3723
rect 8159 3720 8171 3723
rect 9122 3720 9128 3732
rect 8159 3692 9128 3720
rect 8159 3689 8171 3692
rect 8113 3683 8171 3689
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9214 3680 9220 3732
rect 9272 3720 9278 3732
rect 9585 3723 9643 3729
rect 9585 3720 9597 3723
rect 9272 3692 9597 3720
rect 9272 3680 9278 3692
rect 9585 3689 9597 3692
rect 9631 3689 9643 3723
rect 9585 3683 9643 3689
rect 9953 3723 10011 3729
rect 9953 3689 9965 3723
rect 9999 3720 10011 3723
rect 10226 3720 10232 3732
rect 9999 3692 10232 3720
rect 9999 3689 10011 3692
rect 9953 3683 10011 3689
rect 10226 3680 10232 3692
rect 10284 3720 10290 3732
rect 11149 3723 11207 3729
rect 10284 3692 10640 3720
rect 10284 3680 10290 3692
rect 7576 3584 7604 3680
rect 7745 3655 7803 3661
rect 7745 3621 7757 3655
rect 7791 3652 7803 3655
rect 7926 3652 7932 3664
rect 7791 3624 7932 3652
rect 7791 3621 7803 3624
rect 7745 3615 7803 3621
rect 7926 3612 7932 3624
rect 7984 3652 7990 3664
rect 10045 3655 10103 3661
rect 7984 3624 9076 3652
rect 7984 3612 7990 3624
rect 9048 3593 9076 3624
rect 9140 3624 9536 3652
rect 9140 3596 9168 3624
rect 7653 3587 7711 3593
rect 7653 3584 7665 3587
rect 7576 3556 7665 3584
rect 7653 3553 7665 3556
rect 7699 3553 7711 3587
rect 7845 3587 7903 3593
rect 7845 3584 7857 3587
rect 7653 3547 7711 3553
rect 7760 3556 7857 3584
rect 7760 3528 7788 3556
rect 7845 3553 7857 3556
rect 7891 3553 7903 3587
rect 8021 3587 8079 3593
rect 8021 3584 8033 3587
rect 7845 3547 7903 3553
rect 7944 3556 8033 3584
rect 7742 3476 7748 3528
rect 7800 3476 7806 3528
rect 6638 3408 6644 3460
rect 6696 3448 6702 3460
rect 7944 3448 7972 3556
rect 8021 3553 8033 3556
rect 8067 3553 8079 3587
rect 8021 3547 8079 3553
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3584 8263 3587
rect 8297 3587 8355 3593
rect 8297 3584 8309 3587
rect 8251 3556 8309 3584
rect 8251 3553 8263 3556
rect 8205 3547 8263 3553
rect 8297 3553 8309 3556
rect 8343 3553 8355 3587
rect 8297 3547 8355 3553
rect 9033 3587 9091 3593
rect 9033 3553 9045 3587
rect 9079 3553 9091 3587
rect 9033 3547 9091 3553
rect 9122 3544 9128 3596
rect 9180 3544 9186 3596
rect 9398 3544 9404 3596
rect 9456 3544 9462 3596
rect 9508 3584 9536 3624
rect 10045 3621 10057 3655
rect 10091 3652 10103 3655
rect 10502 3652 10508 3664
rect 10091 3624 10508 3652
rect 10091 3621 10103 3624
rect 10045 3615 10103 3621
rect 10502 3612 10508 3624
rect 10560 3612 10566 3664
rect 10612 3652 10640 3692
rect 11149 3689 11161 3723
rect 11195 3720 11207 3723
rect 11238 3720 11244 3732
rect 11195 3692 11244 3720
rect 11195 3689 11207 3692
rect 11149 3683 11207 3689
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 11882 3680 11888 3732
rect 11940 3680 11946 3732
rect 11900 3652 11928 3680
rect 10612 3624 11928 3652
rect 11090 3587 11148 3593
rect 11090 3584 11102 3587
rect 9508 3556 11102 3584
rect 11090 3553 11102 3556
rect 11136 3553 11148 3587
rect 11090 3547 11148 3553
rect 11330 3544 11336 3596
rect 11388 3584 11394 3596
rect 11517 3587 11575 3593
rect 11517 3584 11529 3587
rect 11388 3556 11529 3584
rect 11388 3544 11394 3556
rect 11517 3553 11529 3556
rect 11563 3553 11575 3587
rect 11517 3547 11575 3553
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 8849 3519 8907 3525
rect 8849 3516 8861 3519
rect 8812 3488 8861 3516
rect 8812 3476 8818 3488
rect 8849 3485 8861 3488
rect 8895 3485 8907 3519
rect 8849 3479 8907 3485
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 9030 3448 9036 3460
rect 6696 3420 9036 3448
rect 6696 3408 6702 3420
rect 9030 3408 9036 3420
rect 9088 3408 9094 3460
rect 11624 3448 11652 3479
rect 9140 3420 11652 3448
rect 7558 3340 7564 3392
rect 7616 3380 7622 3392
rect 8294 3380 8300 3392
rect 7616 3352 8300 3380
rect 7616 3340 7622 3352
rect 8294 3340 8300 3352
rect 8352 3380 8358 3392
rect 9140 3389 9168 3420
rect 9125 3383 9183 3389
rect 9125 3380 9137 3383
rect 8352 3352 9137 3380
rect 8352 3340 8358 3352
rect 9125 3349 9137 3352
rect 9171 3349 9183 3383
rect 9125 3343 9183 3349
rect 10962 3340 10968 3392
rect 11020 3340 11026 3392
rect 552 3290 15364 3312
rect 552 3238 2249 3290
rect 2301 3238 2313 3290
rect 2365 3238 2377 3290
rect 2429 3238 2441 3290
rect 2493 3238 2505 3290
rect 2557 3238 5951 3290
rect 6003 3238 6015 3290
rect 6067 3238 6079 3290
rect 6131 3238 6143 3290
rect 6195 3238 6207 3290
rect 6259 3238 9653 3290
rect 9705 3238 9717 3290
rect 9769 3238 9781 3290
rect 9833 3238 9845 3290
rect 9897 3238 9909 3290
rect 9961 3238 13355 3290
rect 13407 3238 13419 3290
rect 13471 3238 13483 3290
rect 13535 3238 13547 3290
rect 13599 3238 13611 3290
rect 13663 3238 15364 3290
rect 552 3216 15364 3238
rect 7650 3136 7656 3188
rect 7708 3176 7714 3188
rect 8389 3179 8447 3185
rect 8389 3176 8401 3179
rect 7708 3148 8401 3176
rect 7708 3136 7714 3148
rect 8389 3145 8401 3148
rect 8435 3176 8447 3179
rect 8754 3176 8760 3188
rect 8435 3148 8760 3176
rect 8435 3145 8447 3148
rect 8389 3139 8447 3145
rect 8754 3136 8760 3148
rect 8812 3136 8818 3188
rect 11238 3136 11244 3188
rect 11296 3176 11302 3188
rect 11333 3179 11391 3185
rect 11333 3176 11345 3179
rect 11296 3148 11345 3176
rect 11296 3136 11302 3148
rect 11333 3145 11345 3148
rect 11379 3145 11391 3179
rect 11333 3139 11391 3145
rect 4522 3000 4528 3052
rect 4580 3040 4586 3052
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 4580 3012 5457 3040
rect 4580 3000 4586 3012
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3040 7527 3043
rect 7653 3043 7711 3049
rect 7653 3040 7665 3043
rect 7515 3012 7665 3040
rect 7515 3009 7527 3012
rect 7469 3003 7527 3009
rect 7653 3009 7665 3012
rect 7699 3009 7711 3043
rect 7653 3003 7711 3009
rect 7926 3000 7932 3052
rect 7984 3000 7990 3052
rect 11974 3000 11980 3052
rect 12032 3000 12038 3052
rect 6638 2932 6644 2984
rect 6696 2972 6702 2984
rect 7042 2975 7100 2981
rect 7042 2972 7054 2975
rect 6696 2944 7054 2972
rect 6696 2932 6702 2944
rect 7042 2941 7054 2944
rect 7088 2941 7100 2975
rect 7042 2935 7100 2941
rect 7558 2932 7564 2984
rect 7616 2932 7622 2984
rect 8021 2975 8079 2981
rect 8021 2941 8033 2975
rect 8067 2972 8079 2975
rect 8202 2972 8208 2984
rect 8067 2944 8208 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 5712 2907 5770 2913
rect 5712 2873 5724 2907
rect 5758 2904 5770 2907
rect 5902 2904 5908 2916
rect 5758 2876 5908 2904
rect 5758 2873 5770 2876
rect 5712 2867 5770 2873
rect 5902 2864 5908 2876
rect 5960 2864 5966 2916
rect 6840 2876 7144 2904
rect 6840 2845 6868 2876
rect 6825 2839 6883 2845
rect 6825 2805 6837 2839
rect 6871 2805 6883 2839
rect 6825 2799 6883 2805
rect 6914 2796 6920 2848
rect 6972 2796 6978 2848
rect 7116 2845 7144 2876
rect 7101 2839 7159 2845
rect 7101 2805 7113 2839
rect 7147 2836 7159 2839
rect 8036 2836 8064 2935
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 8938 2932 8944 2984
rect 8996 2972 9002 2984
rect 9502 2975 9560 2981
rect 9502 2972 9514 2975
rect 8996 2944 9514 2972
rect 8996 2932 9002 2944
rect 9502 2941 9514 2944
rect 9548 2941 9560 2975
rect 9502 2935 9560 2941
rect 9769 2975 9827 2981
rect 9769 2941 9781 2975
rect 9815 2972 9827 2975
rect 9953 2975 10011 2981
rect 9953 2972 9965 2975
rect 9815 2944 9965 2972
rect 9815 2941 9827 2944
rect 9769 2935 9827 2941
rect 9953 2941 9965 2944
rect 9999 2972 10011 2975
rect 11992 2972 12020 3000
rect 9999 2944 12020 2972
rect 9999 2941 10011 2944
rect 9953 2935 10011 2941
rect 10220 2907 10278 2913
rect 10220 2873 10232 2907
rect 10266 2904 10278 2907
rect 10318 2904 10324 2916
rect 10266 2876 10324 2904
rect 10266 2873 10278 2876
rect 10220 2867 10278 2873
rect 10318 2864 10324 2876
rect 10376 2864 10382 2916
rect 7147 2808 8064 2836
rect 7147 2805 7159 2808
rect 7101 2799 7159 2805
rect 552 2746 15520 2768
rect 552 2694 4100 2746
rect 4152 2694 4164 2746
rect 4216 2694 4228 2746
rect 4280 2694 4292 2746
rect 4344 2694 4356 2746
rect 4408 2694 7802 2746
rect 7854 2694 7866 2746
rect 7918 2694 7930 2746
rect 7982 2694 7994 2746
rect 8046 2694 8058 2746
rect 8110 2694 11504 2746
rect 11556 2694 11568 2746
rect 11620 2694 11632 2746
rect 11684 2694 11696 2746
rect 11748 2694 11760 2746
rect 11812 2694 15206 2746
rect 15258 2694 15270 2746
rect 15322 2694 15334 2746
rect 15386 2694 15398 2746
rect 15450 2694 15462 2746
rect 15514 2694 15520 2746
rect 552 2672 15520 2694
rect 5902 2592 5908 2644
rect 5960 2592 5966 2644
rect 10318 2592 10324 2644
rect 10376 2592 10382 2644
rect 5810 2456 5816 2508
rect 5868 2456 5874 2508
rect 5997 2499 6055 2505
rect 5997 2465 6009 2499
rect 6043 2496 6055 2499
rect 6914 2496 6920 2508
rect 6043 2468 6920 2496
rect 6043 2465 6055 2468
rect 5997 2459 6055 2465
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 10226 2456 10232 2508
rect 10284 2456 10290 2508
rect 10413 2499 10471 2505
rect 10413 2465 10425 2499
rect 10459 2496 10471 2499
rect 10962 2496 10968 2508
rect 10459 2468 10968 2496
rect 10459 2465 10471 2468
rect 10413 2459 10471 2465
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 5828 2428 5856 2456
rect 10244 2428 10272 2456
rect 5828 2400 10272 2428
rect 552 2202 15364 2224
rect 552 2150 2249 2202
rect 2301 2150 2313 2202
rect 2365 2150 2377 2202
rect 2429 2150 2441 2202
rect 2493 2150 2505 2202
rect 2557 2150 5951 2202
rect 6003 2150 6015 2202
rect 6067 2150 6079 2202
rect 6131 2150 6143 2202
rect 6195 2150 6207 2202
rect 6259 2150 9653 2202
rect 9705 2150 9717 2202
rect 9769 2150 9781 2202
rect 9833 2150 9845 2202
rect 9897 2150 9909 2202
rect 9961 2150 13355 2202
rect 13407 2150 13419 2202
rect 13471 2150 13483 2202
rect 13535 2150 13547 2202
rect 13599 2150 13611 2202
rect 13663 2150 15364 2202
rect 552 2128 15364 2150
rect 552 1658 15520 1680
rect 552 1606 4100 1658
rect 4152 1606 4164 1658
rect 4216 1606 4228 1658
rect 4280 1606 4292 1658
rect 4344 1606 4356 1658
rect 4408 1606 7802 1658
rect 7854 1606 7866 1658
rect 7918 1606 7930 1658
rect 7982 1606 7994 1658
rect 8046 1606 8058 1658
rect 8110 1606 11504 1658
rect 11556 1606 11568 1658
rect 11620 1606 11632 1658
rect 11684 1606 11696 1658
rect 11748 1606 11760 1658
rect 11812 1606 15206 1658
rect 15258 1606 15270 1658
rect 15322 1606 15334 1658
rect 15386 1606 15398 1658
rect 15450 1606 15462 1658
rect 15514 1606 15520 1658
rect 552 1584 15520 1606
rect 552 1114 15364 1136
rect 552 1062 2249 1114
rect 2301 1062 2313 1114
rect 2365 1062 2377 1114
rect 2429 1062 2441 1114
rect 2493 1062 2505 1114
rect 2557 1062 5951 1114
rect 6003 1062 6015 1114
rect 6067 1062 6079 1114
rect 6131 1062 6143 1114
rect 6195 1062 6207 1114
rect 6259 1062 9653 1114
rect 9705 1062 9717 1114
rect 9769 1062 9781 1114
rect 9833 1062 9845 1114
rect 9897 1062 9909 1114
rect 9961 1062 13355 1114
rect 13407 1062 13419 1114
rect 13471 1062 13483 1114
rect 13535 1062 13547 1114
rect 13599 1062 13611 1114
rect 13663 1062 15364 1114
rect 552 1040 15364 1062
rect 552 570 15520 592
rect 552 518 4100 570
rect 4152 518 4164 570
rect 4216 518 4228 570
rect 4280 518 4292 570
rect 4344 518 4356 570
rect 4408 518 7802 570
rect 7854 518 7866 570
rect 7918 518 7930 570
rect 7982 518 7994 570
rect 8046 518 8058 570
rect 8110 518 11504 570
rect 11556 518 11568 570
rect 11620 518 11632 570
rect 11684 518 11696 570
rect 11748 518 11760 570
rect 11812 518 15206 570
rect 15258 518 15270 570
rect 15322 518 15334 570
rect 15386 518 15398 570
rect 15450 518 15462 570
rect 15514 518 15520 570
rect 552 496 15520 518
<< via1 >>
rect 2249 15206 2301 15258
rect 2313 15206 2365 15258
rect 2377 15206 2429 15258
rect 2441 15206 2493 15258
rect 2505 15206 2557 15258
rect 5951 15206 6003 15258
rect 6015 15206 6067 15258
rect 6079 15206 6131 15258
rect 6143 15206 6195 15258
rect 6207 15206 6259 15258
rect 9653 15206 9705 15258
rect 9717 15206 9769 15258
rect 9781 15206 9833 15258
rect 9845 15206 9897 15258
rect 9909 15206 9961 15258
rect 13355 15206 13407 15258
rect 13419 15206 13471 15258
rect 13483 15206 13535 15258
rect 13547 15206 13599 15258
rect 13611 15206 13663 15258
rect 4896 15147 4948 15156
rect 4896 15113 4905 15147
rect 4905 15113 4939 15147
rect 4939 15113 4948 15147
rect 4896 15104 4948 15113
rect 10876 15104 10928 15156
rect 5540 15036 5592 15088
rect 848 14900 900 14952
rect 2136 14900 2188 14952
rect 3424 14900 3476 14952
rect 4804 14968 4856 15020
rect 5080 14900 5132 14952
rect 8576 14968 8628 15020
rect 4712 14832 4764 14884
rect 5816 14900 5868 14952
rect 7288 14900 7340 14952
rect 7564 14900 7616 14952
rect 8944 14943 8996 14952
rect 8944 14909 8953 14943
rect 8953 14909 8987 14943
rect 8987 14909 8996 14943
rect 8944 14900 8996 14909
rect 10048 14900 10100 14952
rect 11152 14900 11204 14952
rect 12440 14900 12492 14952
rect 13728 14900 13780 14952
rect 10508 14832 10560 14884
rect 4436 14764 4488 14816
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 4620 14764 4672 14773
rect 5448 14807 5500 14816
rect 5448 14773 5457 14807
rect 5457 14773 5491 14807
rect 5491 14773 5500 14807
rect 5448 14764 5500 14773
rect 6276 14807 6328 14816
rect 6276 14773 6285 14807
rect 6285 14773 6319 14807
rect 6319 14773 6328 14807
rect 6276 14764 6328 14773
rect 7656 14764 7708 14816
rect 8392 14807 8444 14816
rect 8392 14773 8401 14807
rect 8401 14773 8435 14807
rect 8435 14773 8444 14807
rect 8392 14764 8444 14773
rect 9036 14764 9088 14816
rect 10784 14764 10836 14816
rect 11336 14764 11388 14816
rect 12808 14807 12860 14816
rect 12808 14773 12817 14807
rect 12817 14773 12851 14807
rect 12851 14773 12860 14807
rect 12808 14764 12860 14773
rect 14004 14807 14056 14816
rect 14004 14773 14013 14807
rect 14013 14773 14047 14807
rect 14047 14773 14056 14807
rect 14004 14764 14056 14773
rect 4100 14662 4152 14714
rect 4164 14662 4216 14714
rect 4228 14662 4280 14714
rect 4292 14662 4344 14714
rect 4356 14662 4408 14714
rect 7802 14662 7854 14714
rect 7866 14662 7918 14714
rect 7930 14662 7982 14714
rect 7994 14662 8046 14714
rect 8058 14662 8110 14714
rect 11504 14662 11556 14714
rect 11568 14662 11620 14714
rect 11632 14662 11684 14714
rect 11696 14662 11748 14714
rect 11760 14662 11812 14714
rect 15206 14662 15258 14714
rect 15270 14662 15322 14714
rect 15334 14662 15386 14714
rect 15398 14662 15450 14714
rect 15462 14662 15514 14714
rect 7472 14560 7524 14612
rect 4988 14424 5040 14476
rect 5264 14492 5316 14544
rect 5172 14424 5224 14476
rect 4804 14220 4856 14272
rect 5172 14220 5224 14272
rect 5356 14220 5408 14272
rect 6920 14467 6972 14476
rect 6920 14433 6938 14467
rect 6938 14433 6972 14467
rect 6920 14424 6972 14433
rect 7564 14467 7616 14476
rect 7564 14433 7573 14467
rect 7573 14433 7607 14467
rect 7607 14433 7616 14467
rect 7564 14424 7616 14433
rect 8208 14560 8260 14612
rect 8944 14560 8996 14612
rect 14004 14560 14056 14612
rect 9220 14467 9272 14476
rect 9220 14433 9238 14467
rect 9238 14433 9272 14467
rect 9220 14424 9272 14433
rect 12808 14492 12860 14544
rect 12440 14467 12492 14476
rect 12440 14433 12449 14467
rect 12449 14433 12483 14467
rect 12483 14433 12492 14467
rect 12440 14424 12492 14433
rect 8484 14356 8536 14408
rect 9496 14399 9548 14408
rect 9496 14365 9505 14399
rect 9505 14365 9539 14399
rect 9539 14365 9548 14399
rect 9496 14356 9548 14365
rect 10140 14399 10192 14408
rect 10140 14365 10149 14399
rect 10149 14365 10183 14399
rect 10183 14365 10192 14399
rect 10140 14356 10192 14365
rect 10232 14356 10284 14408
rect 11336 14356 11388 14408
rect 7288 14263 7340 14272
rect 7288 14229 7297 14263
rect 7297 14229 7331 14263
rect 7331 14229 7340 14263
rect 7288 14220 7340 14229
rect 7380 14220 7432 14272
rect 9128 14220 9180 14272
rect 10968 14263 11020 14272
rect 10968 14229 10977 14263
rect 10977 14229 11011 14263
rect 11011 14229 11020 14263
rect 10968 14220 11020 14229
rect 14188 14263 14240 14272
rect 14188 14229 14197 14263
rect 14197 14229 14231 14263
rect 14231 14229 14240 14263
rect 14188 14220 14240 14229
rect 2249 14118 2301 14170
rect 2313 14118 2365 14170
rect 2377 14118 2429 14170
rect 2441 14118 2493 14170
rect 2505 14118 2557 14170
rect 5951 14118 6003 14170
rect 6015 14118 6067 14170
rect 6079 14118 6131 14170
rect 6143 14118 6195 14170
rect 6207 14118 6259 14170
rect 9653 14118 9705 14170
rect 9717 14118 9769 14170
rect 9781 14118 9833 14170
rect 9845 14118 9897 14170
rect 9909 14118 9961 14170
rect 13355 14118 13407 14170
rect 13419 14118 13471 14170
rect 13483 14118 13535 14170
rect 13547 14118 13599 14170
rect 13611 14118 13663 14170
rect 4896 14016 4948 14068
rect 4988 14059 5040 14068
rect 4988 14025 4997 14059
rect 4997 14025 5031 14059
rect 5031 14025 5040 14059
rect 4988 14016 5040 14025
rect 6920 14016 6972 14068
rect 9220 14059 9272 14068
rect 9220 14025 9229 14059
rect 9229 14025 9263 14059
rect 9263 14025 9272 14059
rect 9220 14016 9272 14025
rect 10140 14016 10192 14068
rect 10876 14059 10928 14068
rect 10876 14025 10885 14059
rect 10885 14025 10919 14059
rect 10919 14025 10928 14059
rect 10876 14016 10928 14025
rect 11060 14016 11112 14068
rect 12072 14016 12124 14068
rect 13912 14016 13964 14068
rect 6184 13948 6236 14000
rect 4620 13880 4672 13932
rect 4528 13812 4580 13864
rect 5172 13880 5224 13932
rect 8760 13948 8812 14000
rect 7288 13880 7340 13932
rect 8392 13880 8444 13932
rect 7656 13812 7708 13864
rect 8852 13812 8904 13864
rect 10784 13948 10836 14000
rect 12900 13991 12952 14000
rect 12900 13957 12909 13991
rect 12909 13957 12943 13991
rect 12943 13957 12952 13991
rect 12900 13948 12952 13957
rect 10232 13812 10284 13864
rect 10968 13855 11020 13864
rect 10968 13821 10971 13855
rect 10971 13821 11005 13855
rect 11005 13821 11020 13855
rect 10968 13812 11020 13821
rect 5448 13744 5500 13796
rect 11428 13744 11480 13796
rect 14188 13880 14240 13932
rect 11888 13855 11940 13864
rect 11888 13821 11897 13855
rect 11897 13821 11931 13855
rect 11931 13821 11940 13855
rect 11888 13812 11940 13821
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 12164 13855 12216 13864
rect 12164 13821 12173 13855
rect 12173 13821 12207 13855
rect 12207 13821 12216 13855
rect 12164 13812 12216 13821
rect 12348 13855 12400 13864
rect 12348 13821 12357 13855
rect 12357 13821 12391 13855
rect 12391 13821 12400 13855
rect 12348 13812 12400 13821
rect 12624 13855 12676 13864
rect 12624 13821 12633 13855
rect 12633 13821 12667 13855
rect 12667 13821 12676 13855
rect 12624 13812 12676 13821
rect 14464 13855 14516 13864
rect 14464 13821 14473 13855
rect 14473 13821 14507 13855
rect 14507 13821 14516 13855
rect 14464 13812 14516 13821
rect 15108 13812 15160 13864
rect 6184 13676 6236 13728
rect 7380 13676 7432 13728
rect 7656 13676 7708 13728
rect 12992 13744 13044 13796
rect 12256 13719 12308 13728
rect 12256 13685 12265 13719
rect 12265 13685 12299 13719
rect 12299 13685 12308 13719
rect 12256 13676 12308 13685
rect 12808 13676 12860 13728
rect 14648 13719 14700 13728
rect 14648 13685 14657 13719
rect 14657 13685 14691 13719
rect 14691 13685 14700 13719
rect 14648 13676 14700 13685
rect 4100 13574 4152 13626
rect 4164 13574 4216 13626
rect 4228 13574 4280 13626
rect 4292 13574 4344 13626
rect 4356 13574 4408 13626
rect 7802 13574 7854 13626
rect 7866 13574 7918 13626
rect 7930 13574 7982 13626
rect 7994 13574 8046 13626
rect 8058 13574 8110 13626
rect 11504 13574 11556 13626
rect 11568 13574 11620 13626
rect 11632 13574 11684 13626
rect 11696 13574 11748 13626
rect 11760 13574 11812 13626
rect 15206 13574 15258 13626
rect 15270 13574 15322 13626
rect 15334 13574 15386 13626
rect 15398 13574 15450 13626
rect 15462 13574 15514 13626
rect 11888 13472 11940 13524
rect 12256 13472 12308 13524
rect 12440 13472 12492 13524
rect 12624 13472 12676 13524
rect 15108 13472 15160 13524
rect 4528 13336 4580 13388
rect 4160 13268 4212 13320
rect 12072 13404 12124 13456
rect 6276 13268 6328 13320
rect 8668 13336 8720 13388
rect 9312 13379 9364 13388
rect 9312 13345 9346 13379
rect 9346 13345 9364 13379
rect 9312 13336 9364 13345
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 8576 13311 8628 13320
rect 8576 13277 8585 13311
rect 8585 13277 8619 13311
rect 8619 13277 8628 13311
rect 8576 13268 8628 13277
rect 4344 13200 4396 13252
rect 4528 13175 4580 13184
rect 4528 13141 4537 13175
rect 4537 13141 4571 13175
rect 4571 13141 4580 13175
rect 4528 13132 4580 13141
rect 5816 13175 5868 13184
rect 5816 13141 5825 13175
rect 5825 13141 5859 13175
rect 5859 13141 5868 13175
rect 5816 13132 5868 13141
rect 7380 13132 7432 13184
rect 11796 13379 11848 13388
rect 11796 13345 11805 13379
rect 11805 13345 11839 13379
rect 11839 13345 11848 13379
rect 11796 13336 11848 13345
rect 11888 13379 11940 13388
rect 11888 13345 11897 13379
rect 11897 13345 11931 13379
rect 11931 13345 11940 13379
rect 11888 13336 11940 13345
rect 13268 13404 13320 13456
rect 12348 13336 12400 13388
rect 12808 13336 12860 13388
rect 12900 13336 12952 13388
rect 11244 13268 11296 13320
rect 10416 13175 10468 13184
rect 10416 13141 10425 13175
rect 10425 13141 10459 13175
rect 10459 13141 10468 13175
rect 10416 13132 10468 13141
rect 12532 13175 12584 13184
rect 12532 13141 12541 13175
rect 12541 13141 12575 13175
rect 12575 13141 12584 13175
rect 12532 13132 12584 13141
rect 2249 13030 2301 13082
rect 2313 13030 2365 13082
rect 2377 13030 2429 13082
rect 2441 13030 2493 13082
rect 2505 13030 2557 13082
rect 5951 13030 6003 13082
rect 6015 13030 6067 13082
rect 6079 13030 6131 13082
rect 6143 13030 6195 13082
rect 6207 13030 6259 13082
rect 9653 13030 9705 13082
rect 9717 13030 9769 13082
rect 9781 13030 9833 13082
rect 9845 13030 9897 13082
rect 9909 13030 9961 13082
rect 13355 13030 13407 13082
rect 13419 13030 13471 13082
rect 13483 13030 13535 13082
rect 13547 13030 13599 13082
rect 13611 13030 13663 13082
rect 6460 12928 6512 12980
rect 7288 12928 7340 12980
rect 7564 12928 7616 12980
rect 7656 12928 7708 12980
rect 8668 12928 8720 12980
rect 9312 12928 9364 12980
rect 10692 12928 10744 12980
rect 11060 12928 11112 12980
rect 11796 12928 11848 12980
rect 5264 12835 5316 12844
rect 5264 12801 5273 12835
rect 5273 12801 5307 12835
rect 5307 12801 5316 12835
rect 5264 12792 5316 12801
rect 4528 12724 4580 12776
rect 5816 12724 5868 12776
rect 7380 12792 7432 12844
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 10232 12835 10284 12844
rect 8760 12792 8812 12801
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 9036 12724 9088 12776
rect 3240 12631 3292 12640
rect 3240 12597 3249 12631
rect 3249 12597 3283 12631
rect 3283 12597 3292 12631
rect 3240 12588 3292 12597
rect 6920 12588 6972 12640
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 10416 12724 10468 12776
rect 10508 12588 10560 12640
rect 11244 12588 11296 12640
rect 11428 12724 11480 12776
rect 11888 12792 11940 12844
rect 12624 12860 12676 12912
rect 12348 12792 12400 12844
rect 12900 12860 12952 12912
rect 12256 12656 12308 12708
rect 11980 12588 12032 12640
rect 12624 12656 12676 12708
rect 12900 12656 12952 12708
rect 13912 12767 13964 12776
rect 13912 12733 13921 12767
rect 13921 12733 13955 12767
rect 13955 12733 13964 12767
rect 13912 12724 13964 12733
rect 14188 12767 14240 12776
rect 14188 12733 14197 12767
rect 14197 12733 14231 12767
rect 14231 12733 14240 12767
rect 14188 12724 14240 12733
rect 14648 12724 14700 12776
rect 15108 12724 15160 12776
rect 13636 12588 13688 12640
rect 4100 12486 4152 12538
rect 4164 12486 4216 12538
rect 4228 12486 4280 12538
rect 4292 12486 4344 12538
rect 4356 12486 4408 12538
rect 7802 12486 7854 12538
rect 7866 12486 7918 12538
rect 7930 12486 7982 12538
rect 7994 12486 8046 12538
rect 8058 12486 8110 12538
rect 11504 12486 11556 12538
rect 11568 12486 11620 12538
rect 11632 12486 11684 12538
rect 11696 12486 11748 12538
rect 11760 12486 11812 12538
rect 15206 12486 15258 12538
rect 15270 12486 15322 12538
rect 15334 12486 15386 12538
rect 15398 12486 15450 12538
rect 15462 12486 15514 12538
rect 4436 12384 4488 12436
rect 8852 12384 8904 12436
rect 11888 12384 11940 12436
rect 11980 12384 12032 12436
rect 12532 12384 12584 12436
rect 5356 12316 5408 12368
rect 7012 12248 7064 12300
rect 8116 12291 8168 12300
rect 8116 12257 8125 12291
rect 8125 12257 8159 12291
rect 8159 12257 8168 12291
rect 8116 12248 8168 12257
rect 8208 12291 8260 12300
rect 8208 12257 8217 12291
rect 8217 12257 8251 12291
rect 8251 12257 8260 12291
rect 8208 12248 8260 12257
rect 15108 12316 15160 12368
rect 13268 12248 13320 12300
rect 13636 12291 13688 12300
rect 13636 12257 13645 12291
rect 13645 12257 13679 12291
rect 13679 12257 13688 12291
rect 13636 12248 13688 12257
rect 7380 12180 7432 12232
rect 8576 12180 8628 12232
rect 8852 12180 8904 12232
rect 11428 12180 11480 12232
rect 12256 12223 12308 12232
rect 12256 12189 12265 12223
rect 12265 12189 12299 12223
rect 12299 12189 12308 12223
rect 12256 12180 12308 12189
rect 8668 12112 8720 12164
rect 8760 12155 8812 12164
rect 8760 12121 8769 12155
rect 8769 12121 8803 12155
rect 8803 12121 8812 12155
rect 8760 12112 8812 12121
rect 9128 12112 9180 12164
rect 10416 12112 10468 12164
rect 3884 12044 3936 12096
rect 3976 12044 4028 12096
rect 4896 12044 4948 12096
rect 8392 12087 8444 12096
rect 8392 12053 8401 12087
rect 8401 12053 8435 12087
rect 8435 12053 8444 12087
rect 8392 12044 8444 12053
rect 9220 12044 9272 12096
rect 9404 12044 9456 12096
rect 2249 11942 2301 11994
rect 2313 11942 2365 11994
rect 2377 11942 2429 11994
rect 2441 11942 2493 11994
rect 2505 11942 2557 11994
rect 5951 11942 6003 11994
rect 6015 11942 6067 11994
rect 6079 11942 6131 11994
rect 6143 11942 6195 11994
rect 6207 11942 6259 11994
rect 9653 11942 9705 11994
rect 9717 11942 9769 11994
rect 9781 11942 9833 11994
rect 9845 11942 9897 11994
rect 9909 11942 9961 11994
rect 13355 11942 13407 11994
rect 13419 11942 13471 11994
rect 13483 11942 13535 11994
rect 13547 11942 13599 11994
rect 13611 11942 13663 11994
rect 6920 11772 6972 11824
rect 3240 11704 3292 11756
rect 3884 11747 3936 11756
rect 3884 11713 3893 11747
rect 3893 11713 3927 11747
rect 3927 11713 3936 11747
rect 3884 11704 3936 11713
rect 4988 11704 5040 11756
rect 3976 11679 4028 11688
rect 3976 11645 3985 11679
rect 3985 11645 4019 11679
rect 4019 11645 4028 11679
rect 3976 11636 4028 11645
rect 4620 11636 4672 11688
rect 5356 11679 5408 11688
rect 5356 11645 5365 11679
rect 5365 11645 5399 11679
rect 5399 11645 5408 11679
rect 5356 11636 5408 11645
rect 5632 11568 5684 11620
rect 6276 11611 6328 11620
rect 6276 11577 6285 11611
rect 6285 11577 6319 11611
rect 6319 11577 6328 11611
rect 6276 11568 6328 11577
rect 5724 11543 5776 11552
rect 5724 11509 5733 11543
rect 5733 11509 5767 11543
rect 5767 11509 5776 11543
rect 5724 11500 5776 11509
rect 6000 11500 6052 11552
rect 7012 11679 7064 11688
rect 7012 11645 7019 11679
rect 7019 11645 7064 11679
rect 7012 11636 7064 11645
rect 7380 11840 7432 11892
rect 8208 11840 8260 11892
rect 8668 11840 8720 11892
rect 9312 11840 9364 11892
rect 7288 11772 7340 11824
rect 8300 11704 8352 11756
rect 7472 11636 7524 11688
rect 8116 11568 8168 11620
rect 9496 11704 9548 11756
rect 12624 11840 12676 11892
rect 12900 11883 12952 11892
rect 12900 11849 12909 11883
rect 12909 11849 12943 11883
rect 12943 11849 12952 11883
rect 12900 11840 12952 11849
rect 9220 11679 9272 11688
rect 9220 11645 9229 11679
rect 9229 11645 9263 11679
rect 9263 11645 9272 11679
rect 9220 11636 9272 11645
rect 9404 11636 9456 11688
rect 7472 11543 7524 11552
rect 7472 11509 7481 11543
rect 7481 11509 7515 11543
rect 7515 11509 7524 11543
rect 7472 11500 7524 11509
rect 7564 11543 7616 11552
rect 7564 11509 7573 11543
rect 7573 11509 7607 11543
rect 7607 11509 7616 11543
rect 7564 11500 7616 11509
rect 7656 11500 7708 11552
rect 8944 11611 8996 11620
rect 8944 11577 8953 11611
rect 8953 11577 8987 11611
rect 8987 11577 8996 11611
rect 8944 11568 8996 11577
rect 9680 11568 9732 11620
rect 11244 11636 11296 11688
rect 8576 11543 8628 11552
rect 8576 11509 8585 11543
rect 8585 11509 8619 11543
rect 8619 11509 8628 11543
rect 8576 11500 8628 11509
rect 13084 11611 13136 11620
rect 13084 11577 13093 11611
rect 13093 11577 13127 11611
rect 13127 11577 13136 11611
rect 13912 11679 13964 11688
rect 13912 11645 13921 11679
rect 13921 11645 13955 11679
rect 13955 11645 13964 11679
rect 13912 11636 13964 11645
rect 14004 11679 14056 11688
rect 14004 11645 14013 11679
rect 14013 11645 14047 11679
rect 14047 11645 14056 11679
rect 14004 11636 14056 11645
rect 14188 11679 14240 11688
rect 14188 11645 14197 11679
rect 14197 11645 14231 11679
rect 14231 11645 14240 11679
rect 14188 11636 14240 11645
rect 13084 11568 13136 11577
rect 11152 11543 11204 11552
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 11152 11500 11204 11509
rect 12440 11500 12492 11552
rect 12900 11543 12952 11552
rect 12900 11509 12927 11543
rect 12927 11509 12952 11543
rect 12900 11500 12952 11509
rect 13636 11500 13688 11552
rect 4100 11398 4152 11450
rect 4164 11398 4216 11450
rect 4228 11398 4280 11450
rect 4292 11398 4344 11450
rect 4356 11398 4408 11450
rect 7802 11398 7854 11450
rect 7866 11398 7918 11450
rect 7930 11398 7982 11450
rect 7994 11398 8046 11450
rect 8058 11398 8110 11450
rect 11504 11398 11556 11450
rect 11568 11398 11620 11450
rect 11632 11398 11684 11450
rect 11696 11398 11748 11450
rect 11760 11398 11812 11450
rect 15206 11398 15258 11450
rect 15270 11398 15322 11450
rect 15334 11398 15386 11450
rect 15398 11398 15450 11450
rect 15462 11398 15514 11450
rect 3976 11296 4028 11348
rect 4620 11296 4672 11348
rect 4344 11203 4396 11212
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 5356 11296 5408 11348
rect 5724 11160 5776 11212
rect 6000 11203 6052 11212
rect 6000 11169 6009 11203
rect 6009 11169 6043 11203
rect 6043 11169 6052 11203
rect 6000 11160 6052 11169
rect 7380 11296 7432 11348
rect 8576 11296 8628 11348
rect 8944 11339 8996 11348
rect 8944 11305 8953 11339
rect 8953 11305 8987 11339
rect 8987 11305 8996 11339
rect 8944 11296 8996 11305
rect 9680 11339 9732 11348
rect 9680 11305 9689 11339
rect 9689 11305 9723 11339
rect 9723 11305 9732 11339
rect 9680 11296 9732 11305
rect 11888 11339 11940 11348
rect 11888 11305 11897 11339
rect 11897 11305 11931 11339
rect 11931 11305 11940 11339
rect 11888 11296 11940 11305
rect 14004 11296 14056 11348
rect 8668 11228 8720 11280
rect 5172 11135 5224 11144
rect 5172 11101 5181 11135
rect 5181 11101 5215 11135
rect 5215 11101 5224 11135
rect 5172 11092 5224 11101
rect 7012 11203 7064 11212
rect 7012 11169 7021 11203
rect 7021 11169 7055 11203
rect 7055 11169 7064 11203
rect 7012 11160 7064 11169
rect 7472 11160 7524 11212
rect 7564 11160 7616 11212
rect 7656 11160 7708 11212
rect 8392 11160 8444 11212
rect 6920 11067 6972 11076
rect 6920 11033 6929 11067
rect 6929 11033 6963 11067
rect 6963 11033 6972 11067
rect 6920 11024 6972 11033
rect 3884 10999 3936 11008
rect 3884 10965 3893 10999
rect 3893 10965 3927 10999
rect 3927 10965 3936 10999
rect 3884 10956 3936 10965
rect 4804 10956 4856 11008
rect 4988 10999 5040 11008
rect 4988 10965 4997 10999
rect 4997 10965 5031 10999
rect 5031 10965 5040 10999
rect 4988 10956 5040 10965
rect 6368 10999 6420 11008
rect 6368 10965 6377 10999
rect 6377 10965 6411 10999
rect 6411 10965 6420 10999
rect 6368 10956 6420 10965
rect 7196 10956 7248 11008
rect 8392 11024 8444 11076
rect 10140 11203 10192 11212
rect 10140 11169 10149 11203
rect 10149 11169 10183 11203
rect 10183 11169 10192 11203
rect 10140 11160 10192 11169
rect 9496 11024 9548 11076
rect 10048 11067 10100 11076
rect 10048 11033 10057 11067
rect 10057 11033 10091 11067
rect 10091 11033 10100 11067
rect 10048 11024 10100 11033
rect 11152 11160 11204 11212
rect 12072 11160 12124 11212
rect 12348 11203 12400 11212
rect 12348 11169 12357 11203
rect 12357 11169 12391 11203
rect 12391 11169 12400 11203
rect 12348 11160 12400 11169
rect 12440 11203 12492 11212
rect 12440 11169 12450 11203
rect 12450 11169 12484 11203
rect 12484 11169 12492 11203
rect 12440 11160 12492 11169
rect 12624 11203 12676 11212
rect 12624 11169 12633 11203
rect 12633 11169 12667 11203
rect 12667 11169 12676 11203
rect 12624 11160 12676 11169
rect 12716 11203 12768 11212
rect 12716 11169 12725 11203
rect 12725 11169 12759 11203
rect 12759 11169 12768 11203
rect 12716 11160 12768 11169
rect 13268 11160 13320 11212
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 11428 11092 11480 11144
rect 13176 11092 13228 11144
rect 13084 11024 13136 11076
rect 15108 11092 15160 11144
rect 8760 10999 8812 11008
rect 8760 10965 8769 10999
rect 8769 10965 8803 10999
rect 8803 10965 8812 10999
rect 8760 10956 8812 10965
rect 9404 10956 9456 11008
rect 10324 10956 10376 11008
rect 12440 10956 12492 11008
rect 15108 10956 15160 11008
rect 2249 10854 2301 10906
rect 2313 10854 2365 10906
rect 2377 10854 2429 10906
rect 2441 10854 2493 10906
rect 2505 10854 2557 10906
rect 5951 10854 6003 10906
rect 6015 10854 6067 10906
rect 6079 10854 6131 10906
rect 6143 10854 6195 10906
rect 6207 10854 6259 10906
rect 9653 10854 9705 10906
rect 9717 10854 9769 10906
rect 9781 10854 9833 10906
rect 9845 10854 9897 10906
rect 9909 10854 9961 10906
rect 13355 10854 13407 10906
rect 13419 10854 13471 10906
rect 13483 10854 13535 10906
rect 13547 10854 13599 10906
rect 13611 10854 13663 10906
rect 5172 10752 5224 10804
rect 5264 10752 5316 10804
rect 10140 10752 10192 10804
rect 12624 10795 12676 10804
rect 12624 10761 12633 10795
rect 12633 10761 12667 10795
rect 12667 10761 12676 10795
rect 12624 10752 12676 10761
rect 4804 10727 4856 10736
rect 4804 10693 4813 10727
rect 4813 10693 4847 10727
rect 4847 10693 4856 10727
rect 4804 10684 4856 10693
rect 8576 10684 8628 10736
rect 4344 10616 4396 10668
rect 8668 10616 8720 10668
rect 12348 10616 12400 10668
rect 9312 10548 9364 10600
rect 10140 10591 10192 10600
rect 10140 10557 10149 10591
rect 10149 10557 10183 10591
rect 10183 10557 10192 10591
rect 10140 10548 10192 10557
rect 13084 10752 13136 10804
rect 13176 10752 13228 10804
rect 12808 10684 12860 10736
rect 12900 10548 12952 10600
rect 13084 10591 13136 10600
rect 13084 10557 13093 10591
rect 13093 10557 13127 10591
rect 13127 10557 13136 10591
rect 13084 10548 13136 10557
rect 8944 10480 8996 10532
rect 12072 10480 12124 10532
rect 13268 10480 13320 10532
rect 6552 10412 6604 10464
rect 10232 10412 10284 10464
rect 12900 10412 12952 10464
rect 13084 10412 13136 10464
rect 4100 10310 4152 10362
rect 4164 10310 4216 10362
rect 4228 10310 4280 10362
rect 4292 10310 4344 10362
rect 4356 10310 4408 10362
rect 7802 10310 7854 10362
rect 7866 10310 7918 10362
rect 7930 10310 7982 10362
rect 7994 10310 8046 10362
rect 8058 10310 8110 10362
rect 11504 10310 11556 10362
rect 11568 10310 11620 10362
rect 11632 10310 11684 10362
rect 11696 10310 11748 10362
rect 11760 10310 11812 10362
rect 15206 10310 15258 10362
rect 15270 10310 15322 10362
rect 15334 10310 15386 10362
rect 15398 10310 15450 10362
rect 15462 10310 15514 10362
rect 5540 10208 5592 10260
rect 6552 10208 6604 10260
rect 7012 10208 7064 10260
rect 7380 10251 7432 10260
rect 7380 10217 7389 10251
rect 7389 10217 7423 10251
rect 7423 10217 7432 10251
rect 7380 10208 7432 10217
rect 7656 10251 7708 10260
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 8576 10251 8628 10260
rect 8576 10217 8585 10251
rect 8585 10217 8619 10251
rect 8619 10217 8628 10251
rect 8576 10208 8628 10217
rect 8668 10208 8720 10260
rect 10876 10208 10928 10260
rect 5632 10140 5684 10192
rect 5816 10072 5868 10124
rect 6276 10072 6328 10124
rect 7564 10140 7616 10192
rect 5448 10004 5500 10056
rect 6920 10004 6972 10056
rect 7748 10115 7800 10124
rect 7748 10081 7757 10115
rect 7757 10081 7791 10115
rect 7791 10081 7800 10115
rect 7748 10072 7800 10081
rect 8484 10115 8536 10124
rect 8484 10081 8493 10115
rect 8493 10081 8527 10115
rect 8527 10081 8536 10115
rect 8484 10072 8536 10081
rect 8668 10072 8720 10124
rect 9404 10115 9456 10124
rect 9404 10081 9413 10115
rect 9413 10081 9447 10115
rect 9447 10081 9456 10115
rect 9404 10072 9456 10081
rect 10140 10140 10192 10192
rect 10232 10140 10284 10192
rect 11152 10140 11204 10192
rect 12164 10140 12216 10192
rect 10324 10072 10376 10124
rect 14096 10208 14148 10260
rect 12440 10115 12492 10124
rect 12440 10081 12449 10115
rect 12449 10081 12483 10115
rect 12483 10081 12492 10115
rect 12440 10072 12492 10081
rect 9312 9936 9364 9988
rect 5172 9868 5224 9920
rect 6644 9868 6696 9920
rect 11060 10004 11112 10056
rect 12808 10115 12860 10124
rect 12808 10081 12817 10115
rect 12817 10081 12851 10115
rect 12851 10081 12860 10115
rect 12808 10072 12860 10081
rect 10140 9936 10192 9988
rect 12808 9936 12860 9988
rect 10048 9911 10100 9920
rect 10048 9877 10057 9911
rect 10057 9877 10091 9911
rect 10091 9877 10100 9911
rect 10048 9868 10100 9877
rect 12440 9868 12492 9920
rect 13176 9936 13228 9988
rect 13452 10072 13504 10124
rect 13360 10047 13412 10056
rect 13360 10013 13369 10047
rect 13369 10013 13403 10047
rect 13403 10013 13412 10047
rect 13360 10004 13412 10013
rect 15108 9868 15160 9920
rect 2249 9766 2301 9818
rect 2313 9766 2365 9818
rect 2377 9766 2429 9818
rect 2441 9766 2493 9818
rect 2505 9766 2557 9818
rect 5951 9766 6003 9818
rect 6015 9766 6067 9818
rect 6079 9766 6131 9818
rect 6143 9766 6195 9818
rect 6207 9766 6259 9818
rect 9653 9766 9705 9818
rect 9717 9766 9769 9818
rect 9781 9766 9833 9818
rect 9845 9766 9897 9818
rect 9909 9766 9961 9818
rect 13355 9766 13407 9818
rect 13419 9766 13471 9818
rect 13483 9766 13535 9818
rect 13547 9766 13599 9818
rect 13611 9766 13663 9818
rect 5264 9664 5316 9716
rect 5816 9664 5868 9716
rect 7564 9707 7616 9716
rect 7564 9673 7573 9707
rect 7573 9673 7607 9707
rect 7607 9673 7616 9707
rect 7564 9664 7616 9673
rect 7748 9707 7800 9716
rect 7748 9673 7757 9707
rect 7757 9673 7791 9707
rect 7791 9673 7800 9707
rect 7748 9664 7800 9673
rect 8484 9664 8536 9716
rect 8576 9707 8628 9716
rect 8576 9673 8585 9707
rect 8585 9673 8619 9707
rect 8619 9673 8628 9707
rect 8576 9664 8628 9673
rect 8668 9664 8720 9716
rect 11244 9664 11296 9716
rect 6276 9639 6328 9648
rect 6276 9605 6285 9639
rect 6285 9605 6319 9639
rect 6319 9605 6328 9639
rect 6276 9596 6328 9605
rect 10876 9596 10928 9648
rect 12624 9596 12676 9648
rect 8576 9528 8628 9580
rect 12072 9528 12124 9580
rect 5172 9503 5224 9512
rect 5172 9469 5206 9503
rect 5206 9469 5224 9503
rect 5172 9460 5224 9469
rect 7012 9503 7064 9512
rect 7012 9469 7021 9503
rect 7021 9469 7055 9503
rect 7055 9469 7064 9503
rect 7012 9460 7064 9469
rect 7288 9460 7340 9512
rect 7380 9503 7432 9512
rect 7380 9469 7389 9503
rect 7389 9469 7423 9503
rect 7423 9469 7432 9503
rect 7380 9460 7432 9469
rect 10140 9460 10192 9512
rect 10784 9503 10836 9512
rect 10784 9469 10793 9503
rect 10793 9469 10827 9503
rect 10827 9469 10836 9503
rect 10784 9460 10836 9469
rect 10876 9460 10928 9512
rect 11152 9503 11204 9512
rect 11152 9469 11161 9503
rect 11161 9469 11195 9503
rect 11195 9469 11204 9503
rect 11152 9460 11204 9469
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 12624 9503 12676 9512
rect 12624 9469 12631 9503
rect 12631 9469 12676 9503
rect 12624 9460 12676 9469
rect 13176 9664 13228 9716
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 8300 9392 8352 9444
rect 9036 9392 9088 9444
rect 6460 9324 6512 9376
rect 6920 9324 6972 9376
rect 7472 9324 7524 9376
rect 9128 9324 9180 9376
rect 9404 9324 9456 9376
rect 10876 9324 10928 9376
rect 10968 9367 11020 9376
rect 10968 9333 10977 9367
rect 10977 9333 11011 9367
rect 11011 9333 11020 9367
rect 10968 9324 11020 9333
rect 13176 9503 13228 9512
rect 13176 9469 13185 9503
rect 13185 9469 13219 9503
rect 13219 9469 13228 9503
rect 13176 9460 13228 9469
rect 13912 9503 13964 9512
rect 13912 9469 13921 9503
rect 13921 9469 13955 9503
rect 13955 9469 13964 9503
rect 13912 9460 13964 9469
rect 14096 9460 14148 9512
rect 14924 9460 14976 9512
rect 13176 9324 13228 9376
rect 13636 9324 13688 9376
rect 4100 9222 4152 9274
rect 4164 9222 4216 9274
rect 4228 9222 4280 9274
rect 4292 9222 4344 9274
rect 4356 9222 4408 9274
rect 7802 9222 7854 9274
rect 7866 9222 7918 9274
rect 7930 9222 7982 9274
rect 7994 9222 8046 9274
rect 8058 9222 8110 9274
rect 11504 9222 11556 9274
rect 11568 9222 11620 9274
rect 11632 9222 11684 9274
rect 11696 9222 11748 9274
rect 11760 9222 11812 9274
rect 15206 9222 15258 9274
rect 15270 9222 15322 9274
rect 15334 9222 15386 9274
rect 15398 9222 15450 9274
rect 15462 9222 15514 9274
rect 5264 9120 5316 9172
rect 5448 9120 5500 9172
rect 6460 9052 6512 9104
rect 7104 9120 7156 9172
rect 8208 9120 8260 9172
rect 6552 8984 6604 9036
rect 6920 9052 6972 9104
rect 11520 9120 11572 9172
rect 6276 8891 6328 8900
rect 6276 8857 6285 8891
rect 6285 8857 6319 8891
rect 6319 8857 6328 8891
rect 6276 8848 6328 8857
rect 6644 8848 6696 8900
rect 7472 8984 7524 9036
rect 7564 9027 7616 9036
rect 7564 8993 7573 9027
rect 7573 8993 7607 9027
rect 7607 8993 7616 9027
rect 7564 8984 7616 8993
rect 8576 8984 8628 9036
rect 10968 8984 11020 9036
rect 11704 9120 11756 9172
rect 15016 9120 15068 9172
rect 12164 9052 12216 9104
rect 12624 9052 12676 9104
rect 13268 9052 13320 9104
rect 11980 9027 12032 9036
rect 11980 8993 11989 9027
rect 11989 8993 12023 9027
rect 12023 8993 12032 9027
rect 11980 8984 12032 8993
rect 12532 9027 12584 9036
rect 12532 8993 12541 9027
rect 12541 8993 12575 9027
rect 12575 8993 12584 9027
rect 12532 8984 12584 8993
rect 13636 9027 13688 9036
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 13912 8984 13964 9036
rect 7012 8916 7064 8968
rect 10692 8916 10744 8968
rect 11152 8959 11204 8968
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 11152 8916 11204 8925
rect 11520 8916 11572 8968
rect 11704 8916 11756 8968
rect 5816 8780 5868 8832
rect 6736 8780 6788 8832
rect 8944 8823 8996 8832
rect 8944 8789 8953 8823
rect 8953 8789 8987 8823
rect 8987 8789 8996 8823
rect 8944 8780 8996 8789
rect 11704 8780 11756 8832
rect 11796 8823 11848 8832
rect 11796 8789 11805 8823
rect 11805 8789 11839 8823
rect 11839 8789 11848 8823
rect 11796 8780 11848 8789
rect 15016 8780 15068 8832
rect 2249 8678 2301 8730
rect 2313 8678 2365 8730
rect 2377 8678 2429 8730
rect 2441 8678 2493 8730
rect 2505 8678 2557 8730
rect 5951 8678 6003 8730
rect 6015 8678 6067 8730
rect 6079 8678 6131 8730
rect 6143 8678 6195 8730
rect 6207 8678 6259 8730
rect 9653 8678 9705 8730
rect 9717 8678 9769 8730
rect 9781 8678 9833 8730
rect 9845 8678 9897 8730
rect 9909 8678 9961 8730
rect 13355 8678 13407 8730
rect 13419 8678 13471 8730
rect 13483 8678 13535 8730
rect 13547 8678 13599 8730
rect 13611 8678 13663 8730
rect 6276 8576 6328 8628
rect 6552 8576 6604 8628
rect 7472 8576 7524 8628
rect 6644 8508 6696 8560
rect 7288 8508 7340 8560
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 11980 8619 12032 8628
rect 11980 8585 11989 8619
rect 11989 8585 12023 8619
rect 12023 8585 12032 8619
rect 11980 8576 12032 8585
rect 4528 8415 4580 8424
rect 4528 8381 4537 8415
rect 4537 8381 4571 8415
rect 4571 8381 4580 8415
rect 4528 8372 4580 8381
rect 5816 8372 5868 8424
rect 8668 8440 8720 8492
rect 10876 8508 10928 8560
rect 11428 8508 11480 8560
rect 12808 8576 12860 8628
rect 13176 8576 13228 8628
rect 6368 8372 6420 8424
rect 7196 8372 7248 8424
rect 8300 8372 8352 8424
rect 8576 8415 8628 8424
rect 8576 8381 8593 8415
rect 8593 8381 8628 8415
rect 8576 8372 8628 8381
rect 5356 8236 5408 8288
rect 5908 8236 5960 8288
rect 6092 8236 6144 8288
rect 7380 8236 7432 8288
rect 7472 8236 7524 8288
rect 8668 8347 8720 8356
rect 8668 8313 8677 8347
rect 8677 8313 8711 8347
rect 8711 8313 8720 8347
rect 8668 8304 8720 8313
rect 9128 8415 9180 8424
rect 9128 8381 9137 8415
rect 9137 8381 9171 8415
rect 9171 8381 9180 8415
rect 9128 8372 9180 8381
rect 10784 8415 10836 8424
rect 10784 8381 10793 8415
rect 10793 8381 10827 8415
rect 10827 8381 10836 8415
rect 10784 8372 10836 8381
rect 12532 8440 12584 8492
rect 15016 8440 15068 8492
rect 9680 8304 9732 8356
rect 9036 8279 9088 8288
rect 9036 8245 9045 8279
rect 9045 8245 9079 8279
rect 9079 8245 9088 8279
rect 9036 8236 9088 8245
rect 11428 8236 11480 8288
rect 11704 8372 11756 8424
rect 13912 8372 13964 8424
rect 15108 8372 15160 8424
rect 12624 8236 12676 8288
rect 12808 8236 12860 8288
rect 13176 8236 13228 8288
rect 13636 8236 13688 8288
rect 4100 8134 4152 8186
rect 4164 8134 4216 8186
rect 4228 8134 4280 8186
rect 4292 8134 4344 8186
rect 4356 8134 4408 8186
rect 7802 8134 7854 8186
rect 7866 8134 7918 8186
rect 7930 8134 7982 8186
rect 7994 8134 8046 8186
rect 8058 8134 8110 8186
rect 11504 8134 11556 8186
rect 11568 8134 11620 8186
rect 11632 8134 11684 8186
rect 11696 8134 11748 8186
rect 11760 8134 11812 8186
rect 15206 8134 15258 8186
rect 15270 8134 15322 8186
rect 15334 8134 15386 8186
rect 15398 8134 15450 8186
rect 15462 8134 15514 8186
rect 4528 8032 4580 8084
rect 4988 7939 5040 7948
rect 4988 7905 4997 7939
rect 4997 7905 5031 7939
rect 5031 7905 5040 7939
rect 4988 7896 5040 7905
rect 5356 7939 5408 7948
rect 5356 7905 5365 7939
rect 5365 7905 5399 7939
rect 5399 7905 5408 7939
rect 5356 7896 5408 7905
rect 5724 7896 5776 7948
rect 5908 7964 5960 8016
rect 6736 8007 6788 8016
rect 6736 7973 6745 8007
rect 6745 7973 6779 8007
rect 6779 7973 6788 8007
rect 6736 7964 6788 7973
rect 4528 7692 4580 7744
rect 6092 7939 6144 7948
rect 6092 7905 6101 7939
rect 6101 7905 6135 7939
rect 6135 7905 6144 7939
rect 6092 7896 6144 7905
rect 6368 7939 6420 7948
rect 6368 7905 6377 7939
rect 6377 7905 6411 7939
rect 6411 7905 6420 7939
rect 6368 7896 6420 7905
rect 6460 7939 6512 7948
rect 6460 7905 6469 7939
rect 6469 7905 6503 7939
rect 6503 7905 6512 7939
rect 6460 7896 6512 7905
rect 7564 8032 7616 8084
rect 8392 8032 8444 8084
rect 9036 8032 9088 8084
rect 9680 8075 9732 8084
rect 9680 8041 9689 8075
rect 9689 8041 9723 8075
rect 9723 8041 9732 8075
rect 9680 8032 9732 8041
rect 7012 8007 7064 8016
rect 7012 7973 7021 8007
rect 7021 7973 7055 8007
rect 7055 7973 7064 8007
rect 7012 7964 7064 7973
rect 5724 7760 5776 7812
rect 8852 7896 8904 7948
rect 11244 7964 11296 8016
rect 10416 7896 10468 7948
rect 11428 7939 11480 7948
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 11428 7896 11480 7905
rect 9036 7871 9088 7880
rect 9036 7837 9045 7871
rect 9045 7837 9079 7871
rect 9079 7837 9088 7871
rect 9036 7828 9088 7837
rect 9312 7828 9364 7880
rect 11336 7828 11388 7880
rect 12256 7939 12308 7948
rect 12256 7905 12265 7939
rect 12265 7905 12299 7939
rect 12299 7905 12308 7939
rect 12256 7896 12308 7905
rect 12808 7896 12860 7948
rect 13636 7939 13688 7948
rect 13636 7905 13645 7939
rect 13645 7905 13679 7939
rect 13679 7905 13688 7939
rect 13636 7896 13688 7905
rect 13268 7828 13320 7880
rect 9404 7760 9456 7812
rect 7288 7735 7340 7744
rect 7288 7701 7297 7735
rect 7297 7701 7331 7735
rect 7331 7701 7340 7735
rect 7288 7692 7340 7701
rect 12164 7692 12216 7744
rect 15108 7692 15160 7744
rect 2249 7590 2301 7642
rect 2313 7590 2365 7642
rect 2377 7590 2429 7642
rect 2441 7590 2493 7642
rect 2505 7590 2557 7642
rect 5951 7590 6003 7642
rect 6015 7590 6067 7642
rect 6079 7590 6131 7642
rect 6143 7590 6195 7642
rect 6207 7590 6259 7642
rect 9653 7590 9705 7642
rect 9717 7590 9769 7642
rect 9781 7590 9833 7642
rect 9845 7590 9897 7642
rect 9909 7590 9961 7642
rect 13355 7590 13407 7642
rect 13419 7590 13471 7642
rect 13483 7590 13535 7642
rect 13547 7590 13599 7642
rect 13611 7590 13663 7642
rect 9128 7488 9180 7540
rect 13084 7420 13136 7472
rect 7288 7352 7340 7404
rect 7656 7327 7708 7336
rect 7656 7293 7665 7327
rect 7665 7293 7699 7327
rect 7699 7293 7708 7327
rect 7656 7284 7708 7293
rect 8300 7352 8352 7404
rect 10416 7352 10468 7404
rect 10508 7352 10560 7404
rect 8208 7284 8260 7336
rect 8852 7327 8904 7336
rect 8852 7293 8887 7327
rect 8887 7293 8904 7327
rect 8852 7284 8904 7293
rect 12072 7284 12124 7336
rect 12624 7352 12676 7404
rect 12256 7327 12308 7336
rect 12256 7293 12265 7327
rect 12265 7293 12299 7327
rect 12299 7293 12308 7327
rect 12256 7284 12308 7293
rect 8300 7216 8352 7268
rect 8760 7259 8812 7268
rect 8760 7225 8769 7259
rect 8769 7225 8803 7259
rect 8803 7225 8812 7259
rect 8760 7216 8812 7225
rect 10232 7216 10284 7268
rect 6276 7148 6328 7200
rect 6644 7148 6696 7200
rect 8392 7191 8444 7200
rect 8392 7157 8401 7191
rect 8401 7157 8435 7191
rect 8435 7157 8444 7191
rect 8392 7148 8444 7157
rect 10508 7148 10560 7200
rect 12624 7259 12676 7268
rect 12624 7225 12633 7259
rect 12633 7225 12667 7259
rect 12667 7225 12676 7259
rect 12624 7216 12676 7225
rect 13176 7284 13228 7336
rect 14924 7284 14976 7336
rect 4100 7046 4152 7098
rect 4164 7046 4216 7098
rect 4228 7046 4280 7098
rect 4292 7046 4344 7098
rect 4356 7046 4408 7098
rect 7802 7046 7854 7098
rect 7866 7046 7918 7098
rect 7930 7046 7982 7098
rect 7994 7046 8046 7098
rect 8058 7046 8110 7098
rect 11504 7046 11556 7098
rect 11568 7046 11620 7098
rect 11632 7046 11684 7098
rect 11696 7046 11748 7098
rect 11760 7046 11812 7098
rect 15206 7046 15258 7098
rect 15270 7046 15322 7098
rect 15334 7046 15386 7098
rect 15398 7046 15450 7098
rect 15462 7046 15514 7098
rect 6460 6944 6512 6996
rect 7656 6944 7708 6996
rect 8300 6944 8352 6996
rect 8392 6944 8444 6996
rect 5448 6808 5500 6860
rect 7012 6876 7064 6928
rect 6276 6851 6328 6860
rect 6276 6817 6285 6851
rect 6285 6817 6319 6851
rect 6319 6817 6328 6851
rect 6276 6808 6328 6817
rect 6460 6851 6512 6860
rect 6460 6817 6469 6851
rect 6469 6817 6503 6851
rect 6503 6817 6512 6851
rect 8208 6876 8260 6928
rect 6460 6808 6512 6817
rect 6368 6740 6420 6792
rect 7656 6851 7708 6860
rect 7656 6817 7665 6851
rect 7665 6817 7699 6851
rect 7699 6817 7708 6851
rect 7656 6808 7708 6817
rect 4436 6604 4488 6656
rect 8852 6944 8904 6996
rect 11704 6944 11756 6996
rect 12072 6944 12124 6996
rect 9496 6808 9548 6860
rect 12440 6876 12492 6928
rect 10232 6808 10284 6860
rect 10508 6808 10560 6860
rect 10600 6851 10652 6860
rect 10600 6817 10609 6851
rect 10609 6817 10643 6851
rect 10643 6817 10652 6851
rect 10600 6808 10652 6817
rect 10784 6808 10836 6860
rect 12624 6851 12676 6860
rect 12624 6817 12633 6851
rect 12633 6817 12667 6851
rect 12667 6817 12676 6851
rect 12624 6808 12676 6817
rect 13912 6944 13964 6996
rect 13268 6876 13320 6928
rect 13084 6851 13136 6860
rect 13084 6817 13093 6851
rect 13093 6817 13127 6851
rect 13127 6817 13136 6851
rect 13084 6808 13136 6817
rect 14096 6808 14148 6860
rect 9036 6672 9088 6724
rect 13728 6740 13780 6792
rect 12808 6672 12860 6724
rect 8576 6647 8628 6656
rect 8576 6613 8585 6647
rect 8585 6613 8619 6647
rect 8619 6613 8628 6647
rect 8576 6604 8628 6613
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 13176 6647 13228 6656
rect 13176 6613 13185 6647
rect 13185 6613 13219 6647
rect 13219 6613 13228 6647
rect 13176 6604 13228 6613
rect 14464 6672 14516 6724
rect 15016 6604 15068 6656
rect 2249 6502 2301 6554
rect 2313 6502 2365 6554
rect 2377 6502 2429 6554
rect 2441 6502 2493 6554
rect 2505 6502 2557 6554
rect 5951 6502 6003 6554
rect 6015 6502 6067 6554
rect 6079 6502 6131 6554
rect 6143 6502 6195 6554
rect 6207 6502 6259 6554
rect 9653 6502 9705 6554
rect 9717 6502 9769 6554
rect 9781 6502 9833 6554
rect 9845 6502 9897 6554
rect 9909 6502 9961 6554
rect 13355 6502 13407 6554
rect 13419 6502 13471 6554
rect 13483 6502 13535 6554
rect 13547 6502 13599 6554
rect 13611 6502 13663 6554
rect 6460 6400 6512 6452
rect 9496 6400 9548 6452
rect 10600 6443 10652 6452
rect 10600 6409 10609 6443
rect 10609 6409 10643 6443
rect 10643 6409 10652 6443
rect 10600 6400 10652 6409
rect 7472 6332 7524 6384
rect 7564 6332 7616 6384
rect 13728 6400 13780 6452
rect 4436 6171 4488 6180
rect 4436 6137 4470 6171
rect 4470 6137 4488 6171
rect 4436 6128 4488 6137
rect 7012 6196 7064 6248
rect 6920 6128 6972 6180
rect 11888 6264 11940 6316
rect 4528 6060 4580 6112
rect 7288 6060 7340 6112
rect 8576 6196 8628 6248
rect 12164 6239 12216 6248
rect 12164 6205 12197 6239
rect 12197 6205 12216 6239
rect 8208 6128 8260 6180
rect 10508 6128 10560 6180
rect 10692 6128 10744 6180
rect 12164 6196 12216 6205
rect 12992 6332 13044 6384
rect 11336 6128 11388 6180
rect 11704 6128 11756 6180
rect 7748 6103 7800 6112
rect 7748 6069 7757 6103
rect 7757 6069 7791 6103
rect 7791 6069 7800 6103
rect 7748 6060 7800 6069
rect 10876 6060 10928 6112
rect 11888 6060 11940 6112
rect 12532 6239 12584 6248
rect 12532 6205 12541 6239
rect 12541 6205 12575 6239
rect 12575 6205 12584 6239
rect 12532 6196 12584 6205
rect 12900 6196 12952 6248
rect 13084 6196 13136 6248
rect 13176 6196 13228 6248
rect 13912 6196 13964 6248
rect 4100 5958 4152 6010
rect 4164 5958 4216 6010
rect 4228 5958 4280 6010
rect 4292 5958 4344 6010
rect 4356 5958 4408 6010
rect 7802 5958 7854 6010
rect 7866 5958 7918 6010
rect 7930 5958 7982 6010
rect 7994 5958 8046 6010
rect 8058 5958 8110 6010
rect 11504 5958 11556 6010
rect 11568 5958 11620 6010
rect 11632 5958 11684 6010
rect 11696 5958 11748 6010
rect 11760 5958 11812 6010
rect 15206 5958 15258 6010
rect 15270 5958 15322 6010
rect 15334 5958 15386 6010
rect 15398 5958 15450 6010
rect 15462 5958 15514 6010
rect 10784 5856 10836 5908
rect 11980 5856 12032 5908
rect 8944 5788 8996 5840
rect 5540 5720 5592 5772
rect 7380 5720 7432 5772
rect 8208 5720 8260 5772
rect 8024 5652 8076 5704
rect 12992 5652 13044 5704
rect 13268 5652 13320 5704
rect 4528 5516 4580 5568
rect 6368 5584 6420 5636
rect 6920 5516 6972 5568
rect 8208 5516 8260 5568
rect 10876 5516 10928 5568
rect 12072 5516 12124 5568
rect 14464 5516 14516 5568
rect 2249 5414 2301 5466
rect 2313 5414 2365 5466
rect 2377 5414 2429 5466
rect 2441 5414 2493 5466
rect 2505 5414 2557 5466
rect 5951 5414 6003 5466
rect 6015 5414 6067 5466
rect 6079 5414 6131 5466
rect 6143 5414 6195 5466
rect 6207 5414 6259 5466
rect 9653 5414 9705 5466
rect 9717 5414 9769 5466
rect 9781 5414 9833 5466
rect 9845 5414 9897 5466
rect 9909 5414 9961 5466
rect 13355 5414 13407 5466
rect 13419 5414 13471 5466
rect 13483 5414 13535 5466
rect 13547 5414 13599 5466
rect 13611 5414 13663 5466
rect 5540 5312 5592 5364
rect 8208 5244 8260 5296
rect 11336 5312 11388 5364
rect 12440 5312 12492 5364
rect 6920 5219 6972 5228
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 6920 5176 6972 5185
rect 8024 5176 8076 5228
rect 5632 5108 5684 5160
rect 5816 5151 5868 5160
rect 5816 5117 5825 5151
rect 5825 5117 5859 5151
rect 5859 5117 5868 5151
rect 5816 5108 5868 5117
rect 6000 5151 6052 5160
rect 6000 5117 6009 5151
rect 6009 5117 6043 5151
rect 6043 5117 6052 5151
rect 6000 5108 6052 5117
rect 8300 5108 8352 5160
rect 7748 5040 7800 5092
rect 6552 4972 6604 5024
rect 7288 4972 7340 5024
rect 7472 4972 7524 5024
rect 7656 5015 7708 5024
rect 7656 4981 7665 5015
rect 7665 4981 7699 5015
rect 7699 4981 7708 5015
rect 7656 4972 7708 4981
rect 10416 5151 10468 5160
rect 10416 5117 10425 5151
rect 10425 5117 10459 5151
rect 10459 5117 10468 5151
rect 10416 5108 10468 5117
rect 10600 5219 10652 5228
rect 10600 5185 10609 5219
rect 10609 5185 10643 5219
rect 10643 5185 10652 5219
rect 10600 5176 10652 5185
rect 10692 5108 10744 5160
rect 10784 5151 10836 5160
rect 10784 5117 10793 5151
rect 10793 5117 10827 5151
rect 10827 5117 10836 5151
rect 10784 5108 10836 5117
rect 12072 5219 12124 5228
rect 12072 5185 12081 5219
rect 12081 5185 12115 5219
rect 12115 5185 12124 5219
rect 12072 5176 12124 5185
rect 11888 5151 11940 5160
rect 11888 5117 11897 5151
rect 11897 5117 11931 5151
rect 11931 5117 11940 5151
rect 11888 5108 11940 5117
rect 11244 5040 11296 5092
rect 12348 5151 12400 5160
rect 12348 5117 12357 5151
rect 12357 5117 12391 5151
rect 12391 5117 12400 5151
rect 12348 5108 12400 5117
rect 12440 5108 12492 5160
rect 9956 4972 10008 5024
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 11428 4972 11480 5024
rect 11888 4972 11940 5024
rect 13360 5083 13412 5092
rect 13360 5049 13369 5083
rect 13369 5049 13403 5083
rect 13403 5049 13412 5083
rect 13360 5040 13412 5049
rect 4100 4870 4152 4922
rect 4164 4870 4216 4922
rect 4228 4870 4280 4922
rect 4292 4870 4344 4922
rect 4356 4870 4408 4922
rect 7802 4870 7854 4922
rect 7866 4870 7918 4922
rect 7930 4870 7982 4922
rect 7994 4870 8046 4922
rect 8058 4870 8110 4922
rect 11504 4870 11556 4922
rect 11568 4870 11620 4922
rect 11632 4870 11684 4922
rect 11696 4870 11748 4922
rect 11760 4870 11812 4922
rect 15206 4870 15258 4922
rect 15270 4870 15322 4922
rect 15334 4870 15386 4922
rect 15398 4870 15450 4922
rect 15462 4870 15514 4922
rect 6000 4768 6052 4820
rect 6552 4768 6604 4820
rect 7564 4811 7616 4820
rect 7564 4777 7573 4811
rect 7573 4777 7607 4811
rect 7607 4777 7616 4811
rect 7564 4768 7616 4777
rect 7656 4768 7708 4820
rect 8300 4768 8352 4820
rect 6276 4700 6328 4752
rect 4988 4632 5040 4684
rect 5356 4632 5408 4684
rect 5264 4471 5316 4480
rect 5264 4437 5273 4471
rect 5273 4437 5307 4471
rect 5307 4437 5316 4471
rect 5264 4428 5316 4437
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 6644 4675 6696 4684
rect 6644 4641 6653 4675
rect 6653 4641 6687 4675
rect 6687 4641 6696 4675
rect 6644 4632 6696 4641
rect 7840 4743 7892 4752
rect 7840 4709 7849 4743
rect 7849 4709 7883 4743
rect 7883 4709 7892 4743
rect 7840 4700 7892 4709
rect 7380 4632 7432 4684
rect 7288 4564 7340 4616
rect 7564 4632 7616 4684
rect 7472 4496 7524 4548
rect 7196 4471 7248 4480
rect 7196 4437 7205 4471
rect 7205 4437 7239 4471
rect 7239 4437 7248 4471
rect 7196 4428 7248 4437
rect 7932 4675 7984 4684
rect 7932 4641 7941 4675
rect 7941 4641 7975 4675
rect 7975 4641 7984 4675
rect 7932 4632 7984 4641
rect 10048 4632 10100 4684
rect 10876 4768 10928 4820
rect 11244 4811 11296 4820
rect 11244 4777 11253 4811
rect 11253 4777 11287 4811
rect 11287 4777 11296 4811
rect 11244 4768 11296 4777
rect 11336 4811 11388 4820
rect 11336 4777 11345 4811
rect 11345 4777 11379 4811
rect 11379 4777 11388 4811
rect 11336 4768 11388 4777
rect 12348 4768 12400 4820
rect 13360 4811 13412 4820
rect 13360 4777 13369 4811
rect 13369 4777 13403 4811
rect 13403 4777 13412 4811
rect 13360 4768 13412 4777
rect 11796 4700 11848 4752
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 11336 4632 11388 4684
rect 11428 4632 11480 4684
rect 11980 4675 12032 4684
rect 11980 4641 11989 4675
rect 11989 4641 12023 4675
rect 12023 4641 12032 4675
rect 11980 4632 12032 4641
rect 10692 4496 10744 4548
rect 10784 4496 10836 4548
rect 11520 4539 11572 4548
rect 11520 4505 11529 4539
rect 11529 4505 11563 4539
rect 11563 4505 11572 4539
rect 11520 4496 11572 4505
rect 9496 4428 9548 4480
rect 11244 4428 11296 4480
rect 2249 4326 2301 4378
rect 2313 4326 2365 4378
rect 2377 4326 2429 4378
rect 2441 4326 2493 4378
rect 2505 4326 2557 4378
rect 5951 4326 6003 4378
rect 6015 4326 6067 4378
rect 6079 4326 6131 4378
rect 6143 4326 6195 4378
rect 6207 4326 6259 4378
rect 9653 4326 9705 4378
rect 9717 4326 9769 4378
rect 9781 4326 9833 4378
rect 9845 4326 9897 4378
rect 9909 4326 9961 4378
rect 13355 4326 13407 4378
rect 13419 4326 13471 4378
rect 13483 4326 13535 4378
rect 13547 4326 13599 4378
rect 13611 4326 13663 4378
rect 5356 4224 5408 4276
rect 6276 4224 6328 4276
rect 7472 4224 7524 4276
rect 11336 4224 11388 4276
rect 11796 4224 11848 4276
rect 11888 4224 11940 4276
rect 8760 4156 8812 4208
rect 8944 4199 8996 4208
rect 8944 4165 8953 4199
rect 8953 4165 8987 4199
rect 8987 4165 8996 4199
rect 8944 4156 8996 4165
rect 8116 4088 8168 4140
rect 5264 4020 5316 4072
rect 5724 4020 5776 4072
rect 6644 3952 6696 4004
rect 4528 3884 4580 3936
rect 7932 4020 7984 4072
rect 8208 4020 8260 4072
rect 7656 3952 7708 4004
rect 7840 3952 7892 4004
rect 9220 4063 9272 4072
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 9220 4020 9272 4029
rect 9496 4063 9548 4072
rect 9496 4029 9505 4063
rect 9505 4029 9539 4063
rect 9539 4029 9548 4063
rect 9496 4020 9548 4029
rect 10416 4020 10468 4072
rect 10508 4020 10560 4072
rect 11244 4020 11296 4072
rect 11888 4063 11940 4072
rect 11888 4029 11897 4063
rect 11897 4029 11931 4063
rect 11931 4029 11940 4063
rect 11888 4020 11940 4029
rect 12900 4020 12952 4072
rect 8760 3952 8812 4004
rect 7564 3884 7616 3936
rect 9128 3927 9180 3936
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 9404 3927 9456 3936
rect 9404 3893 9413 3927
rect 9413 3893 9447 3927
rect 9447 3893 9456 3927
rect 9404 3884 9456 3893
rect 11336 3927 11388 3936
rect 11336 3893 11345 3927
rect 11345 3893 11379 3927
rect 11379 3893 11388 3927
rect 11336 3884 11388 3893
rect 4100 3782 4152 3834
rect 4164 3782 4216 3834
rect 4228 3782 4280 3834
rect 4292 3782 4344 3834
rect 4356 3782 4408 3834
rect 7802 3782 7854 3834
rect 7866 3782 7918 3834
rect 7930 3782 7982 3834
rect 7994 3782 8046 3834
rect 8058 3782 8110 3834
rect 11504 3782 11556 3834
rect 11568 3782 11620 3834
rect 11632 3782 11684 3834
rect 11696 3782 11748 3834
rect 11760 3782 11812 3834
rect 15206 3782 15258 3834
rect 15270 3782 15322 3834
rect 15334 3782 15386 3834
rect 15398 3782 15450 3834
rect 15462 3782 15514 3834
rect 7564 3680 7616 3732
rect 9128 3680 9180 3732
rect 9220 3680 9272 3732
rect 10232 3680 10284 3732
rect 7932 3612 7984 3664
rect 7748 3476 7800 3528
rect 6644 3408 6696 3460
rect 9128 3544 9180 3596
rect 9404 3587 9456 3596
rect 9404 3553 9413 3587
rect 9413 3553 9447 3587
rect 9447 3553 9456 3587
rect 9404 3544 9456 3553
rect 10508 3612 10560 3664
rect 11244 3680 11296 3732
rect 11888 3680 11940 3732
rect 11336 3544 11388 3596
rect 8760 3476 8812 3528
rect 9036 3408 9088 3460
rect 7564 3340 7616 3392
rect 8300 3340 8352 3392
rect 10968 3383 11020 3392
rect 10968 3349 10977 3383
rect 10977 3349 11011 3383
rect 11011 3349 11020 3383
rect 10968 3340 11020 3349
rect 2249 3238 2301 3290
rect 2313 3238 2365 3290
rect 2377 3238 2429 3290
rect 2441 3238 2493 3290
rect 2505 3238 2557 3290
rect 5951 3238 6003 3290
rect 6015 3238 6067 3290
rect 6079 3238 6131 3290
rect 6143 3238 6195 3290
rect 6207 3238 6259 3290
rect 9653 3238 9705 3290
rect 9717 3238 9769 3290
rect 9781 3238 9833 3290
rect 9845 3238 9897 3290
rect 9909 3238 9961 3290
rect 13355 3238 13407 3290
rect 13419 3238 13471 3290
rect 13483 3238 13535 3290
rect 13547 3238 13599 3290
rect 13611 3238 13663 3290
rect 7656 3136 7708 3188
rect 8760 3136 8812 3188
rect 11244 3136 11296 3188
rect 4528 3000 4580 3052
rect 7932 3043 7984 3052
rect 7932 3009 7941 3043
rect 7941 3009 7975 3043
rect 7975 3009 7984 3043
rect 7932 3000 7984 3009
rect 11980 3000 12032 3052
rect 6644 2932 6696 2984
rect 7564 2975 7616 2984
rect 7564 2941 7573 2975
rect 7573 2941 7607 2975
rect 7607 2941 7616 2975
rect 7564 2932 7616 2941
rect 5908 2864 5960 2916
rect 6920 2839 6972 2848
rect 6920 2805 6929 2839
rect 6929 2805 6963 2839
rect 6963 2805 6972 2839
rect 6920 2796 6972 2805
rect 8208 2932 8260 2984
rect 8944 2932 8996 2984
rect 10324 2864 10376 2916
rect 4100 2694 4152 2746
rect 4164 2694 4216 2746
rect 4228 2694 4280 2746
rect 4292 2694 4344 2746
rect 4356 2694 4408 2746
rect 7802 2694 7854 2746
rect 7866 2694 7918 2746
rect 7930 2694 7982 2746
rect 7994 2694 8046 2746
rect 8058 2694 8110 2746
rect 11504 2694 11556 2746
rect 11568 2694 11620 2746
rect 11632 2694 11684 2746
rect 11696 2694 11748 2746
rect 11760 2694 11812 2746
rect 15206 2694 15258 2746
rect 15270 2694 15322 2746
rect 15334 2694 15386 2746
rect 15398 2694 15450 2746
rect 15462 2694 15514 2746
rect 5908 2635 5960 2644
rect 5908 2601 5917 2635
rect 5917 2601 5951 2635
rect 5951 2601 5960 2635
rect 5908 2592 5960 2601
rect 10324 2635 10376 2644
rect 10324 2601 10333 2635
rect 10333 2601 10367 2635
rect 10367 2601 10376 2635
rect 10324 2592 10376 2601
rect 5816 2499 5868 2508
rect 5816 2465 5825 2499
rect 5825 2465 5859 2499
rect 5859 2465 5868 2499
rect 5816 2456 5868 2465
rect 6920 2456 6972 2508
rect 10232 2499 10284 2508
rect 10232 2465 10241 2499
rect 10241 2465 10275 2499
rect 10275 2465 10284 2499
rect 10232 2456 10284 2465
rect 10968 2456 11020 2508
rect 2249 2150 2301 2202
rect 2313 2150 2365 2202
rect 2377 2150 2429 2202
rect 2441 2150 2493 2202
rect 2505 2150 2557 2202
rect 5951 2150 6003 2202
rect 6015 2150 6067 2202
rect 6079 2150 6131 2202
rect 6143 2150 6195 2202
rect 6207 2150 6259 2202
rect 9653 2150 9705 2202
rect 9717 2150 9769 2202
rect 9781 2150 9833 2202
rect 9845 2150 9897 2202
rect 9909 2150 9961 2202
rect 13355 2150 13407 2202
rect 13419 2150 13471 2202
rect 13483 2150 13535 2202
rect 13547 2150 13599 2202
rect 13611 2150 13663 2202
rect 4100 1606 4152 1658
rect 4164 1606 4216 1658
rect 4228 1606 4280 1658
rect 4292 1606 4344 1658
rect 4356 1606 4408 1658
rect 7802 1606 7854 1658
rect 7866 1606 7918 1658
rect 7930 1606 7982 1658
rect 7994 1606 8046 1658
rect 8058 1606 8110 1658
rect 11504 1606 11556 1658
rect 11568 1606 11620 1658
rect 11632 1606 11684 1658
rect 11696 1606 11748 1658
rect 11760 1606 11812 1658
rect 15206 1606 15258 1658
rect 15270 1606 15322 1658
rect 15334 1606 15386 1658
rect 15398 1606 15450 1658
rect 15462 1606 15514 1658
rect 2249 1062 2301 1114
rect 2313 1062 2365 1114
rect 2377 1062 2429 1114
rect 2441 1062 2493 1114
rect 2505 1062 2557 1114
rect 5951 1062 6003 1114
rect 6015 1062 6067 1114
rect 6079 1062 6131 1114
rect 6143 1062 6195 1114
rect 6207 1062 6259 1114
rect 9653 1062 9705 1114
rect 9717 1062 9769 1114
rect 9781 1062 9833 1114
rect 9845 1062 9897 1114
rect 9909 1062 9961 1114
rect 13355 1062 13407 1114
rect 13419 1062 13471 1114
rect 13483 1062 13535 1114
rect 13547 1062 13599 1114
rect 13611 1062 13663 1114
rect 4100 518 4152 570
rect 4164 518 4216 570
rect 4228 518 4280 570
rect 4292 518 4344 570
rect 4356 518 4408 570
rect 7802 518 7854 570
rect 7866 518 7918 570
rect 7930 518 7982 570
rect 7994 518 8046 570
rect 8058 518 8110 570
rect 11504 518 11556 570
rect 11568 518 11620 570
rect 11632 518 11684 570
rect 11696 518 11748 570
rect 11760 518 11812 570
rect 15206 518 15258 570
rect 15270 518 15322 570
rect 15334 518 15386 570
rect 15398 518 15450 570
rect 15462 518 15514 570
<< metal2 >>
rect 846 15600 902 16000
rect 2134 15600 2190 16000
rect 3422 15600 3478 16000
rect 4710 15600 4766 16000
rect 5998 15600 6054 16000
rect 7286 15600 7342 16000
rect 8574 15600 8630 16000
rect 9862 15600 9918 16000
rect 11150 15600 11206 16000
rect 12438 15600 12494 16000
rect 13726 15600 13782 16000
rect 15014 15600 15070 16000
rect 860 14958 888 15600
rect 2148 14958 2176 15600
rect 2249 15260 2557 15269
rect 2249 15258 2255 15260
rect 2311 15258 2335 15260
rect 2391 15258 2415 15260
rect 2471 15258 2495 15260
rect 2551 15258 2557 15260
rect 2311 15206 2313 15258
rect 2493 15206 2495 15258
rect 2249 15204 2255 15206
rect 2311 15204 2335 15206
rect 2391 15204 2415 15206
rect 2471 15204 2495 15206
rect 2551 15204 2557 15206
rect 2249 15195 2557 15204
rect 3436 14958 3464 15600
rect 848 14952 900 14958
rect 848 14894 900 14900
rect 2136 14952 2188 14958
rect 2136 14894 2188 14900
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 4724 14890 4752 15600
rect 6012 15450 6040 15600
rect 5828 15422 6040 15450
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4712 14884 4764 14890
rect 4712 14826 4764 14832
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4100 14716 4408 14725
rect 4100 14714 4106 14716
rect 4162 14714 4186 14716
rect 4242 14714 4266 14716
rect 4322 14714 4346 14716
rect 4402 14714 4408 14716
rect 4162 14662 4164 14714
rect 4344 14662 4346 14714
rect 4100 14660 4106 14662
rect 4162 14660 4186 14662
rect 4242 14660 4266 14662
rect 4322 14660 4346 14662
rect 4402 14660 4408 14662
rect 4100 14651 4408 14660
rect 2249 14172 2557 14181
rect 2249 14170 2255 14172
rect 2311 14170 2335 14172
rect 2391 14170 2415 14172
rect 2471 14170 2495 14172
rect 2551 14170 2557 14172
rect 2311 14118 2313 14170
rect 2493 14118 2495 14170
rect 2249 14116 2255 14118
rect 2311 14116 2335 14118
rect 2391 14116 2415 14118
rect 2471 14116 2495 14118
rect 2551 14116 2557 14118
rect 2249 14107 2557 14116
rect 4100 13628 4408 13637
rect 4100 13626 4106 13628
rect 4162 13626 4186 13628
rect 4242 13626 4266 13628
rect 4322 13626 4346 13628
rect 4402 13626 4408 13628
rect 4162 13574 4164 13626
rect 4344 13574 4346 13626
rect 4100 13572 4106 13574
rect 4162 13572 4186 13574
rect 4242 13572 4266 13574
rect 4322 13572 4346 13574
rect 4402 13572 4408 13574
rect 4100 13563 4408 13572
rect 4448 13512 4476 14758
rect 4632 13938 4660 14758
rect 4816 14278 4844 14962
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4528 13864 4580 13870
rect 4528 13806 4580 13812
rect 4356 13484 4476 13512
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 2249 13084 2557 13093
rect 2249 13082 2255 13084
rect 2311 13082 2335 13084
rect 2391 13082 2415 13084
rect 2471 13082 2495 13084
rect 2551 13082 2557 13084
rect 2311 13030 2313 13082
rect 2493 13030 2495 13082
rect 2249 13028 2255 13030
rect 2311 13028 2335 13030
rect 2391 13028 2415 13030
rect 2471 13028 2495 13030
rect 2551 13028 2557 13030
rect 2249 13019 2557 13028
rect 4172 12866 4200 13262
rect 4356 13258 4384 13484
rect 4540 13394 4568 13806
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4172 12838 4476 12866
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 2249 11996 2557 12005
rect 2249 11994 2255 11996
rect 2311 11994 2335 11996
rect 2391 11994 2415 11996
rect 2471 11994 2495 11996
rect 2551 11994 2557 11996
rect 2311 11942 2313 11994
rect 2493 11942 2495 11994
rect 2249 11940 2255 11942
rect 2311 11940 2335 11942
rect 2391 11940 2415 11942
rect 2471 11940 2495 11942
rect 2551 11940 2557 11942
rect 2249 11931 2557 11940
rect 3252 11762 3280 12582
rect 4100 12540 4408 12549
rect 4100 12538 4106 12540
rect 4162 12538 4186 12540
rect 4242 12538 4266 12540
rect 4322 12538 4346 12540
rect 4402 12538 4408 12540
rect 4162 12486 4164 12538
rect 4344 12486 4346 12538
rect 4100 12484 4106 12486
rect 4162 12484 4186 12486
rect 4242 12484 4266 12486
rect 4322 12484 4346 12486
rect 4402 12484 4408 12486
rect 4100 12475 4408 12484
rect 4448 12442 4476 12838
rect 4540 12782 4568 13126
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3896 11762 3924 12038
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3896 11014 3924 11698
rect 3988 11694 4016 12038
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 3988 11354 4016 11630
rect 4100 11452 4408 11461
rect 4100 11450 4106 11452
rect 4162 11450 4186 11452
rect 4242 11450 4266 11452
rect 4322 11450 4346 11452
rect 4402 11450 4408 11452
rect 4162 11398 4164 11450
rect 4344 11398 4346 11450
rect 4100 11396 4106 11398
rect 4162 11396 4186 11398
rect 4242 11396 4266 11398
rect 4322 11396 4346 11398
rect 4402 11396 4408 11398
rect 4100 11387 4408 11396
rect 4632 11354 4660 11630
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 2249 10908 2557 10917
rect 2249 10906 2255 10908
rect 2311 10906 2335 10908
rect 2391 10906 2415 10908
rect 2471 10906 2495 10908
rect 2551 10906 2557 10908
rect 2311 10854 2313 10906
rect 2493 10854 2495 10906
rect 2249 10852 2255 10854
rect 2311 10852 2335 10854
rect 2391 10852 2415 10854
rect 2471 10852 2495 10854
rect 2551 10852 2557 10854
rect 2249 10843 2557 10852
rect 4356 10674 4384 11154
rect 4816 11014 4844 14214
rect 4908 14074 4936 15098
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5080 14952 5132 14958
rect 5132 14912 5212 14940
rect 5080 14894 5132 14900
rect 5184 14482 5212 14912
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5264 14544 5316 14550
rect 5264 14486 5316 14492
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 5000 14074 5028 14418
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 4908 12102 4936 14010
rect 5184 13938 5212 14214
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 5276 12850 5304 14486
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5000 11014 5028 11698
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 4816 10742 4844 10950
rect 5184 10810 5212 11086
rect 5276 10810 5304 12786
rect 5368 12374 5396 14214
rect 5460 13802 5488 14758
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5368 11354 5396 11630
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4100 10364 4408 10373
rect 4100 10362 4106 10364
rect 4162 10362 4186 10364
rect 4242 10362 4266 10364
rect 4322 10362 4346 10364
rect 4402 10362 4408 10364
rect 4162 10310 4164 10362
rect 4344 10310 4346 10362
rect 4100 10308 4106 10310
rect 4162 10308 4186 10310
rect 4242 10308 4266 10310
rect 4322 10308 4346 10310
rect 4402 10308 4408 10310
rect 4100 10299 4408 10308
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 2249 9820 2557 9829
rect 2249 9818 2255 9820
rect 2311 9818 2335 9820
rect 2391 9818 2415 9820
rect 2471 9818 2495 9820
rect 2551 9818 2557 9820
rect 2311 9766 2313 9818
rect 2493 9766 2495 9818
rect 2249 9764 2255 9766
rect 2311 9764 2335 9766
rect 2391 9764 2415 9766
rect 2471 9764 2495 9766
rect 2551 9764 2557 9766
rect 2249 9755 2557 9764
rect 5184 9518 5212 9862
rect 5276 9722 5304 10746
rect 5552 10266 5580 15030
rect 5828 14958 5856 15422
rect 5951 15260 6259 15269
rect 5951 15258 5957 15260
rect 6013 15258 6037 15260
rect 6093 15258 6117 15260
rect 6173 15258 6197 15260
rect 6253 15258 6259 15260
rect 6013 15206 6015 15258
rect 6195 15206 6197 15258
rect 5951 15204 5957 15206
rect 6013 15204 6037 15206
rect 6093 15204 6117 15206
rect 6173 15204 6197 15206
rect 6253 15204 6259 15206
rect 5951 15195 6259 15204
rect 7300 14958 7328 15600
rect 8588 15026 8616 15600
rect 9876 15450 9904 15600
rect 9876 15422 10088 15450
rect 9653 15260 9961 15269
rect 9653 15258 9659 15260
rect 9715 15258 9739 15260
rect 9795 15258 9819 15260
rect 9875 15258 9899 15260
rect 9955 15258 9961 15260
rect 9715 15206 9717 15258
rect 9897 15206 9899 15258
rect 9653 15204 9659 15206
rect 9715 15204 9739 15206
rect 9795 15204 9819 15206
rect 9875 15204 9899 15206
rect 9955 15204 9961 15206
rect 9653 15195 9961 15204
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 10060 14958 10088 15422
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 5951 14172 6259 14181
rect 5951 14170 5957 14172
rect 6013 14170 6037 14172
rect 6093 14170 6117 14172
rect 6173 14170 6197 14172
rect 6253 14170 6259 14172
rect 6013 14118 6015 14170
rect 6195 14118 6197 14170
rect 5951 14116 5957 14118
rect 6013 14116 6037 14118
rect 6093 14116 6117 14118
rect 6173 14116 6197 14118
rect 6253 14116 6259 14118
rect 5951 14107 6259 14116
rect 6184 14000 6236 14006
rect 6184 13942 6236 13948
rect 6196 13734 6224 13942
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6288 13326 6316 14758
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6932 14074 6960 14418
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 7300 13938 7328 14214
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7392 13734 7420 14214
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5828 12782 5856 13126
rect 5951 13084 6259 13093
rect 5951 13082 5957 13084
rect 6013 13082 6037 13084
rect 6093 13082 6117 13084
rect 6173 13082 6197 13084
rect 6253 13082 6259 13084
rect 6013 13030 6015 13082
rect 6195 13030 6197 13082
rect 5951 13028 5957 13030
rect 6013 13028 6037 13030
rect 6093 13028 6117 13030
rect 6173 13028 6197 13030
rect 6253 13028 6259 13030
rect 5951 13019 6259 13028
rect 6472 12986 6500 13262
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 7300 12646 7328 12922
rect 7392 12850 7420 13126
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 5951 11996 6259 12005
rect 5951 11994 5957 11996
rect 6013 11994 6037 11996
rect 6093 11994 6117 11996
rect 6173 11994 6197 11996
rect 6253 11994 6259 11996
rect 6013 11942 6015 11994
rect 6195 11942 6197 11994
rect 5951 11940 5957 11942
rect 6013 11940 6037 11942
rect 6093 11940 6117 11942
rect 6173 11940 6197 11942
rect 6253 11940 6259 11942
rect 5951 11931 6259 11940
rect 6932 11830 6960 12582
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5644 10198 5672 11562
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 5736 11218 5764 11494
rect 6012 11218 6040 11494
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 5951 10908 6259 10917
rect 5951 10906 5957 10908
rect 6013 10906 6037 10908
rect 6093 10906 6117 10908
rect 6173 10906 6197 10908
rect 6253 10906 6259 10908
rect 6013 10854 6015 10906
rect 6195 10854 6197 10906
rect 5951 10852 5957 10854
rect 6013 10852 6037 10854
rect 6093 10852 6117 10854
rect 6173 10852 6197 10854
rect 6253 10852 6259 10854
rect 5951 10843 6259 10852
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 6288 10130 6316 11562
rect 6932 11082 6960 11766
rect 7024 11694 7052 12242
rect 7300 11830 7328 12582
rect 7392 12238 7420 12786
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7392 11898 7420 12174
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7288 11824 7340 11830
rect 7288 11766 7340 11772
rect 7484 11694 7512 14554
rect 7576 14482 7604 14894
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7576 12986 7604 14418
rect 7668 13870 7696 14758
rect 7802 14716 8110 14725
rect 7802 14714 7808 14716
rect 7864 14714 7888 14716
rect 7944 14714 7968 14716
rect 8024 14714 8048 14716
rect 8104 14714 8110 14716
rect 7864 14662 7866 14714
rect 8046 14662 8048 14714
rect 7802 14660 7808 14662
rect 7864 14660 7888 14662
rect 7944 14660 7968 14662
rect 8024 14660 8048 14662
rect 8104 14660 8110 14662
rect 7802 14651 8110 14660
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 12986 7696 13670
rect 7802 13628 8110 13637
rect 7802 13626 7808 13628
rect 7864 13626 7888 13628
rect 7944 13626 7968 13628
rect 8024 13626 8048 13628
rect 8104 13626 8110 13628
rect 7864 13574 7866 13626
rect 8046 13574 8048 13626
rect 7802 13572 7808 13574
rect 7864 13572 7888 13574
rect 7944 13572 7968 13574
rect 8024 13572 8048 13574
rect 8104 13572 8110 13574
rect 7802 13563 8110 13572
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7802 12540 8110 12549
rect 7802 12538 7808 12540
rect 7864 12538 7888 12540
rect 7944 12538 7968 12540
rect 8024 12538 8048 12540
rect 8104 12538 8110 12540
rect 7864 12486 7866 12538
rect 8046 12486 8048 12538
rect 7802 12484 7808 12486
rect 7864 12484 7888 12486
rect 7944 12484 7968 12486
rect 8024 12484 8048 12486
rect 8104 12484 8110 12486
rect 7802 12475 8110 12484
rect 8220 12306 8248 14554
rect 8404 13938 8432 14758
rect 8956 14618 8984 14894
rect 10508 14884 10560 14890
rect 10508 14826 10560 14832
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8496 13954 8524 14350
rect 8760 14000 8812 14006
rect 8392 13932 8444 13938
rect 8496 13926 8616 13954
rect 8760 13942 8812 13948
rect 8392 13874 8444 13880
rect 8588 13326 8616 13926
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8680 12986 8708 13330
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8772 12850 8800 13942
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8864 12442 8892 13806
rect 9048 12782 9076 14758
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 7012 11688 7064 11694
rect 7472 11688 7524 11694
rect 7064 11648 7144 11676
rect 7012 11630 7064 11636
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 4100 9276 4408 9285
rect 4100 9274 4106 9276
rect 4162 9274 4186 9276
rect 4242 9274 4266 9276
rect 4322 9274 4346 9276
rect 4402 9274 4408 9276
rect 4162 9222 4164 9274
rect 4344 9222 4346 9274
rect 4100 9220 4106 9222
rect 4162 9220 4186 9222
rect 4242 9220 4266 9222
rect 4322 9220 4346 9222
rect 4402 9220 4408 9222
rect 4100 9211 4408 9220
rect 5276 9178 5304 9658
rect 5460 9178 5488 9998
rect 5828 9722 5856 10066
rect 5951 9820 6259 9829
rect 5951 9818 5957 9820
rect 6013 9818 6037 9820
rect 6093 9818 6117 9820
rect 6173 9818 6197 9820
rect 6253 9818 6259 9820
rect 6013 9766 6015 9818
rect 6195 9766 6197 9818
rect 5951 9764 5957 9766
rect 6013 9764 6037 9766
rect 6093 9764 6117 9766
rect 6173 9764 6197 9766
rect 6253 9764 6259 9766
rect 5951 9755 6259 9764
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 6288 9654 6316 10066
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 2249 8732 2557 8741
rect 2249 8730 2255 8732
rect 2311 8730 2335 8732
rect 2391 8730 2415 8732
rect 2471 8730 2495 8732
rect 2551 8730 2557 8732
rect 2311 8678 2313 8730
rect 2493 8678 2495 8730
rect 2249 8676 2255 8678
rect 2311 8676 2335 8678
rect 2391 8676 2415 8678
rect 2471 8676 2495 8678
rect 2551 8676 2557 8678
rect 2249 8667 2557 8676
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4100 8188 4408 8197
rect 4100 8186 4106 8188
rect 4162 8186 4186 8188
rect 4242 8186 4266 8188
rect 4322 8186 4346 8188
rect 4402 8186 4408 8188
rect 4162 8134 4164 8186
rect 4344 8134 4346 8186
rect 4100 8132 4106 8134
rect 4162 8132 4186 8134
rect 4242 8132 4266 8134
rect 4322 8132 4346 8134
rect 4402 8132 4408 8134
rect 4100 8123 4408 8132
rect 4540 8090 4568 8366
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 5368 7954 5396 8230
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 2249 7644 2557 7653
rect 2249 7642 2255 7644
rect 2311 7642 2335 7644
rect 2391 7642 2415 7644
rect 2471 7642 2495 7644
rect 2551 7642 2557 7644
rect 2311 7590 2313 7642
rect 2493 7590 2495 7642
rect 2249 7588 2255 7590
rect 2311 7588 2335 7590
rect 2391 7588 2415 7590
rect 2471 7588 2495 7590
rect 2551 7588 2557 7590
rect 2249 7579 2557 7588
rect 4100 7100 4408 7109
rect 4100 7098 4106 7100
rect 4162 7098 4186 7100
rect 4242 7098 4266 7100
rect 4322 7098 4346 7100
rect 4402 7098 4408 7100
rect 4162 7046 4164 7098
rect 4344 7046 4346 7098
rect 4100 7044 4106 7046
rect 4162 7044 4186 7046
rect 4242 7044 4266 7046
rect 4322 7044 4346 7046
rect 4402 7044 4408 7046
rect 4100 7035 4408 7044
rect 4436 6656 4488 6662
rect 4436 6598 4488 6604
rect 2249 6556 2557 6565
rect 2249 6554 2255 6556
rect 2311 6554 2335 6556
rect 2391 6554 2415 6556
rect 2471 6554 2495 6556
rect 2551 6554 2557 6556
rect 2311 6502 2313 6554
rect 2493 6502 2495 6554
rect 2249 6500 2255 6502
rect 2311 6500 2335 6502
rect 2391 6500 2415 6502
rect 2471 6500 2495 6502
rect 2551 6500 2557 6502
rect 2249 6491 2557 6500
rect 4448 6186 4476 6598
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 4540 6118 4568 7686
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4100 6012 4408 6021
rect 4100 6010 4106 6012
rect 4162 6010 4186 6012
rect 4242 6010 4266 6012
rect 4322 6010 4346 6012
rect 4402 6010 4408 6012
rect 4162 5958 4164 6010
rect 4344 5958 4346 6010
rect 4100 5956 4106 5958
rect 4162 5956 4186 5958
rect 4242 5956 4266 5958
rect 4322 5956 4346 5958
rect 4402 5956 4408 5958
rect 4100 5947 4408 5956
rect 4540 5574 4568 6054
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 2249 5468 2557 5477
rect 2249 5466 2255 5468
rect 2311 5466 2335 5468
rect 2391 5466 2415 5468
rect 2471 5466 2495 5468
rect 2551 5466 2557 5468
rect 2311 5414 2313 5466
rect 2493 5414 2495 5466
rect 2249 5412 2255 5414
rect 2311 5412 2335 5414
rect 2391 5412 2415 5414
rect 2471 5412 2495 5414
rect 2551 5412 2557 5414
rect 2249 5403 2557 5412
rect 4100 4924 4408 4933
rect 4100 4922 4106 4924
rect 4162 4922 4186 4924
rect 4242 4922 4266 4924
rect 4322 4922 4346 4924
rect 4402 4922 4408 4924
rect 4162 4870 4164 4922
rect 4344 4870 4346 4922
rect 4100 4868 4106 4870
rect 4162 4868 4186 4870
rect 4242 4868 4266 4870
rect 4322 4868 4346 4870
rect 4402 4868 4408 4870
rect 4100 4859 4408 4868
rect 2249 4380 2557 4389
rect 2249 4378 2255 4380
rect 2311 4378 2335 4380
rect 2391 4378 2415 4380
rect 2471 4378 2495 4380
rect 2551 4378 2557 4380
rect 2311 4326 2313 4378
rect 2493 4326 2495 4378
rect 2249 4324 2255 4326
rect 2311 4324 2335 4326
rect 2391 4324 2415 4326
rect 2471 4324 2495 4326
rect 2551 4324 2557 4326
rect 2249 4315 2557 4324
rect 4540 3942 4568 5510
rect 5000 4690 5028 7890
rect 5460 6866 5488 9114
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8430 5856 8774
rect 5951 8732 6259 8741
rect 5951 8730 5957 8732
rect 6013 8730 6037 8732
rect 6093 8730 6117 8732
rect 6173 8730 6197 8732
rect 6253 8730 6259 8732
rect 6013 8678 6015 8730
rect 6195 8678 6197 8730
rect 5951 8676 5957 8678
rect 6013 8676 6037 8678
rect 6093 8676 6117 8678
rect 6173 8676 6197 8678
rect 6253 8676 6259 8678
rect 5951 8667 6259 8676
rect 6288 8634 6316 8842
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6380 8430 6408 10950
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6564 10266 6592 10406
rect 7024 10266 7052 11154
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6472 9110 6500 9318
rect 6460 9104 6512 9110
rect 6460 9046 6512 9052
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 6092 8288 6144 8294
rect 6472 8242 6500 9046
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6564 8634 6592 8978
rect 6656 8906 6684 9862
rect 6932 9382 6960 9998
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 9110 6960 9318
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 7024 8974 7052 9454
rect 7116 9178 7144 11648
rect 7392 11648 7472 11676
rect 7392 11354 7420 11648
rect 7472 11630 7524 11636
rect 8128 11642 8156 12242
rect 8220 11898 8248 12242
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8128 11626 8248 11642
rect 8116 11620 8248 11626
rect 8168 11614 8248 11620
rect 8116 11562 8168 11568
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7484 11218 7512 11494
rect 7576 11218 7604 11494
rect 7668 11218 7696 11494
rect 7802 11452 8110 11461
rect 7802 11450 7808 11452
rect 7864 11450 7888 11452
rect 7944 11450 7968 11452
rect 8024 11450 8048 11452
rect 8104 11450 8110 11452
rect 7864 11398 7866 11450
rect 8046 11398 8048 11450
rect 7802 11396 7808 11398
rect 7864 11396 7888 11398
rect 7944 11396 7968 11398
rect 8024 11396 8048 11398
rect 8104 11396 8110 11398
rect 7802 11387 8110 11396
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 6644 8900 6696 8906
rect 6644 8842 6696 8848
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6656 8566 6684 8842
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6092 8230 6144 8236
rect 5920 8022 5948 8230
rect 5908 8016 5960 8022
rect 5908 7958 5960 7964
rect 6104 7954 6132 8230
rect 6380 8214 6500 8242
rect 6380 7954 6408 8214
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 5736 7818 5764 7890
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5448 6860 5500 6866
rect 5500 6820 5672 6848
rect 5448 6802 5500 6808
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5552 5370 5580 5714
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5644 5166 5672 6820
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5276 4078 5304 4422
rect 5368 4282 5396 4626
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5736 4078 5764 7754
rect 5951 7644 6259 7653
rect 5951 7642 5957 7644
rect 6013 7642 6037 7644
rect 6093 7642 6117 7644
rect 6173 7642 6197 7644
rect 6253 7642 6259 7644
rect 6013 7590 6015 7642
rect 6195 7590 6197 7642
rect 5951 7588 5957 7590
rect 6013 7588 6037 7590
rect 6093 7588 6117 7590
rect 6173 7588 6197 7590
rect 6253 7588 6259 7590
rect 5951 7579 6259 7588
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6288 6866 6316 7142
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6380 6798 6408 7890
rect 6472 7002 6500 7890
rect 6656 7206 6684 8502
rect 6748 8022 6776 8774
rect 7208 8430 7236 10950
rect 7668 10266 7696 11154
rect 7802 10364 8110 10373
rect 7802 10362 7808 10364
rect 7864 10362 7888 10364
rect 7944 10362 7968 10364
rect 8024 10362 8048 10364
rect 8104 10362 8110 10364
rect 7864 10310 7866 10362
rect 8046 10310 8048 10362
rect 7802 10308 7808 10310
rect 7864 10308 7888 10310
rect 7944 10308 7968 10310
rect 8024 10308 8048 10310
rect 8104 10308 8110 10310
rect 7802 10299 8110 10308
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7392 9518 7420 10202
rect 7564 10192 7616 10198
rect 7564 10134 7616 10140
rect 7576 9722 7604 10134
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7760 9722 7788 10066
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7300 8566 7328 9454
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7484 9042 7512 9318
rect 7802 9276 8110 9285
rect 7802 9274 7808 9276
rect 7864 9274 7888 9276
rect 7944 9274 7968 9276
rect 8024 9274 8048 9276
rect 8104 9274 8110 9276
rect 7864 9222 7866 9274
rect 8046 9222 8048 9274
rect 7802 9220 7808 9222
rect 7864 9220 7888 9222
rect 7944 9220 7968 9222
rect 8024 9220 8048 9222
rect 8104 9220 8110 9222
rect 7802 9211 8110 9220
rect 8220 9178 8248 11614
rect 8312 9450 8340 11698
rect 8404 11218 8432 12038
rect 8588 11642 8616 12174
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8680 11898 8708 12106
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8588 11614 8708 11642
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8588 11354 8616 11494
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8680 11286 8708 11614
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7484 8634 7512 8978
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7484 8294 7512 8570
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 5951 6556 6259 6565
rect 5951 6554 5957 6556
rect 6013 6554 6037 6556
rect 6093 6554 6117 6556
rect 6173 6554 6197 6556
rect 6253 6554 6259 6556
rect 6013 6502 6015 6554
rect 6195 6502 6197 6554
rect 5951 6500 5957 6502
rect 6013 6500 6037 6502
rect 6093 6500 6117 6502
rect 6173 6500 6197 6502
rect 6253 6500 6259 6502
rect 5951 6491 6259 6500
rect 6380 5642 6408 6734
rect 6472 6458 6500 6802
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 5951 5468 6259 5477
rect 5951 5466 5957 5468
rect 6013 5466 6037 5468
rect 6093 5466 6117 5468
rect 6173 5466 6197 5468
rect 6253 5466 6259 5468
rect 6013 5414 6015 5466
rect 6195 5414 6197 5466
rect 5951 5412 5957 5414
rect 6013 5412 6037 5414
rect 6093 5412 6117 5414
rect 6173 5412 6197 5414
rect 6253 5412 6259 5414
rect 5951 5403 6259 5412
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4100 3836 4408 3845
rect 4100 3834 4106 3836
rect 4162 3834 4186 3836
rect 4242 3834 4266 3836
rect 4322 3834 4346 3836
rect 4402 3834 4408 3836
rect 4162 3782 4164 3834
rect 4344 3782 4346 3834
rect 4100 3780 4106 3782
rect 4162 3780 4186 3782
rect 4242 3780 4266 3782
rect 4322 3780 4346 3782
rect 4402 3780 4408 3782
rect 4100 3771 4408 3780
rect 2249 3292 2557 3301
rect 2249 3290 2255 3292
rect 2311 3290 2335 3292
rect 2391 3290 2415 3292
rect 2471 3290 2495 3292
rect 2551 3290 2557 3292
rect 2311 3238 2313 3290
rect 2493 3238 2495 3290
rect 2249 3236 2255 3238
rect 2311 3236 2335 3238
rect 2391 3236 2415 3238
rect 2471 3236 2495 3238
rect 2551 3236 2557 3238
rect 2249 3227 2557 3236
rect 4540 3058 4568 3878
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4100 2748 4408 2757
rect 4100 2746 4106 2748
rect 4162 2746 4186 2748
rect 4242 2746 4266 2748
rect 4322 2746 4346 2748
rect 4402 2746 4408 2748
rect 4162 2694 4164 2746
rect 4344 2694 4346 2746
rect 4100 2692 4106 2694
rect 4162 2692 4186 2694
rect 4242 2692 4266 2694
rect 4322 2692 4346 2694
rect 4402 2692 4408 2694
rect 4100 2683 4408 2692
rect 5828 2514 5856 5102
rect 6012 4826 6040 5102
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 5951 4380 6259 4389
rect 5951 4378 5957 4380
rect 6013 4378 6037 4380
rect 6093 4378 6117 4380
rect 6173 4378 6197 4380
rect 6253 4378 6259 4380
rect 6013 4326 6015 4378
rect 6195 4326 6197 4378
rect 5951 4324 5957 4326
rect 6013 4324 6037 4326
rect 6093 4324 6117 4326
rect 6173 4324 6197 4326
rect 6253 4324 6259 4326
rect 5951 4315 6259 4324
rect 6288 4282 6316 4694
rect 6380 4690 6408 5578
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6564 4826 6592 4966
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6656 4690 6684 7142
rect 7024 6934 7052 7958
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7300 7410 7328 7686
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 7024 6254 7052 6870
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6932 5574 6960 6122
rect 7300 6118 7328 7346
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7392 5778 7420 8230
rect 7484 6390 7512 8230
rect 7576 8090 7604 8978
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 7802 8188 8110 8197
rect 7802 8186 7808 8188
rect 7864 8186 7888 8188
rect 7944 8186 7968 8188
rect 8024 8186 8048 8188
rect 8104 8186 8110 8188
rect 7864 8134 7866 8186
rect 8046 8134 8048 8186
rect 7802 8132 7808 8134
rect 7864 8132 7888 8134
rect 7944 8132 7968 8134
rect 8024 8132 8048 8134
rect 8104 8132 8110 8134
rect 7802 8123 8110 8132
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 8312 7410 8340 8366
rect 8404 8090 8432 11018
rect 8772 11014 8800 12106
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8588 10266 8616 10678
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8680 10266 8708 10610
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8680 10130 8708 10202
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8496 9722 8524 10066
rect 8680 9722 8708 10066
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8588 9586 8616 9658
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8588 9042 8616 9522
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8588 8430 8616 8978
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8680 8362 8708 8434
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8680 7290 8708 8298
rect 8864 7954 8892 12174
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8956 11354 8984 11562
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8944 10532 8996 10538
rect 8944 10474 8996 10480
rect 8956 8838 8984 10474
rect 9048 9450 9076 12718
rect 9140 12170 9168 14214
rect 9232 14074 9260 14418
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9324 12986 9352 13330
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9128 12164 9180 12170
rect 9128 12106 9180 12112
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9232 11694 9260 12038
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9324 10606 9352 11834
rect 9416 11694 9444 12038
rect 9508 11762 9536 14350
rect 9653 14172 9961 14181
rect 9653 14170 9659 14172
rect 9715 14170 9739 14172
rect 9795 14170 9819 14172
rect 9875 14170 9899 14172
rect 9955 14170 9961 14172
rect 9715 14118 9717 14170
rect 9897 14118 9899 14170
rect 9653 14116 9659 14118
rect 9715 14116 9739 14118
rect 9795 14116 9819 14118
rect 9875 14116 9899 14118
rect 9955 14116 9961 14118
rect 9653 14107 9961 14116
rect 10152 14074 10180 14350
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10244 13870 10272 14350
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 9653 13084 9961 13093
rect 9653 13082 9659 13084
rect 9715 13082 9739 13084
rect 9795 13082 9819 13084
rect 9875 13082 9899 13084
rect 9955 13082 9961 13084
rect 9715 13030 9717 13082
rect 9897 13030 9899 13082
rect 9653 13028 9659 13030
rect 9715 13028 9739 13030
rect 9795 13028 9819 13030
rect 9875 13028 9899 13030
rect 9955 13028 9961 13030
rect 9653 13019 9961 13028
rect 10244 12850 10272 13806
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10428 12782 10456 13126
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10428 12170 10456 12718
rect 10520 12646 10548 14826
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10796 14006 10824 14758
rect 10888 14074 10916 15098
rect 11164 14958 11192 15600
rect 12452 14958 12480 15600
rect 13355 15260 13663 15269
rect 13355 15258 13361 15260
rect 13417 15258 13441 15260
rect 13497 15258 13521 15260
rect 13577 15258 13601 15260
rect 13657 15258 13663 15260
rect 13417 15206 13419 15258
rect 13599 15206 13601 15258
rect 13355 15204 13361 15206
rect 13417 15204 13441 15206
rect 13497 15204 13521 15206
rect 13577 15204 13601 15206
rect 13657 15204 13663 15206
rect 13355 15195 13663 15204
rect 13740 14958 13768 15600
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 11348 14414 11376 14758
rect 11504 14716 11812 14725
rect 11504 14714 11510 14716
rect 11566 14714 11590 14716
rect 11646 14714 11670 14716
rect 11726 14714 11750 14716
rect 11806 14714 11812 14716
rect 11566 14662 11568 14714
rect 11748 14662 11750 14714
rect 11504 14660 11510 14662
rect 11566 14660 11590 14662
rect 11646 14660 11670 14662
rect 11726 14660 11750 14662
rect 11806 14660 11812 14662
rect 11504 14651 11812 14660
rect 12820 14550 12848 14758
rect 14016 14618 14044 14758
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 12808 14544 12860 14550
rect 12808 14486 12860 14492
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10784 14000 10836 14006
rect 10784 13942 10836 13948
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 9653 11996 9961 12005
rect 9653 11994 9659 11996
rect 9715 11994 9739 11996
rect 9795 11994 9819 11996
rect 9875 11994 9899 11996
rect 9955 11994 9961 11996
rect 9715 11942 9717 11994
rect 9897 11942 9899 11994
rect 9653 11940 9659 11942
rect 9715 11940 9739 11942
rect 9795 11940 9819 11942
rect 9875 11940 9899 11942
rect 9955 11940 9961 11942
rect 9653 11931 9961 11940
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9692 11354 9720 11562
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9416 10418 9444 10950
rect 9324 10390 9444 10418
rect 9324 9994 9352 10390
rect 9508 10282 9536 11018
rect 9653 10908 9961 10917
rect 9653 10906 9659 10908
rect 9715 10906 9739 10908
rect 9795 10906 9819 10908
rect 9875 10906 9899 10908
rect 9955 10906 9961 10908
rect 9715 10854 9717 10906
rect 9897 10854 9899 10906
rect 9653 10852 9659 10854
rect 9715 10852 9739 10854
rect 9795 10852 9819 10854
rect 9875 10852 9899 10854
rect 9955 10852 9961 10854
rect 9653 10843 9961 10852
rect 9416 10254 9536 10282
rect 9416 10130 9444 10254
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9036 9444 9088 9450
rect 9036 9386 9088 9392
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8864 7342 8892 7890
rect 8852 7336 8904 7342
rect 7668 7002 7696 7278
rect 7802 7100 8110 7109
rect 7802 7098 7808 7100
rect 7864 7098 7888 7100
rect 7944 7098 7968 7100
rect 8024 7098 8048 7100
rect 8104 7098 8110 7100
rect 7864 7046 7866 7098
rect 8046 7046 8048 7098
rect 7802 7044 7808 7046
rect 7864 7044 7888 7046
rect 7944 7044 7968 7046
rect 8024 7044 8048 7046
rect 8104 7044 8110 7046
rect 7802 7035 8110 7044
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7668 6866 7696 6938
rect 8220 6934 8248 7278
rect 8680 7274 8800 7290
rect 8852 7278 8904 7284
rect 8300 7268 8352 7274
rect 8680 7268 8812 7274
rect 8680 7262 8760 7268
rect 8300 7210 8352 7216
rect 8760 7210 8812 7216
rect 8312 7002 8340 7210
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8404 7002 8432 7142
rect 8864 7002 8892 7278
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7470 6216 7526 6225
rect 7470 6151 7526 6160
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7392 5658 7420 5714
rect 7208 5630 7420 5658
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6932 5234 6960 5510
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 7208 4486 7236 5630
rect 7484 5534 7512 6151
rect 7392 5506 7512 5534
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7300 4622 7328 4966
rect 7392 4690 7420 5506
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7484 4706 7512 4966
rect 7576 4826 7604 6326
rect 7668 5534 7696 6802
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8588 6254 8616 6598
rect 8576 6248 8628 6254
rect 7746 6216 7802 6225
rect 8576 6190 8628 6196
rect 7746 6151 7802 6160
rect 8208 6180 8260 6186
rect 7760 6118 7788 6151
rect 8208 6122 8260 6128
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7802 6012 8110 6021
rect 7802 6010 7808 6012
rect 7864 6010 7888 6012
rect 7944 6010 7968 6012
rect 8024 6010 8048 6012
rect 8104 6010 8110 6012
rect 7864 5958 7866 6010
rect 8046 5958 8048 6010
rect 7802 5956 7808 5958
rect 7864 5956 7888 5958
rect 7944 5956 7968 5958
rect 8024 5956 8048 5958
rect 8104 5956 8110 5958
rect 7802 5947 8110 5956
rect 8220 5778 8248 6122
rect 8956 5846 8984 8774
rect 9140 8430 9168 9318
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9048 8090 9076 8230
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 9048 6730 9076 7822
rect 9140 7546 9168 8366
rect 9324 7886 9352 9930
rect 9416 9382 9444 10066
rect 10060 9926 10088 11018
rect 10152 10810 10180 11154
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10152 10198 10180 10542
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10244 10198 10272 10406
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10232 10192 10284 10198
rect 10232 10134 10284 10140
rect 10336 10130 10364 10950
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9653 9820 9961 9829
rect 9653 9818 9659 9820
rect 9715 9818 9739 9820
rect 9795 9818 9819 9820
rect 9875 9818 9899 9820
rect 9955 9818 9961 9820
rect 9715 9766 9717 9818
rect 9897 9766 9899 9818
rect 9653 9764 9659 9766
rect 9715 9764 9739 9766
rect 9795 9764 9819 9766
rect 9875 9764 9899 9766
rect 9955 9764 9961 9766
rect 9653 9755 9961 9764
rect 10152 9518 10180 9930
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9416 7818 9444 9318
rect 9653 8732 9961 8741
rect 9653 8730 9659 8732
rect 9715 8730 9739 8732
rect 9795 8730 9819 8732
rect 9875 8730 9899 8732
rect 9955 8730 9961 8732
rect 9715 8678 9717 8730
rect 9897 8678 9899 8730
rect 9653 8676 9659 8678
rect 9715 8676 9739 8678
rect 9795 8676 9819 8678
rect 9875 8676 9899 8678
rect 9955 8676 9961 8678
rect 9653 8667 9961 8676
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9692 8090 9720 8298
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9653 7644 9961 7653
rect 9653 7642 9659 7644
rect 9715 7642 9739 7644
rect 9795 7642 9819 7644
rect 9875 7642 9899 7644
rect 9955 7642 9961 7644
rect 9715 7590 9717 7642
rect 9897 7590 9899 7642
rect 9653 7588 9659 7590
rect 9715 7588 9739 7590
rect 9795 7588 9819 7590
rect 9875 7588 9899 7590
rect 9955 7588 9961 7590
rect 9653 7579 9961 7588
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 10428 7410 10456 7890
rect 10520 7410 10548 12582
rect 10704 8974 10732 12922
rect 10796 9518 10824 13942
rect 10980 13870 11008 14214
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 11072 12986 11100 14010
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11256 12646 11284 13262
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11256 11694 11284 12582
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11164 11218 11192 11494
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10888 9654 10916 10202
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10888 9518 10916 9590
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10888 9382 10916 9454
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10980 9042 11008 9318
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10692 8968 10744 8974
rect 11072 8956 11100 9998
rect 11164 9518 11192 10134
rect 11256 9722 11284 11630
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11152 9512 11204 9518
rect 11256 9489 11284 9658
rect 11152 9454 11204 9460
rect 11242 9480 11298 9489
rect 11242 9415 11298 9424
rect 11152 8968 11204 8974
rect 11072 8928 11152 8956
rect 10692 8910 10744 8916
rect 11152 8910 11204 8916
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10244 6866 10272 7210
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10520 6866 10548 7142
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 9508 6458 9536 6802
rect 9653 6556 9961 6565
rect 9653 6554 9659 6556
rect 9715 6554 9739 6556
rect 9795 6554 9819 6556
rect 9875 6554 9899 6556
rect 9955 6554 9961 6556
rect 9715 6502 9717 6554
rect 9897 6502 9899 6554
rect 9653 6500 9659 6502
rect 9715 6500 9739 6502
rect 9795 6500 9819 6502
rect 9875 6500 9899 6502
rect 9955 6500 9961 6502
rect 9653 6491 9961 6500
rect 10612 6458 10640 6802
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10704 6186 10732 8910
rect 10876 8560 10928 8566
rect 10876 8502 10928 8508
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10796 6866 10824 8366
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 7668 5506 7788 5534
rect 7760 5098 7788 5506
rect 8036 5234 8064 5646
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8220 5302 8248 5510
rect 9653 5468 9961 5477
rect 9653 5466 9659 5468
rect 9715 5466 9739 5468
rect 9795 5466 9819 5468
rect 9875 5466 9899 5468
rect 9955 5466 9961 5468
rect 9715 5414 9717 5466
rect 9897 5414 9899 5466
rect 9653 5412 9659 5414
rect 9715 5412 9739 5414
rect 9795 5412 9819 5414
rect 9875 5412 9899 5414
rect 9955 5412 9961 5414
rect 9653 5403 9961 5412
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7668 4826 7696 4966
rect 7802 4924 8110 4933
rect 7802 4922 7808 4924
rect 7864 4922 7888 4924
rect 7944 4922 7968 4924
rect 8024 4922 8048 4924
rect 8104 4922 8110 4924
rect 7864 4870 7866 4922
rect 8046 4870 8048 4922
rect 7802 4868 7808 4870
rect 7864 4868 7888 4870
rect 7944 4868 7968 4870
rect 8024 4868 8048 4870
rect 8104 4868 8110 4870
rect 7802 4859 8110 4868
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7840 4752 7892 4758
rect 7484 4690 7604 4706
rect 7840 4694 7892 4700
rect 8220 4706 8248 5238
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 8312 4826 8340 5102
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 7380 4684 7432 4690
rect 7484 4684 7616 4690
rect 7484 4678 7564 4684
rect 7380 4626 7432 4632
rect 7564 4626 7616 4632
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7484 4282 7512 4490
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6656 3466 6684 3946
rect 7576 3942 7604 4626
rect 7852 4010 7880 4694
rect 7932 4684 7984 4690
rect 8220 4678 8340 4706
rect 7932 4626 7984 4632
rect 7944 4078 7972 4626
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8128 4146 8156 4558
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7840 4004 7892 4010
rect 7840 3946 7892 3952
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7576 3738 7604 3878
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7668 3482 7696 3946
rect 7802 3836 8110 3845
rect 7802 3834 7808 3836
rect 7864 3834 7888 3836
rect 7944 3834 7968 3836
rect 8024 3834 8048 3836
rect 8104 3834 8110 3836
rect 7864 3782 7866 3834
rect 8046 3782 8048 3834
rect 7802 3780 7808 3782
rect 7864 3780 7888 3782
rect 7944 3780 7968 3782
rect 8024 3780 8048 3782
rect 8104 3780 8110 3782
rect 7802 3771 8110 3780
rect 7932 3664 7984 3670
rect 7932 3606 7984 3612
rect 7748 3528 7800 3534
rect 7668 3476 7748 3482
rect 7668 3470 7800 3476
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 7668 3454 7788 3470
rect 5951 3292 6259 3301
rect 5951 3290 5957 3292
rect 6013 3290 6037 3292
rect 6093 3290 6117 3292
rect 6173 3290 6197 3292
rect 6253 3290 6259 3292
rect 6013 3238 6015 3290
rect 6195 3238 6197 3290
rect 5951 3236 5957 3238
rect 6013 3236 6037 3238
rect 6093 3236 6117 3238
rect 6173 3236 6197 3238
rect 6253 3236 6259 3238
rect 5951 3227 6259 3236
rect 6656 2990 6684 3402
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7576 2990 7604 3334
rect 7668 3194 7696 3454
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7944 3058 7972 3606
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 8220 2990 8248 4014
rect 8312 3398 8340 4678
rect 9968 4570 9996 4966
rect 10060 4690 10088 4966
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10428 4593 10456 5102
rect 10414 4584 10470 4593
rect 9968 4542 10272 4570
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8944 4208 8996 4214
rect 8944 4150 8996 4156
rect 8772 4010 8800 4150
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8772 3194 8800 3470
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8956 2990 8984 4150
rect 9508 4078 9536 4422
rect 9653 4380 9961 4389
rect 9653 4378 9659 4380
rect 9715 4378 9739 4380
rect 9795 4378 9819 4380
rect 9875 4378 9899 4380
rect 9955 4378 9961 4380
rect 9715 4326 9717 4378
rect 9897 4326 9899 4378
rect 9653 4324 9659 4326
rect 9715 4324 9739 4326
rect 9795 4324 9819 4326
rect 9875 4324 9899 4326
rect 9955 4324 9961 4326
rect 9653 4315 9961 4324
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9140 3738 9168 3878
rect 9232 3738 9260 4014
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 9416 3602 9444 3878
rect 10244 3738 10272 4542
rect 10414 4519 10470 4528
rect 10428 4078 10456 4519
rect 10520 4078 10548 6122
rect 10796 5914 10824 6802
rect 10888 6118 10916 8502
rect 11256 8022 11284 9415
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11348 7886 11376 14350
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12084 13870 12112 14010
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12164 13864 12216 13870
rect 12348 13864 12400 13870
rect 12164 13806 12216 13812
rect 12346 13832 12348 13841
rect 12400 13832 12402 13841
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 11440 12782 11468 13738
rect 11504 13628 11812 13637
rect 11504 13626 11510 13628
rect 11566 13626 11590 13628
rect 11646 13626 11670 13628
rect 11726 13626 11750 13628
rect 11806 13626 11812 13628
rect 11566 13574 11568 13626
rect 11748 13574 11750 13626
rect 11504 13572 11510 13574
rect 11566 13572 11590 13574
rect 11646 13572 11670 13574
rect 11726 13572 11750 13574
rect 11806 13572 11812 13574
rect 11504 13563 11812 13572
rect 11900 13530 11928 13806
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11808 12986 11836 13330
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11900 12850 11928 13330
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11504 12540 11812 12549
rect 11504 12538 11510 12540
rect 11566 12538 11590 12540
rect 11646 12538 11670 12540
rect 11726 12538 11750 12540
rect 11806 12538 11812 12540
rect 11566 12486 11568 12538
rect 11748 12486 11750 12538
rect 11504 12484 11510 12486
rect 11566 12484 11590 12486
rect 11646 12484 11670 12486
rect 11726 12484 11750 12486
rect 11806 12484 11812 12486
rect 11504 12475 11812 12484
rect 11992 12442 12020 12582
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11440 11150 11468 12174
rect 11504 11452 11812 11461
rect 11504 11450 11510 11452
rect 11566 11450 11590 11452
rect 11646 11450 11670 11452
rect 11726 11450 11750 11452
rect 11806 11450 11812 11452
rect 11566 11398 11568 11450
rect 11748 11398 11750 11450
rect 11504 11396 11510 11398
rect 11566 11396 11590 11398
rect 11646 11396 11670 11398
rect 11726 11396 11750 11398
rect 11806 11396 11812 11398
rect 11504 11387 11812 11396
rect 11900 11354 11928 12378
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 12084 11218 12112 13398
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11440 8566 11468 11086
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 11504 10364 11812 10373
rect 11504 10362 11510 10364
rect 11566 10362 11590 10364
rect 11646 10362 11670 10364
rect 11726 10362 11750 10364
rect 11806 10362 11812 10364
rect 11566 10310 11568 10362
rect 11748 10310 11750 10362
rect 11504 10308 11510 10310
rect 11566 10308 11590 10310
rect 11646 10308 11670 10310
rect 11726 10308 11750 10310
rect 11806 10308 11812 10310
rect 11504 10299 11812 10308
rect 12084 9586 12112 10474
rect 12176 10198 12204 13806
rect 12346 13767 12402 13776
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12268 13530 12296 13670
rect 12452 13530 12480 14418
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 13355 14172 13663 14181
rect 13355 14170 13361 14172
rect 13417 14170 13441 14172
rect 13497 14170 13521 14172
rect 13577 14170 13601 14172
rect 13657 14170 13663 14172
rect 13417 14118 13419 14170
rect 13599 14118 13601 14170
rect 13355 14116 13361 14118
rect 13417 14116 13441 14118
rect 13497 14116 13521 14118
rect 13577 14116 13601 14118
rect 13657 14116 13663 14118
rect 13355 14107 13663 14116
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 12900 14000 12952 14006
rect 12900 13942 12952 13948
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12636 13530 12664 13806
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12820 13394 12848 13670
rect 12912 13394 12940 13942
rect 12992 13796 13044 13802
rect 12992 13738 13044 13744
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12360 12850 12388 13330
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12256 12708 12308 12714
rect 12256 12650 12308 12656
rect 12268 12238 12296 12650
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12360 11218 12388 12786
rect 12544 12442 12572 13126
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12900 12912 12952 12918
rect 12900 12854 12952 12860
rect 12636 12714 12664 12854
rect 12912 12714 12940 12854
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12636 11898 12664 12650
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12912 11642 12940 11834
rect 12820 11614 12940 11642
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12452 11218 12480 11494
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12360 10674 12388 11154
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12164 10192 12216 10198
rect 12164 10134 12216 10140
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 11504 9276 11812 9285
rect 11504 9274 11510 9276
rect 11566 9274 11590 9276
rect 11646 9274 11670 9276
rect 11726 9274 11750 9276
rect 11806 9274 11812 9276
rect 11566 9222 11568 9274
rect 11748 9222 11750 9274
rect 11504 9220 11510 9222
rect 11566 9220 11590 9222
rect 11646 9220 11670 9222
rect 11726 9220 11750 9222
rect 11806 9220 11812 9222
rect 11504 9211 11812 9220
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11532 9058 11560 9114
rect 11716 9058 11744 9114
rect 12176 9110 12204 10134
rect 12360 10010 12388 10610
rect 12452 10130 12480 10950
rect 12636 10810 12664 11154
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12360 9982 12480 10010
rect 12452 9926 12480 9982
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12452 9518 12480 9862
rect 12624 9648 12676 9654
rect 12728 9602 12756 11154
rect 12820 10742 12848 11614
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12820 10146 12848 10678
rect 12912 10606 12940 11494
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12912 10169 12940 10406
rect 12898 10160 12954 10169
rect 12820 10130 12898 10146
rect 12808 10124 12898 10130
rect 12860 10118 12898 10124
rect 12898 10095 12954 10104
rect 12808 10066 12860 10072
rect 12806 10024 12862 10033
rect 12806 9959 12808 9968
rect 12860 9959 12862 9968
rect 12808 9930 12860 9936
rect 12676 9596 12756 9602
rect 12624 9590 12756 9596
rect 12636 9574 12756 9590
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12624 9512 12676 9518
rect 12728 9500 12756 9574
rect 12808 9512 12860 9518
rect 12728 9472 12808 9500
rect 12624 9454 12676 9460
rect 12808 9454 12860 9460
rect 11532 9030 11744 9058
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11520 8968 11572 8974
rect 11704 8968 11756 8974
rect 11572 8928 11704 8956
rect 11520 8910 11572 8916
rect 11704 8910 11756 8916
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11716 8430 11744 8774
rect 11808 8634 11836 8774
rect 11992 8634 12020 8978
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11440 7954 11468 8230
rect 11504 8188 11812 8197
rect 11504 8186 11510 8188
rect 11566 8186 11590 8188
rect 11646 8186 11670 8188
rect 11726 8186 11750 8188
rect 11806 8186 11812 8188
rect 11566 8134 11568 8186
rect 11748 8134 11750 8186
rect 11504 8132 11510 8134
rect 11566 8132 11590 8134
rect 11646 8132 11670 8134
rect 11726 8132 11750 8134
rect 11806 8132 11812 8134
rect 11504 8123 11812 8132
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 12256 7948 12308 7954
rect 12256 7890 12308 7896
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 11504 7100 11812 7109
rect 11504 7098 11510 7100
rect 11566 7098 11590 7100
rect 11646 7098 11670 7100
rect 11726 7098 11750 7100
rect 11806 7098 11812 7100
rect 11566 7046 11568 7098
rect 11748 7046 11750 7098
rect 11504 7044 11510 7046
rect 11566 7044 11590 7046
rect 11646 7044 11670 7046
rect 11726 7044 11750 7046
rect 11806 7044 11812 7046
rect 11504 7035 11812 7044
rect 12084 7002 12112 7278
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 11716 6186 11744 6938
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11704 6180 11756 6186
rect 11704 6122 11756 6128
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10888 5574 10916 6054
rect 10876 5568 10928 5574
rect 10704 5516 10876 5534
rect 10704 5510 10928 5516
rect 10704 5506 10916 5510
rect 10704 5386 10732 5506
rect 10612 5358 10732 5386
rect 11348 5370 11376 6122
rect 11900 6118 11928 6258
rect 12176 6254 12204 7686
rect 12268 7342 12296 7890
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12452 6934 12480 9454
rect 12636 9110 12664 9454
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12544 8498 12572 8978
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12820 8294 12848 8570
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12636 7410 12664 8230
rect 12820 7954 12848 8230
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12636 6866 12664 7210
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12820 6730 12848 7890
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 12532 6656 12584 6662
rect 13004 6610 13032 13738
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 13280 12306 13308 13398
rect 13355 13084 13663 13093
rect 13355 13082 13361 13084
rect 13417 13082 13441 13084
rect 13497 13082 13521 13084
rect 13577 13082 13601 13084
rect 13657 13082 13663 13084
rect 13417 13030 13419 13082
rect 13599 13030 13601 13082
rect 13355 13028 13361 13030
rect 13417 13028 13441 13030
rect 13497 13028 13521 13030
rect 13577 13028 13601 13030
rect 13657 13028 13663 13030
rect 13355 13019 13663 13028
rect 13924 12782 13952 14010
rect 14200 13938 14228 14214
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14464 13864 14516 13870
rect 14462 13832 14464 13841
rect 14516 13832 14518 13841
rect 14462 13767 14518 13776
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14660 12782 14688 13670
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13648 12306 13676 12582
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 13096 11082 13124 11562
rect 13280 11218 13308 12242
rect 13355 11996 13663 12005
rect 13355 11994 13361 11996
rect 13417 11994 13441 11996
rect 13497 11994 13521 11996
rect 13577 11994 13601 11996
rect 13657 11994 13663 11996
rect 13417 11942 13419 11994
rect 13599 11942 13601 11994
rect 13355 11940 13361 11942
rect 13417 11940 13441 11942
rect 13497 11940 13521 11942
rect 13577 11940 13601 11942
rect 13657 11940 13663 11942
rect 13355 11931 13663 11940
rect 13924 11694 13952 12718
rect 14200 11694 14228 12718
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 11218 13676 11494
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 13096 10810 13124 11018
rect 13188 10810 13216 11086
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13084 10600 13136 10606
rect 13084 10542 13136 10548
rect 13096 10470 13124 10542
rect 13280 10538 13308 11154
rect 13355 10908 13663 10917
rect 13355 10906 13361 10908
rect 13417 10906 13441 10908
rect 13497 10906 13521 10908
rect 13577 10906 13601 10908
rect 13657 10906 13663 10908
rect 13417 10854 13419 10906
rect 13599 10854 13601 10906
rect 13355 10852 13361 10854
rect 13417 10852 13441 10854
rect 13497 10852 13521 10854
rect 13577 10852 13601 10854
rect 13657 10852 13663 10854
rect 13355 10843 13663 10852
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13096 9364 13124 10406
rect 13280 10010 13308 10474
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13360 10056 13412 10062
rect 13280 10004 13360 10010
rect 13464 10033 13492 10066
rect 13280 9998 13412 10004
rect 13450 10024 13506 10033
rect 13176 9988 13228 9994
rect 13176 9930 13228 9936
rect 13280 9982 13400 9998
rect 13188 9722 13216 9930
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13176 9512 13228 9518
rect 13174 9480 13176 9489
rect 13228 9480 13230 9489
rect 13174 9415 13230 9424
rect 13176 9376 13228 9382
rect 13096 9336 13176 9364
rect 13176 9318 13228 9324
rect 13188 8634 13216 9318
rect 13280 9110 13308 9982
rect 13450 9959 13506 9968
rect 13355 9820 13663 9829
rect 13355 9818 13361 9820
rect 13417 9818 13441 9820
rect 13497 9818 13521 9820
rect 13577 9818 13601 9820
rect 13657 9818 13663 9820
rect 13417 9766 13419 9818
rect 13599 9766 13601 9818
rect 13355 9764 13361 9766
rect 13417 9764 13441 9766
rect 13497 9764 13521 9766
rect 13577 9764 13601 9766
rect 13657 9764 13663 9766
rect 13355 9755 13663 9764
rect 13924 9518 13952 11630
rect 14016 11354 14044 11630
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 14200 11054 14228 11630
rect 14108 11026 14228 11054
rect 14108 10266 14136 11026
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14108 9518 14136 10202
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13648 9042 13676 9318
rect 13924 9042 13952 9454
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13355 8732 13663 8741
rect 13355 8730 13361 8732
rect 13417 8730 13441 8732
rect 13497 8730 13521 8732
rect 13577 8730 13601 8732
rect 13657 8730 13663 8732
rect 13417 8678 13419 8730
rect 13599 8678 13601 8730
rect 13355 8676 13361 8678
rect 13417 8676 13441 8678
rect 13497 8676 13521 8678
rect 13577 8676 13601 8678
rect 13657 8676 13663 8678
rect 13355 8667 13663 8676
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13924 8430 13952 8978
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13084 7472 13136 7478
rect 13084 7414 13136 7420
rect 13096 6866 13124 7414
rect 13188 7342 13216 8230
rect 13648 7954 13676 8230
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 13280 6934 13308 7822
rect 13355 7644 13663 7653
rect 13355 7642 13361 7644
rect 13417 7642 13441 7644
rect 13497 7642 13521 7644
rect 13577 7642 13601 7644
rect 13657 7642 13663 7644
rect 13417 7590 13419 7642
rect 13599 7590 13601 7642
rect 13355 7588 13361 7590
rect 13417 7588 13441 7590
rect 13497 7588 13521 7590
rect 13577 7588 13601 7590
rect 13657 7588 13663 7590
rect 13355 7579 13663 7588
rect 13924 7002 13952 8366
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 12532 6598 12584 6604
rect 12544 6254 12572 6598
rect 12912 6582 13032 6610
rect 12912 6254 12940 6582
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11504 6012 11812 6021
rect 11504 6010 11510 6012
rect 11566 6010 11590 6012
rect 11646 6010 11670 6012
rect 11726 6010 11750 6012
rect 11806 6010 11812 6012
rect 11566 5958 11568 6010
rect 11748 5958 11750 6010
rect 11504 5956 11510 5958
rect 11566 5956 11590 5958
rect 11646 5956 11670 5958
rect 11726 5956 11750 5958
rect 11806 5956 11812 5958
rect 11504 5947 11812 5956
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11336 5364 11388 5370
rect 10612 5234 10640 5358
rect 11336 5306 11388 5312
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10874 5128 10930 5137
rect 10704 4554 10732 5102
rect 10796 4554 10824 5102
rect 10874 5063 10930 5072
rect 11244 5092 11296 5098
rect 10888 4826 10916 5063
rect 11244 5034 11296 5040
rect 11256 4826 11284 5034
rect 11348 4826 11376 5306
rect 11888 5160 11940 5166
rect 11886 5128 11888 5137
rect 11940 5128 11942 5137
rect 11886 5063 11942 5072
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 11256 4486 11284 4762
rect 11348 4690 11376 4762
rect 11440 4690 11468 4966
rect 11504 4924 11812 4933
rect 11504 4922 11510 4924
rect 11566 4922 11590 4924
rect 11646 4922 11670 4924
rect 11726 4922 11750 4924
rect 11806 4922 11812 4924
rect 11566 4870 11568 4922
rect 11748 4870 11750 4922
rect 11504 4868 11510 4870
rect 11566 4868 11590 4870
rect 11646 4868 11670 4870
rect 11726 4868 11750 4870
rect 11806 4868 11812 4870
rect 11504 4859 11812 4868
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11256 4078 11284 4422
rect 11348 4282 11376 4626
rect 11518 4584 11574 4593
rect 11518 4519 11520 4528
rect 11572 4519 11574 4528
rect 11520 4490 11572 4496
rect 11808 4282 11836 4694
rect 11900 4282 11928 4966
rect 11992 4690 12020 5850
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 12084 5234 12112 5510
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 12452 5166 12480 5306
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12360 4826 12388 5102
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9140 3482 9168 3538
rect 9048 3466 9168 3482
rect 9036 3460 9168 3466
rect 9088 3454 9168 3460
rect 9036 3402 9088 3408
rect 9653 3292 9961 3301
rect 9653 3290 9659 3292
rect 9715 3290 9739 3292
rect 9795 3290 9819 3292
rect 9875 3290 9899 3292
rect 9955 3290 9961 3292
rect 9715 3238 9717 3290
rect 9897 3238 9899 3290
rect 9653 3236 9659 3238
rect 9715 3236 9739 3238
rect 9795 3236 9819 3238
rect 9875 3236 9899 3238
rect 9955 3236 9961 3238
rect 9653 3227 9961 3236
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 5908 2916 5960 2922
rect 5908 2858 5960 2864
rect 5920 2650 5948 2858
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 6932 2514 6960 2790
rect 7802 2748 8110 2757
rect 7802 2746 7808 2748
rect 7864 2746 7888 2748
rect 7944 2746 7968 2748
rect 8024 2746 8048 2748
rect 8104 2746 8110 2748
rect 7864 2694 7866 2746
rect 8046 2694 8048 2746
rect 7802 2692 7808 2694
rect 7864 2692 7888 2694
rect 7944 2692 7968 2694
rect 8024 2692 8048 2694
rect 8104 2692 8110 2694
rect 7802 2683 8110 2692
rect 10244 2514 10272 3674
rect 10520 3670 10548 4014
rect 11256 3738 11284 4014
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 10336 2650 10364 2858
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10980 2514 11008 3334
rect 11256 3194 11284 3674
rect 11348 3602 11376 3878
rect 11504 3836 11812 3845
rect 11504 3834 11510 3836
rect 11566 3834 11590 3836
rect 11646 3834 11670 3836
rect 11726 3834 11750 3836
rect 11806 3834 11812 3836
rect 11566 3782 11568 3834
rect 11748 3782 11750 3834
rect 11504 3780 11510 3782
rect 11566 3780 11590 3782
rect 11646 3780 11670 3782
rect 11726 3780 11750 3782
rect 11806 3780 11812 3782
rect 11504 3771 11812 3780
rect 11900 3738 11928 4014
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11992 3058 12020 4626
rect 12912 4078 12940 6190
rect 13004 5710 13032 6326
rect 13096 6254 13124 6802
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13188 6254 13216 6598
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13280 5710 13308 6870
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13355 6556 13663 6565
rect 13355 6554 13361 6556
rect 13417 6554 13441 6556
rect 13497 6554 13521 6556
rect 13577 6554 13601 6556
rect 13657 6554 13663 6556
rect 13417 6502 13419 6554
rect 13599 6502 13601 6554
rect 13355 6500 13361 6502
rect 13417 6500 13441 6502
rect 13497 6500 13521 6502
rect 13577 6500 13601 6502
rect 13657 6500 13663 6502
rect 13355 6491 13663 6500
rect 13740 6458 13768 6734
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13924 6254 13952 6938
rect 14108 6866 14136 9454
rect 14936 9058 14964 9454
rect 15028 9178 15056 15600
rect 15206 14716 15514 14725
rect 15206 14714 15212 14716
rect 15268 14714 15292 14716
rect 15348 14714 15372 14716
rect 15428 14714 15452 14716
rect 15508 14714 15514 14716
rect 15268 14662 15270 14714
rect 15450 14662 15452 14714
rect 15206 14660 15212 14662
rect 15268 14660 15292 14662
rect 15348 14660 15372 14662
rect 15428 14660 15452 14662
rect 15508 14660 15514 14662
rect 15206 14651 15514 14660
rect 15106 14512 15162 14521
rect 15106 14447 15162 14456
rect 15120 13870 15148 14447
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15120 13530 15148 13806
rect 15206 13628 15514 13637
rect 15206 13626 15212 13628
rect 15268 13626 15292 13628
rect 15348 13626 15372 13628
rect 15428 13626 15452 13628
rect 15508 13626 15514 13628
rect 15268 13574 15270 13626
rect 15450 13574 15452 13626
rect 15206 13572 15212 13574
rect 15268 13572 15292 13574
rect 15348 13572 15372 13574
rect 15428 13572 15452 13574
rect 15508 13572 15514 13574
rect 15206 13563 15514 13572
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15120 12374 15148 12718
rect 15206 12540 15514 12549
rect 15206 12538 15212 12540
rect 15268 12538 15292 12540
rect 15348 12538 15372 12540
rect 15428 12538 15452 12540
rect 15508 12538 15514 12540
rect 15268 12486 15270 12538
rect 15450 12486 15452 12538
rect 15206 12484 15212 12486
rect 15268 12484 15292 12486
rect 15348 12484 15372 12486
rect 15428 12484 15452 12486
rect 15508 12484 15514 12486
rect 15206 12475 15514 12484
rect 15108 12368 15160 12374
rect 15106 12336 15108 12345
rect 15160 12336 15162 12345
rect 15106 12271 15162 12280
rect 15206 11452 15514 11461
rect 15206 11450 15212 11452
rect 15268 11450 15292 11452
rect 15348 11450 15372 11452
rect 15428 11450 15452 11452
rect 15508 11450 15514 11452
rect 15268 11398 15270 11450
rect 15450 11398 15452 11450
rect 15206 11396 15212 11398
rect 15268 11396 15292 11398
rect 15348 11396 15372 11398
rect 15428 11396 15452 11398
rect 15508 11396 15514 11398
rect 15206 11387 15514 11396
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15120 11014 15148 11086
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15120 10713 15148 10950
rect 15106 10704 15162 10713
rect 15106 10639 15162 10648
rect 15206 10364 15514 10373
rect 15206 10362 15212 10364
rect 15268 10362 15292 10364
rect 15348 10362 15372 10364
rect 15428 10362 15452 10364
rect 15508 10362 15514 10364
rect 15268 10310 15270 10362
rect 15450 10310 15452 10362
rect 15206 10308 15212 10310
rect 15268 10308 15292 10310
rect 15348 10308 15372 10310
rect 15428 10308 15452 10310
rect 15508 10308 15514 10310
rect 15206 10299 15514 10308
rect 15106 10160 15162 10169
rect 15106 10095 15162 10104
rect 15120 9926 15148 10095
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 14936 9030 15056 9058
rect 15028 8838 15056 9030
rect 15016 8832 15068 8838
rect 15120 8809 15148 9862
rect 15206 9276 15514 9285
rect 15206 9274 15212 9276
rect 15268 9274 15292 9276
rect 15348 9274 15372 9276
rect 15428 9274 15452 9276
rect 15508 9274 15514 9276
rect 15268 9222 15270 9274
rect 15450 9222 15452 9274
rect 15206 9220 15212 9222
rect 15268 9220 15292 9222
rect 15348 9220 15372 9222
rect 15428 9220 15452 9222
rect 15508 9220 15514 9222
rect 15206 9211 15514 9220
rect 15016 8774 15068 8780
rect 15106 8800 15162 8809
rect 15028 8498 15056 8774
rect 15106 8735 15162 8744
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14936 6746 14964 7278
rect 15028 6905 15056 8434
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15120 7750 15148 8366
rect 15206 8188 15514 8197
rect 15206 8186 15212 8188
rect 15268 8186 15292 8188
rect 15348 8186 15372 8188
rect 15428 8186 15452 8188
rect 15508 8186 15514 8188
rect 15268 8134 15270 8186
rect 15450 8134 15452 8186
rect 15206 8132 15212 8134
rect 15268 8132 15292 8134
rect 15348 8132 15372 8134
rect 15428 8132 15452 8134
rect 15508 8132 15514 8134
rect 15206 8123 15514 8132
rect 15108 7744 15160 7750
rect 15108 7686 15160 7692
rect 15014 6896 15070 6905
rect 15014 6831 15070 6840
rect 14464 6724 14516 6730
rect 14936 6718 15056 6746
rect 14464 6666 14516 6672
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 14476 5574 14504 6666
rect 15028 6662 15056 6718
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 13355 5468 13663 5477
rect 13355 5466 13361 5468
rect 13417 5466 13441 5468
rect 13497 5466 13521 5468
rect 13577 5466 13601 5468
rect 13657 5466 13663 5468
rect 13417 5414 13419 5466
rect 13599 5414 13601 5466
rect 13355 5412 13361 5414
rect 13417 5412 13441 5414
rect 13497 5412 13521 5414
rect 13577 5412 13601 5414
rect 13657 5412 13663 5414
rect 13355 5403 13663 5412
rect 13360 5092 13412 5098
rect 13360 5034 13412 5040
rect 13372 4826 13400 5034
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13355 4380 13663 4389
rect 13355 4378 13361 4380
rect 13417 4378 13441 4380
rect 13497 4378 13521 4380
rect 13577 4378 13601 4380
rect 13657 4378 13663 4380
rect 13417 4326 13419 4378
rect 13599 4326 13601 4378
rect 13355 4324 13361 4326
rect 13417 4324 13441 4326
rect 13497 4324 13521 4326
rect 13577 4324 13601 4326
rect 13657 4324 13663 4326
rect 13355 4315 13663 4324
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 13355 3292 13663 3301
rect 13355 3290 13361 3292
rect 13417 3290 13441 3292
rect 13497 3290 13521 3292
rect 13577 3290 13601 3292
rect 13657 3290 13663 3292
rect 13417 3238 13419 3290
rect 13599 3238 13601 3290
rect 13355 3236 13361 3238
rect 13417 3236 13441 3238
rect 13497 3236 13521 3238
rect 13577 3236 13601 3238
rect 13657 3236 13663 3238
rect 13355 3227 13663 3236
rect 14476 3097 14504 5510
rect 14462 3088 14518 3097
rect 11980 3052 12032 3058
rect 14462 3023 14518 3032
rect 11980 2994 12032 3000
rect 11504 2748 11812 2757
rect 11504 2746 11510 2748
rect 11566 2746 11590 2748
rect 11646 2746 11670 2748
rect 11726 2746 11750 2748
rect 11806 2746 11812 2748
rect 11566 2694 11568 2746
rect 11748 2694 11750 2746
rect 11504 2692 11510 2694
rect 11566 2692 11590 2694
rect 11646 2692 11670 2694
rect 11726 2692 11750 2694
rect 11806 2692 11812 2694
rect 11504 2683 11812 2692
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 2249 2204 2557 2213
rect 2249 2202 2255 2204
rect 2311 2202 2335 2204
rect 2391 2202 2415 2204
rect 2471 2202 2495 2204
rect 2551 2202 2557 2204
rect 2311 2150 2313 2202
rect 2493 2150 2495 2202
rect 2249 2148 2255 2150
rect 2311 2148 2335 2150
rect 2391 2148 2415 2150
rect 2471 2148 2495 2150
rect 2551 2148 2557 2150
rect 2249 2139 2557 2148
rect 5951 2204 6259 2213
rect 5951 2202 5957 2204
rect 6013 2202 6037 2204
rect 6093 2202 6117 2204
rect 6173 2202 6197 2204
rect 6253 2202 6259 2204
rect 6013 2150 6015 2202
rect 6195 2150 6197 2202
rect 5951 2148 5957 2150
rect 6013 2148 6037 2150
rect 6093 2148 6117 2150
rect 6173 2148 6197 2150
rect 6253 2148 6259 2150
rect 5951 2139 6259 2148
rect 9653 2204 9961 2213
rect 9653 2202 9659 2204
rect 9715 2202 9739 2204
rect 9795 2202 9819 2204
rect 9875 2202 9899 2204
rect 9955 2202 9961 2204
rect 9715 2150 9717 2202
rect 9897 2150 9899 2202
rect 9653 2148 9659 2150
rect 9715 2148 9739 2150
rect 9795 2148 9819 2150
rect 9875 2148 9899 2150
rect 9955 2148 9961 2150
rect 9653 2139 9961 2148
rect 13355 2204 13663 2213
rect 13355 2202 13361 2204
rect 13417 2202 13441 2204
rect 13497 2202 13521 2204
rect 13577 2202 13601 2204
rect 13657 2202 13663 2204
rect 13417 2150 13419 2202
rect 13599 2150 13601 2202
rect 13355 2148 13361 2150
rect 13417 2148 13441 2150
rect 13497 2148 13521 2150
rect 13577 2148 13601 2150
rect 13657 2148 13663 2150
rect 13355 2139 13663 2148
rect 4100 1660 4408 1669
rect 4100 1658 4106 1660
rect 4162 1658 4186 1660
rect 4242 1658 4266 1660
rect 4322 1658 4346 1660
rect 4402 1658 4408 1660
rect 4162 1606 4164 1658
rect 4344 1606 4346 1658
rect 4100 1604 4106 1606
rect 4162 1604 4186 1606
rect 4242 1604 4266 1606
rect 4322 1604 4346 1606
rect 4402 1604 4408 1606
rect 4100 1595 4408 1604
rect 7802 1660 8110 1669
rect 7802 1658 7808 1660
rect 7864 1658 7888 1660
rect 7944 1658 7968 1660
rect 8024 1658 8048 1660
rect 8104 1658 8110 1660
rect 7864 1606 7866 1658
rect 8046 1606 8048 1658
rect 7802 1604 7808 1606
rect 7864 1604 7888 1606
rect 7944 1604 7968 1606
rect 8024 1604 8048 1606
rect 8104 1604 8110 1606
rect 7802 1595 8110 1604
rect 11504 1660 11812 1669
rect 11504 1658 11510 1660
rect 11566 1658 11590 1660
rect 11646 1658 11670 1660
rect 11726 1658 11750 1660
rect 11806 1658 11812 1660
rect 11566 1606 11568 1658
rect 11748 1606 11750 1658
rect 11504 1604 11510 1606
rect 11566 1604 11590 1606
rect 11646 1604 11670 1606
rect 11726 1604 11750 1606
rect 11806 1604 11812 1606
rect 11504 1595 11812 1604
rect 15028 1193 15056 6598
rect 15120 5545 15148 7686
rect 15206 7100 15514 7109
rect 15206 7098 15212 7100
rect 15268 7098 15292 7100
rect 15348 7098 15372 7100
rect 15428 7098 15452 7100
rect 15508 7098 15514 7100
rect 15268 7046 15270 7098
rect 15450 7046 15452 7098
rect 15206 7044 15212 7046
rect 15268 7044 15292 7046
rect 15348 7044 15372 7046
rect 15428 7044 15452 7046
rect 15508 7044 15514 7046
rect 15206 7035 15514 7044
rect 15206 6012 15514 6021
rect 15206 6010 15212 6012
rect 15268 6010 15292 6012
rect 15348 6010 15372 6012
rect 15428 6010 15452 6012
rect 15508 6010 15514 6012
rect 15268 5958 15270 6010
rect 15450 5958 15452 6010
rect 15206 5956 15212 5958
rect 15268 5956 15292 5958
rect 15348 5956 15372 5958
rect 15428 5956 15452 5958
rect 15508 5956 15514 5958
rect 15206 5947 15514 5956
rect 15106 5536 15162 5545
rect 15106 5471 15162 5480
rect 15206 4924 15514 4933
rect 15206 4922 15212 4924
rect 15268 4922 15292 4924
rect 15348 4922 15372 4924
rect 15428 4922 15452 4924
rect 15508 4922 15514 4924
rect 15268 4870 15270 4922
rect 15450 4870 15452 4922
rect 15206 4868 15212 4870
rect 15268 4868 15292 4870
rect 15348 4868 15372 4870
rect 15428 4868 15452 4870
rect 15508 4868 15514 4870
rect 15206 4859 15514 4868
rect 15206 3836 15514 3845
rect 15206 3834 15212 3836
rect 15268 3834 15292 3836
rect 15348 3834 15372 3836
rect 15428 3834 15452 3836
rect 15508 3834 15514 3836
rect 15268 3782 15270 3834
rect 15450 3782 15452 3834
rect 15206 3780 15212 3782
rect 15268 3780 15292 3782
rect 15348 3780 15372 3782
rect 15428 3780 15452 3782
rect 15508 3780 15514 3782
rect 15206 3771 15514 3780
rect 15206 2748 15514 2757
rect 15206 2746 15212 2748
rect 15268 2746 15292 2748
rect 15348 2746 15372 2748
rect 15428 2746 15452 2748
rect 15508 2746 15514 2748
rect 15268 2694 15270 2746
rect 15450 2694 15452 2746
rect 15206 2692 15212 2694
rect 15268 2692 15292 2694
rect 15348 2692 15372 2694
rect 15428 2692 15452 2694
rect 15508 2692 15514 2694
rect 15206 2683 15514 2692
rect 15206 1660 15514 1669
rect 15206 1658 15212 1660
rect 15268 1658 15292 1660
rect 15348 1658 15372 1660
rect 15428 1658 15452 1660
rect 15508 1658 15514 1660
rect 15268 1606 15270 1658
rect 15450 1606 15452 1658
rect 15206 1604 15212 1606
rect 15268 1604 15292 1606
rect 15348 1604 15372 1606
rect 15428 1604 15452 1606
rect 15508 1604 15514 1606
rect 15206 1595 15514 1604
rect 15014 1184 15070 1193
rect 2249 1116 2557 1125
rect 2249 1114 2255 1116
rect 2311 1114 2335 1116
rect 2391 1114 2415 1116
rect 2471 1114 2495 1116
rect 2551 1114 2557 1116
rect 2311 1062 2313 1114
rect 2493 1062 2495 1114
rect 2249 1060 2255 1062
rect 2311 1060 2335 1062
rect 2391 1060 2415 1062
rect 2471 1060 2495 1062
rect 2551 1060 2557 1062
rect 2249 1051 2557 1060
rect 5951 1116 6259 1125
rect 5951 1114 5957 1116
rect 6013 1114 6037 1116
rect 6093 1114 6117 1116
rect 6173 1114 6197 1116
rect 6253 1114 6259 1116
rect 6013 1062 6015 1114
rect 6195 1062 6197 1114
rect 5951 1060 5957 1062
rect 6013 1060 6037 1062
rect 6093 1060 6117 1062
rect 6173 1060 6197 1062
rect 6253 1060 6259 1062
rect 5951 1051 6259 1060
rect 9653 1116 9961 1125
rect 9653 1114 9659 1116
rect 9715 1114 9739 1116
rect 9795 1114 9819 1116
rect 9875 1114 9899 1116
rect 9955 1114 9961 1116
rect 9715 1062 9717 1114
rect 9897 1062 9899 1114
rect 9653 1060 9659 1062
rect 9715 1060 9739 1062
rect 9795 1060 9819 1062
rect 9875 1060 9899 1062
rect 9955 1060 9961 1062
rect 9653 1051 9961 1060
rect 13355 1116 13663 1125
rect 15014 1119 15070 1128
rect 13355 1114 13361 1116
rect 13417 1114 13441 1116
rect 13497 1114 13521 1116
rect 13577 1114 13601 1116
rect 13657 1114 13663 1116
rect 13417 1062 13419 1114
rect 13599 1062 13601 1114
rect 13355 1060 13361 1062
rect 13417 1060 13441 1062
rect 13497 1060 13521 1062
rect 13577 1060 13601 1062
rect 13657 1060 13663 1062
rect 13355 1051 13663 1060
rect 4100 572 4408 581
rect 4100 570 4106 572
rect 4162 570 4186 572
rect 4242 570 4266 572
rect 4322 570 4346 572
rect 4402 570 4408 572
rect 4162 518 4164 570
rect 4344 518 4346 570
rect 4100 516 4106 518
rect 4162 516 4186 518
rect 4242 516 4266 518
rect 4322 516 4346 518
rect 4402 516 4408 518
rect 4100 507 4408 516
rect 7802 572 8110 581
rect 7802 570 7808 572
rect 7864 570 7888 572
rect 7944 570 7968 572
rect 8024 570 8048 572
rect 8104 570 8110 572
rect 7864 518 7866 570
rect 8046 518 8048 570
rect 7802 516 7808 518
rect 7864 516 7888 518
rect 7944 516 7968 518
rect 8024 516 8048 518
rect 8104 516 8110 518
rect 7802 507 8110 516
rect 11504 572 11812 581
rect 11504 570 11510 572
rect 11566 570 11590 572
rect 11646 570 11670 572
rect 11726 570 11750 572
rect 11806 570 11812 572
rect 11566 518 11568 570
rect 11748 518 11750 570
rect 11504 516 11510 518
rect 11566 516 11590 518
rect 11646 516 11670 518
rect 11726 516 11750 518
rect 11806 516 11812 518
rect 11504 507 11812 516
rect 15206 572 15514 581
rect 15206 570 15212 572
rect 15268 570 15292 572
rect 15348 570 15372 572
rect 15428 570 15452 572
rect 15508 570 15514 572
rect 15268 518 15270 570
rect 15450 518 15452 570
rect 15206 516 15212 518
rect 15268 516 15292 518
rect 15348 516 15372 518
rect 15428 516 15452 518
rect 15508 516 15514 518
rect 15206 507 15514 516
<< via2 >>
rect 2255 15258 2311 15260
rect 2335 15258 2391 15260
rect 2415 15258 2471 15260
rect 2495 15258 2551 15260
rect 2255 15206 2301 15258
rect 2301 15206 2311 15258
rect 2335 15206 2365 15258
rect 2365 15206 2377 15258
rect 2377 15206 2391 15258
rect 2415 15206 2429 15258
rect 2429 15206 2441 15258
rect 2441 15206 2471 15258
rect 2495 15206 2505 15258
rect 2505 15206 2551 15258
rect 2255 15204 2311 15206
rect 2335 15204 2391 15206
rect 2415 15204 2471 15206
rect 2495 15204 2551 15206
rect 4106 14714 4162 14716
rect 4186 14714 4242 14716
rect 4266 14714 4322 14716
rect 4346 14714 4402 14716
rect 4106 14662 4152 14714
rect 4152 14662 4162 14714
rect 4186 14662 4216 14714
rect 4216 14662 4228 14714
rect 4228 14662 4242 14714
rect 4266 14662 4280 14714
rect 4280 14662 4292 14714
rect 4292 14662 4322 14714
rect 4346 14662 4356 14714
rect 4356 14662 4402 14714
rect 4106 14660 4162 14662
rect 4186 14660 4242 14662
rect 4266 14660 4322 14662
rect 4346 14660 4402 14662
rect 2255 14170 2311 14172
rect 2335 14170 2391 14172
rect 2415 14170 2471 14172
rect 2495 14170 2551 14172
rect 2255 14118 2301 14170
rect 2301 14118 2311 14170
rect 2335 14118 2365 14170
rect 2365 14118 2377 14170
rect 2377 14118 2391 14170
rect 2415 14118 2429 14170
rect 2429 14118 2441 14170
rect 2441 14118 2471 14170
rect 2495 14118 2505 14170
rect 2505 14118 2551 14170
rect 2255 14116 2311 14118
rect 2335 14116 2391 14118
rect 2415 14116 2471 14118
rect 2495 14116 2551 14118
rect 4106 13626 4162 13628
rect 4186 13626 4242 13628
rect 4266 13626 4322 13628
rect 4346 13626 4402 13628
rect 4106 13574 4152 13626
rect 4152 13574 4162 13626
rect 4186 13574 4216 13626
rect 4216 13574 4228 13626
rect 4228 13574 4242 13626
rect 4266 13574 4280 13626
rect 4280 13574 4292 13626
rect 4292 13574 4322 13626
rect 4346 13574 4356 13626
rect 4356 13574 4402 13626
rect 4106 13572 4162 13574
rect 4186 13572 4242 13574
rect 4266 13572 4322 13574
rect 4346 13572 4402 13574
rect 2255 13082 2311 13084
rect 2335 13082 2391 13084
rect 2415 13082 2471 13084
rect 2495 13082 2551 13084
rect 2255 13030 2301 13082
rect 2301 13030 2311 13082
rect 2335 13030 2365 13082
rect 2365 13030 2377 13082
rect 2377 13030 2391 13082
rect 2415 13030 2429 13082
rect 2429 13030 2441 13082
rect 2441 13030 2471 13082
rect 2495 13030 2505 13082
rect 2505 13030 2551 13082
rect 2255 13028 2311 13030
rect 2335 13028 2391 13030
rect 2415 13028 2471 13030
rect 2495 13028 2551 13030
rect 2255 11994 2311 11996
rect 2335 11994 2391 11996
rect 2415 11994 2471 11996
rect 2495 11994 2551 11996
rect 2255 11942 2301 11994
rect 2301 11942 2311 11994
rect 2335 11942 2365 11994
rect 2365 11942 2377 11994
rect 2377 11942 2391 11994
rect 2415 11942 2429 11994
rect 2429 11942 2441 11994
rect 2441 11942 2471 11994
rect 2495 11942 2505 11994
rect 2505 11942 2551 11994
rect 2255 11940 2311 11942
rect 2335 11940 2391 11942
rect 2415 11940 2471 11942
rect 2495 11940 2551 11942
rect 4106 12538 4162 12540
rect 4186 12538 4242 12540
rect 4266 12538 4322 12540
rect 4346 12538 4402 12540
rect 4106 12486 4152 12538
rect 4152 12486 4162 12538
rect 4186 12486 4216 12538
rect 4216 12486 4228 12538
rect 4228 12486 4242 12538
rect 4266 12486 4280 12538
rect 4280 12486 4292 12538
rect 4292 12486 4322 12538
rect 4346 12486 4356 12538
rect 4356 12486 4402 12538
rect 4106 12484 4162 12486
rect 4186 12484 4242 12486
rect 4266 12484 4322 12486
rect 4346 12484 4402 12486
rect 4106 11450 4162 11452
rect 4186 11450 4242 11452
rect 4266 11450 4322 11452
rect 4346 11450 4402 11452
rect 4106 11398 4152 11450
rect 4152 11398 4162 11450
rect 4186 11398 4216 11450
rect 4216 11398 4228 11450
rect 4228 11398 4242 11450
rect 4266 11398 4280 11450
rect 4280 11398 4292 11450
rect 4292 11398 4322 11450
rect 4346 11398 4356 11450
rect 4356 11398 4402 11450
rect 4106 11396 4162 11398
rect 4186 11396 4242 11398
rect 4266 11396 4322 11398
rect 4346 11396 4402 11398
rect 2255 10906 2311 10908
rect 2335 10906 2391 10908
rect 2415 10906 2471 10908
rect 2495 10906 2551 10908
rect 2255 10854 2301 10906
rect 2301 10854 2311 10906
rect 2335 10854 2365 10906
rect 2365 10854 2377 10906
rect 2377 10854 2391 10906
rect 2415 10854 2429 10906
rect 2429 10854 2441 10906
rect 2441 10854 2471 10906
rect 2495 10854 2505 10906
rect 2505 10854 2551 10906
rect 2255 10852 2311 10854
rect 2335 10852 2391 10854
rect 2415 10852 2471 10854
rect 2495 10852 2551 10854
rect 4106 10362 4162 10364
rect 4186 10362 4242 10364
rect 4266 10362 4322 10364
rect 4346 10362 4402 10364
rect 4106 10310 4152 10362
rect 4152 10310 4162 10362
rect 4186 10310 4216 10362
rect 4216 10310 4228 10362
rect 4228 10310 4242 10362
rect 4266 10310 4280 10362
rect 4280 10310 4292 10362
rect 4292 10310 4322 10362
rect 4346 10310 4356 10362
rect 4356 10310 4402 10362
rect 4106 10308 4162 10310
rect 4186 10308 4242 10310
rect 4266 10308 4322 10310
rect 4346 10308 4402 10310
rect 2255 9818 2311 9820
rect 2335 9818 2391 9820
rect 2415 9818 2471 9820
rect 2495 9818 2551 9820
rect 2255 9766 2301 9818
rect 2301 9766 2311 9818
rect 2335 9766 2365 9818
rect 2365 9766 2377 9818
rect 2377 9766 2391 9818
rect 2415 9766 2429 9818
rect 2429 9766 2441 9818
rect 2441 9766 2471 9818
rect 2495 9766 2505 9818
rect 2505 9766 2551 9818
rect 2255 9764 2311 9766
rect 2335 9764 2391 9766
rect 2415 9764 2471 9766
rect 2495 9764 2551 9766
rect 5957 15258 6013 15260
rect 6037 15258 6093 15260
rect 6117 15258 6173 15260
rect 6197 15258 6253 15260
rect 5957 15206 6003 15258
rect 6003 15206 6013 15258
rect 6037 15206 6067 15258
rect 6067 15206 6079 15258
rect 6079 15206 6093 15258
rect 6117 15206 6131 15258
rect 6131 15206 6143 15258
rect 6143 15206 6173 15258
rect 6197 15206 6207 15258
rect 6207 15206 6253 15258
rect 5957 15204 6013 15206
rect 6037 15204 6093 15206
rect 6117 15204 6173 15206
rect 6197 15204 6253 15206
rect 9659 15258 9715 15260
rect 9739 15258 9795 15260
rect 9819 15258 9875 15260
rect 9899 15258 9955 15260
rect 9659 15206 9705 15258
rect 9705 15206 9715 15258
rect 9739 15206 9769 15258
rect 9769 15206 9781 15258
rect 9781 15206 9795 15258
rect 9819 15206 9833 15258
rect 9833 15206 9845 15258
rect 9845 15206 9875 15258
rect 9899 15206 9909 15258
rect 9909 15206 9955 15258
rect 9659 15204 9715 15206
rect 9739 15204 9795 15206
rect 9819 15204 9875 15206
rect 9899 15204 9955 15206
rect 5957 14170 6013 14172
rect 6037 14170 6093 14172
rect 6117 14170 6173 14172
rect 6197 14170 6253 14172
rect 5957 14118 6003 14170
rect 6003 14118 6013 14170
rect 6037 14118 6067 14170
rect 6067 14118 6079 14170
rect 6079 14118 6093 14170
rect 6117 14118 6131 14170
rect 6131 14118 6143 14170
rect 6143 14118 6173 14170
rect 6197 14118 6207 14170
rect 6207 14118 6253 14170
rect 5957 14116 6013 14118
rect 6037 14116 6093 14118
rect 6117 14116 6173 14118
rect 6197 14116 6253 14118
rect 5957 13082 6013 13084
rect 6037 13082 6093 13084
rect 6117 13082 6173 13084
rect 6197 13082 6253 13084
rect 5957 13030 6003 13082
rect 6003 13030 6013 13082
rect 6037 13030 6067 13082
rect 6067 13030 6079 13082
rect 6079 13030 6093 13082
rect 6117 13030 6131 13082
rect 6131 13030 6143 13082
rect 6143 13030 6173 13082
rect 6197 13030 6207 13082
rect 6207 13030 6253 13082
rect 5957 13028 6013 13030
rect 6037 13028 6093 13030
rect 6117 13028 6173 13030
rect 6197 13028 6253 13030
rect 5957 11994 6013 11996
rect 6037 11994 6093 11996
rect 6117 11994 6173 11996
rect 6197 11994 6253 11996
rect 5957 11942 6003 11994
rect 6003 11942 6013 11994
rect 6037 11942 6067 11994
rect 6067 11942 6079 11994
rect 6079 11942 6093 11994
rect 6117 11942 6131 11994
rect 6131 11942 6143 11994
rect 6143 11942 6173 11994
rect 6197 11942 6207 11994
rect 6207 11942 6253 11994
rect 5957 11940 6013 11942
rect 6037 11940 6093 11942
rect 6117 11940 6173 11942
rect 6197 11940 6253 11942
rect 5957 10906 6013 10908
rect 6037 10906 6093 10908
rect 6117 10906 6173 10908
rect 6197 10906 6253 10908
rect 5957 10854 6003 10906
rect 6003 10854 6013 10906
rect 6037 10854 6067 10906
rect 6067 10854 6079 10906
rect 6079 10854 6093 10906
rect 6117 10854 6131 10906
rect 6131 10854 6143 10906
rect 6143 10854 6173 10906
rect 6197 10854 6207 10906
rect 6207 10854 6253 10906
rect 5957 10852 6013 10854
rect 6037 10852 6093 10854
rect 6117 10852 6173 10854
rect 6197 10852 6253 10854
rect 7808 14714 7864 14716
rect 7888 14714 7944 14716
rect 7968 14714 8024 14716
rect 8048 14714 8104 14716
rect 7808 14662 7854 14714
rect 7854 14662 7864 14714
rect 7888 14662 7918 14714
rect 7918 14662 7930 14714
rect 7930 14662 7944 14714
rect 7968 14662 7982 14714
rect 7982 14662 7994 14714
rect 7994 14662 8024 14714
rect 8048 14662 8058 14714
rect 8058 14662 8104 14714
rect 7808 14660 7864 14662
rect 7888 14660 7944 14662
rect 7968 14660 8024 14662
rect 8048 14660 8104 14662
rect 7808 13626 7864 13628
rect 7888 13626 7944 13628
rect 7968 13626 8024 13628
rect 8048 13626 8104 13628
rect 7808 13574 7854 13626
rect 7854 13574 7864 13626
rect 7888 13574 7918 13626
rect 7918 13574 7930 13626
rect 7930 13574 7944 13626
rect 7968 13574 7982 13626
rect 7982 13574 7994 13626
rect 7994 13574 8024 13626
rect 8048 13574 8058 13626
rect 8058 13574 8104 13626
rect 7808 13572 7864 13574
rect 7888 13572 7944 13574
rect 7968 13572 8024 13574
rect 8048 13572 8104 13574
rect 7808 12538 7864 12540
rect 7888 12538 7944 12540
rect 7968 12538 8024 12540
rect 8048 12538 8104 12540
rect 7808 12486 7854 12538
rect 7854 12486 7864 12538
rect 7888 12486 7918 12538
rect 7918 12486 7930 12538
rect 7930 12486 7944 12538
rect 7968 12486 7982 12538
rect 7982 12486 7994 12538
rect 7994 12486 8024 12538
rect 8048 12486 8058 12538
rect 8058 12486 8104 12538
rect 7808 12484 7864 12486
rect 7888 12484 7944 12486
rect 7968 12484 8024 12486
rect 8048 12484 8104 12486
rect 4106 9274 4162 9276
rect 4186 9274 4242 9276
rect 4266 9274 4322 9276
rect 4346 9274 4402 9276
rect 4106 9222 4152 9274
rect 4152 9222 4162 9274
rect 4186 9222 4216 9274
rect 4216 9222 4228 9274
rect 4228 9222 4242 9274
rect 4266 9222 4280 9274
rect 4280 9222 4292 9274
rect 4292 9222 4322 9274
rect 4346 9222 4356 9274
rect 4356 9222 4402 9274
rect 4106 9220 4162 9222
rect 4186 9220 4242 9222
rect 4266 9220 4322 9222
rect 4346 9220 4402 9222
rect 5957 9818 6013 9820
rect 6037 9818 6093 9820
rect 6117 9818 6173 9820
rect 6197 9818 6253 9820
rect 5957 9766 6003 9818
rect 6003 9766 6013 9818
rect 6037 9766 6067 9818
rect 6067 9766 6079 9818
rect 6079 9766 6093 9818
rect 6117 9766 6131 9818
rect 6131 9766 6143 9818
rect 6143 9766 6173 9818
rect 6197 9766 6207 9818
rect 6207 9766 6253 9818
rect 5957 9764 6013 9766
rect 6037 9764 6093 9766
rect 6117 9764 6173 9766
rect 6197 9764 6253 9766
rect 2255 8730 2311 8732
rect 2335 8730 2391 8732
rect 2415 8730 2471 8732
rect 2495 8730 2551 8732
rect 2255 8678 2301 8730
rect 2301 8678 2311 8730
rect 2335 8678 2365 8730
rect 2365 8678 2377 8730
rect 2377 8678 2391 8730
rect 2415 8678 2429 8730
rect 2429 8678 2441 8730
rect 2441 8678 2471 8730
rect 2495 8678 2505 8730
rect 2505 8678 2551 8730
rect 2255 8676 2311 8678
rect 2335 8676 2391 8678
rect 2415 8676 2471 8678
rect 2495 8676 2551 8678
rect 4106 8186 4162 8188
rect 4186 8186 4242 8188
rect 4266 8186 4322 8188
rect 4346 8186 4402 8188
rect 4106 8134 4152 8186
rect 4152 8134 4162 8186
rect 4186 8134 4216 8186
rect 4216 8134 4228 8186
rect 4228 8134 4242 8186
rect 4266 8134 4280 8186
rect 4280 8134 4292 8186
rect 4292 8134 4322 8186
rect 4346 8134 4356 8186
rect 4356 8134 4402 8186
rect 4106 8132 4162 8134
rect 4186 8132 4242 8134
rect 4266 8132 4322 8134
rect 4346 8132 4402 8134
rect 2255 7642 2311 7644
rect 2335 7642 2391 7644
rect 2415 7642 2471 7644
rect 2495 7642 2551 7644
rect 2255 7590 2301 7642
rect 2301 7590 2311 7642
rect 2335 7590 2365 7642
rect 2365 7590 2377 7642
rect 2377 7590 2391 7642
rect 2415 7590 2429 7642
rect 2429 7590 2441 7642
rect 2441 7590 2471 7642
rect 2495 7590 2505 7642
rect 2505 7590 2551 7642
rect 2255 7588 2311 7590
rect 2335 7588 2391 7590
rect 2415 7588 2471 7590
rect 2495 7588 2551 7590
rect 4106 7098 4162 7100
rect 4186 7098 4242 7100
rect 4266 7098 4322 7100
rect 4346 7098 4402 7100
rect 4106 7046 4152 7098
rect 4152 7046 4162 7098
rect 4186 7046 4216 7098
rect 4216 7046 4228 7098
rect 4228 7046 4242 7098
rect 4266 7046 4280 7098
rect 4280 7046 4292 7098
rect 4292 7046 4322 7098
rect 4346 7046 4356 7098
rect 4356 7046 4402 7098
rect 4106 7044 4162 7046
rect 4186 7044 4242 7046
rect 4266 7044 4322 7046
rect 4346 7044 4402 7046
rect 2255 6554 2311 6556
rect 2335 6554 2391 6556
rect 2415 6554 2471 6556
rect 2495 6554 2551 6556
rect 2255 6502 2301 6554
rect 2301 6502 2311 6554
rect 2335 6502 2365 6554
rect 2365 6502 2377 6554
rect 2377 6502 2391 6554
rect 2415 6502 2429 6554
rect 2429 6502 2441 6554
rect 2441 6502 2471 6554
rect 2495 6502 2505 6554
rect 2505 6502 2551 6554
rect 2255 6500 2311 6502
rect 2335 6500 2391 6502
rect 2415 6500 2471 6502
rect 2495 6500 2551 6502
rect 4106 6010 4162 6012
rect 4186 6010 4242 6012
rect 4266 6010 4322 6012
rect 4346 6010 4402 6012
rect 4106 5958 4152 6010
rect 4152 5958 4162 6010
rect 4186 5958 4216 6010
rect 4216 5958 4228 6010
rect 4228 5958 4242 6010
rect 4266 5958 4280 6010
rect 4280 5958 4292 6010
rect 4292 5958 4322 6010
rect 4346 5958 4356 6010
rect 4356 5958 4402 6010
rect 4106 5956 4162 5958
rect 4186 5956 4242 5958
rect 4266 5956 4322 5958
rect 4346 5956 4402 5958
rect 2255 5466 2311 5468
rect 2335 5466 2391 5468
rect 2415 5466 2471 5468
rect 2495 5466 2551 5468
rect 2255 5414 2301 5466
rect 2301 5414 2311 5466
rect 2335 5414 2365 5466
rect 2365 5414 2377 5466
rect 2377 5414 2391 5466
rect 2415 5414 2429 5466
rect 2429 5414 2441 5466
rect 2441 5414 2471 5466
rect 2495 5414 2505 5466
rect 2505 5414 2551 5466
rect 2255 5412 2311 5414
rect 2335 5412 2391 5414
rect 2415 5412 2471 5414
rect 2495 5412 2551 5414
rect 4106 4922 4162 4924
rect 4186 4922 4242 4924
rect 4266 4922 4322 4924
rect 4346 4922 4402 4924
rect 4106 4870 4152 4922
rect 4152 4870 4162 4922
rect 4186 4870 4216 4922
rect 4216 4870 4228 4922
rect 4228 4870 4242 4922
rect 4266 4870 4280 4922
rect 4280 4870 4292 4922
rect 4292 4870 4322 4922
rect 4346 4870 4356 4922
rect 4356 4870 4402 4922
rect 4106 4868 4162 4870
rect 4186 4868 4242 4870
rect 4266 4868 4322 4870
rect 4346 4868 4402 4870
rect 2255 4378 2311 4380
rect 2335 4378 2391 4380
rect 2415 4378 2471 4380
rect 2495 4378 2551 4380
rect 2255 4326 2301 4378
rect 2301 4326 2311 4378
rect 2335 4326 2365 4378
rect 2365 4326 2377 4378
rect 2377 4326 2391 4378
rect 2415 4326 2429 4378
rect 2429 4326 2441 4378
rect 2441 4326 2471 4378
rect 2495 4326 2505 4378
rect 2505 4326 2551 4378
rect 2255 4324 2311 4326
rect 2335 4324 2391 4326
rect 2415 4324 2471 4326
rect 2495 4324 2551 4326
rect 5957 8730 6013 8732
rect 6037 8730 6093 8732
rect 6117 8730 6173 8732
rect 6197 8730 6253 8732
rect 5957 8678 6003 8730
rect 6003 8678 6013 8730
rect 6037 8678 6067 8730
rect 6067 8678 6079 8730
rect 6079 8678 6093 8730
rect 6117 8678 6131 8730
rect 6131 8678 6143 8730
rect 6143 8678 6173 8730
rect 6197 8678 6207 8730
rect 6207 8678 6253 8730
rect 5957 8676 6013 8678
rect 6037 8676 6093 8678
rect 6117 8676 6173 8678
rect 6197 8676 6253 8678
rect 7808 11450 7864 11452
rect 7888 11450 7944 11452
rect 7968 11450 8024 11452
rect 8048 11450 8104 11452
rect 7808 11398 7854 11450
rect 7854 11398 7864 11450
rect 7888 11398 7918 11450
rect 7918 11398 7930 11450
rect 7930 11398 7944 11450
rect 7968 11398 7982 11450
rect 7982 11398 7994 11450
rect 7994 11398 8024 11450
rect 8048 11398 8058 11450
rect 8058 11398 8104 11450
rect 7808 11396 7864 11398
rect 7888 11396 7944 11398
rect 7968 11396 8024 11398
rect 8048 11396 8104 11398
rect 5957 7642 6013 7644
rect 6037 7642 6093 7644
rect 6117 7642 6173 7644
rect 6197 7642 6253 7644
rect 5957 7590 6003 7642
rect 6003 7590 6013 7642
rect 6037 7590 6067 7642
rect 6067 7590 6079 7642
rect 6079 7590 6093 7642
rect 6117 7590 6131 7642
rect 6131 7590 6143 7642
rect 6143 7590 6173 7642
rect 6197 7590 6207 7642
rect 6207 7590 6253 7642
rect 5957 7588 6013 7590
rect 6037 7588 6093 7590
rect 6117 7588 6173 7590
rect 6197 7588 6253 7590
rect 7808 10362 7864 10364
rect 7888 10362 7944 10364
rect 7968 10362 8024 10364
rect 8048 10362 8104 10364
rect 7808 10310 7854 10362
rect 7854 10310 7864 10362
rect 7888 10310 7918 10362
rect 7918 10310 7930 10362
rect 7930 10310 7944 10362
rect 7968 10310 7982 10362
rect 7982 10310 7994 10362
rect 7994 10310 8024 10362
rect 8048 10310 8058 10362
rect 8058 10310 8104 10362
rect 7808 10308 7864 10310
rect 7888 10308 7944 10310
rect 7968 10308 8024 10310
rect 8048 10308 8104 10310
rect 7808 9274 7864 9276
rect 7888 9274 7944 9276
rect 7968 9274 8024 9276
rect 8048 9274 8104 9276
rect 7808 9222 7854 9274
rect 7854 9222 7864 9274
rect 7888 9222 7918 9274
rect 7918 9222 7930 9274
rect 7930 9222 7944 9274
rect 7968 9222 7982 9274
rect 7982 9222 7994 9274
rect 7994 9222 8024 9274
rect 8048 9222 8058 9274
rect 8058 9222 8104 9274
rect 7808 9220 7864 9222
rect 7888 9220 7944 9222
rect 7968 9220 8024 9222
rect 8048 9220 8104 9222
rect 5957 6554 6013 6556
rect 6037 6554 6093 6556
rect 6117 6554 6173 6556
rect 6197 6554 6253 6556
rect 5957 6502 6003 6554
rect 6003 6502 6013 6554
rect 6037 6502 6067 6554
rect 6067 6502 6079 6554
rect 6079 6502 6093 6554
rect 6117 6502 6131 6554
rect 6131 6502 6143 6554
rect 6143 6502 6173 6554
rect 6197 6502 6207 6554
rect 6207 6502 6253 6554
rect 5957 6500 6013 6502
rect 6037 6500 6093 6502
rect 6117 6500 6173 6502
rect 6197 6500 6253 6502
rect 5957 5466 6013 5468
rect 6037 5466 6093 5468
rect 6117 5466 6173 5468
rect 6197 5466 6253 5468
rect 5957 5414 6003 5466
rect 6003 5414 6013 5466
rect 6037 5414 6067 5466
rect 6067 5414 6079 5466
rect 6079 5414 6093 5466
rect 6117 5414 6131 5466
rect 6131 5414 6143 5466
rect 6143 5414 6173 5466
rect 6197 5414 6207 5466
rect 6207 5414 6253 5466
rect 5957 5412 6013 5414
rect 6037 5412 6093 5414
rect 6117 5412 6173 5414
rect 6197 5412 6253 5414
rect 4106 3834 4162 3836
rect 4186 3834 4242 3836
rect 4266 3834 4322 3836
rect 4346 3834 4402 3836
rect 4106 3782 4152 3834
rect 4152 3782 4162 3834
rect 4186 3782 4216 3834
rect 4216 3782 4228 3834
rect 4228 3782 4242 3834
rect 4266 3782 4280 3834
rect 4280 3782 4292 3834
rect 4292 3782 4322 3834
rect 4346 3782 4356 3834
rect 4356 3782 4402 3834
rect 4106 3780 4162 3782
rect 4186 3780 4242 3782
rect 4266 3780 4322 3782
rect 4346 3780 4402 3782
rect 2255 3290 2311 3292
rect 2335 3290 2391 3292
rect 2415 3290 2471 3292
rect 2495 3290 2551 3292
rect 2255 3238 2301 3290
rect 2301 3238 2311 3290
rect 2335 3238 2365 3290
rect 2365 3238 2377 3290
rect 2377 3238 2391 3290
rect 2415 3238 2429 3290
rect 2429 3238 2441 3290
rect 2441 3238 2471 3290
rect 2495 3238 2505 3290
rect 2505 3238 2551 3290
rect 2255 3236 2311 3238
rect 2335 3236 2391 3238
rect 2415 3236 2471 3238
rect 2495 3236 2551 3238
rect 4106 2746 4162 2748
rect 4186 2746 4242 2748
rect 4266 2746 4322 2748
rect 4346 2746 4402 2748
rect 4106 2694 4152 2746
rect 4152 2694 4162 2746
rect 4186 2694 4216 2746
rect 4216 2694 4228 2746
rect 4228 2694 4242 2746
rect 4266 2694 4280 2746
rect 4280 2694 4292 2746
rect 4292 2694 4322 2746
rect 4346 2694 4356 2746
rect 4356 2694 4402 2746
rect 4106 2692 4162 2694
rect 4186 2692 4242 2694
rect 4266 2692 4322 2694
rect 4346 2692 4402 2694
rect 5957 4378 6013 4380
rect 6037 4378 6093 4380
rect 6117 4378 6173 4380
rect 6197 4378 6253 4380
rect 5957 4326 6003 4378
rect 6003 4326 6013 4378
rect 6037 4326 6067 4378
rect 6067 4326 6079 4378
rect 6079 4326 6093 4378
rect 6117 4326 6131 4378
rect 6131 4326 6143 4378
rect 6143 4326 6173 4378
rect 6197 4326 6207 4378
rect 6207 4326 6253 4378
rect 5957 4324 6013 4326
rect 6037 4324 6093 4326
rect 6117 4324 6173 4326
rect 6197 4324 6253 4326
rect 7808 8186 7864 8188
rect 7888 8186 7944 8188
rect 7968 8186 8024 8188
rect 8048 8186 8104 8188
rect 7808 8134 7854 8186
rect 7854 8134 7864 8186
rect 7888 8134 7918 8186
rect 7918 8134 7930 8186
rect 7930 8134 7944 8186
rect 7968 8134 7982 8186
rect 7982 8134 7994 8186
rect 7994 8134 8024 8186
rect 8048 8134 8058 8186
rect 8058 8134 8104 8186
rect 7808 8132 7864 8134
rect 7888 8132 7944 8134
rect 7968 8132 8024 8134
rect 8048 8132 8104 8134
rect 9659 14170 9715 14172
rect 9739 14170 9795 14172
rect 9819 14170 9875 14172
rect 9899 14170 9955 14172
rect 9659 14118 9705 14170
rect 9705 14118 9715 14170
rect 9739 14118 9769 14170
rect 9769 14118 9781 14170
rect 9781 14118 9795 14170
rect 9819 14118 9833 14170
rect 9833 14118 9845 14170
rect 9845 14118 9875 14170
rect 9899 14118 9909 14170
rect 9909 14118 9955 14170
rect 9659 14116 9715 14118
rect 9739 14116 9795 14118
rect 9819 14116 9875 14118
rect 9899 14116 9955 14118
rect 9659 13082 9715 13084
rect 9739 13082 9795 13084
rect 9819 13082 9875 13084
rect 9899 13082 9955 13084
rect 9659 13030 9705 13082
rect 9705 13030 9715 13082
rect 9739 13030 9769 13082
rect 9769 13030 9781 13082
rect 9781 13030 9795 13082
rect 9819 13030 9833 13082
rect 9833 13030 9845 13082
rect 9845 13030 9875 13082
rect 9899 13030 9909 13082
rect 9909 13030 9955 13082
rect 9659 13028 9715 13030
rect 9739 13028 9795 13030
rect 9819 13028 9875 13030
rect 9899 13028 9955 13030
rect 13361 15258 13417 15260
rect 13441 15258 13497 15260
rect 13521 15258 13577 15260
rect 13601 15258 13657 15260
rect 13361 15206 13407 15258
rect 13407 15206 13417 15258
rect 13441 15206 13471 15258
rect 13471 15206 13483 15258
rect 13483 15206 13497 15258
rect 13521 15206 13535 15258
rect 13535 15206 13547 15258
rect 13547 15206 13577 15258
rect 13601 15206 13611 15258
rect 13611 15206 13657 15258
rect 13361 15204 13417 15206
rect 13441 15204 13497 15206
rect 13521 15204 13577 15206
rect 13601 15204 13657 15206
rect 11510 14714 11566 14716
rect 11590 14714 11646 14716
rect 11670 14714 11726 14716
rect 11750 14714 11806 14716
rect 11510 14662 11556 14714
rect 11556 14662 11566 14714
rect 11590 14662 11620 14714
rect 11620 14662 11632 14714
rect 11632 14662 11646 14714
rect 11670 14662 11684 14714
rect 11684 14662 11696 14714
rect 11696 14662 11726 14714
rect 11750 14662 11760 14714
rect 11760 14662 11806 14714
rect 11510 14660 11566 14662
rect 11590 14660 11646 14662
rect 11670 14660 11726 14662
rect 11750 14660 11806 14662
rect 9659 11994 9715 11996
rect 9739 11994 9795 11996
rect 9819 11994 9875 11996
rect 9899 11994 9955 11996
rect 9659 11942 9705 11994
rect 9705 11942 9715 11994
rect 9739 11942 9769 11994
rect 9769 11942 9781 11994
rect 9781 11942 9795 11994
rect 9819 11942 9833 11994
rect 9833 11942 9845 11994
rect 9845 11942 9875 11994
rect 9899 11942 9909 11994
rect 9909 11942 9955 11994
rect 9659 11940 9715 11942
rect 9739 11940 9795 11942
rect 9819 11940 9875 11942
rect 9899 11940 9955 11942
rect 9659 10906 9715 10908
rect 9739 10906 9795 10908
rect 9819 10906 9875 10908
rect 9899 10906 9955 10908
rect 9659 10854 9705 10906
rect 9705 10854 9715 10906
rect 9739 10854 9769 10906
rect 9769 10854 9781 10906
rect 9781 10854 9795 10906
rect 9819 10854 9833 10906
rect 9833 10854 9845 10906
rect 9845 10854 9875 10906
rect 9899 10854 9909 10906
rect 9909 10854 9955 10906
rect 9659 10852 9715 10854
rect 9739 10852 9795 10854
rect 9819 10852 9875 10854
rect 9899 10852 9955 10854
rect 7808 7098 7864 7100
rect 7888 7098 7944 7100
rect 7968 7098 8024 7100
rect 8048 7098 8104 7100
rect 7808 7046 7854 7098
rect 7854 7046 7864 7098
rect 7888 7046 7918 7098
rect 7918 7046 7930 7098
rect 7930 7046 7944 7098
rect 7968 7046 7982 7098
rect 7982 7046 7994 7098
rect 7994 7046 8024 7098
rect 8048 7046 8058 7098
rect 8058 7046 8104 7098
rect 7808 7044 7864 7046
rect 7888 7044 7944 7046
rect 7968 7044 8024 7046
rect 8048 7044 8104 7046
rect 7470 6160 7526 6216
rect 7746 6160 7802 6216
rect 7808 6010 7864 6012
rect 7888 6010 7944 6012
rect 7968 6010 8024 6012
rect 8048 6010 8104 6012
rect 7808 5958 7854 6010
rect 7854 5958 7864 6010
rect 7888 5958 7918 6010
rect 7918 5958 7930 6010
rect 7930 5958 7944 6010
rect 7968 5958 7982 6010
rect 7982 5958 7994 6010
rect 7994 5958 8024 6010
rect 8048 5958 8058 6010
rect 8058 5958 8104 6010
rect 7808 5956 7864 5958
rect 7888 5956 7944 5958
rect 7968 5956 8024 5958
rect 8048 5956 8104 5958
rect 9659 9818 9715 9820
rect 9739 9818 9795 9820
rect 9819 9818 9875 9820
rect 9899 9818 9955 9820
rect 9659 9766 9705 9818
rect 9705 9766 9715 9818
rect 9739 9766 9769 9818
rect 9769 9766 9781 9818
rect 9781 9766 9795 9818
rect 9819 9766 9833 9818
rect 9833 9766 9845 9818
rect 9845 9766 9875 9818
rect 9899 9766 9909 9818
rect 9909 9766 9955 9818
rect 9659 9764 9715 9766
rect 9739 9764 9795 9766
rect 9819 9764 9875 9766
rect 9899 9764 9955 9766
rect 9659 8730 9715 8732
rect 9739 8730 9795 8732
rect 9819 8730 9875 8732
rect 9899 8730 9955 8732
rect 9659 8678 9705 8730
rect 9705 8678 9715 8730
rect 9739 8678 9769 8730
rect 9769 8678 9781 8730
rect 9781 8678 9795 8730
rect 9819 8678 9833 8730
rect 9833 8678 9845 8730
rect 9845 8678 9875 8730
rect 9899 8678 9909 8730
rect 9909 8678 9955 8730
rect 9659 8676 9715 8678
rect 9739 8676 9795 8678
rect 9819 8676 9875 8678
rect 9899 8676 9955 8678
rect 9659 7642 9715 7644
rect 9739 7642 9795 7644
rect 9819 7642 9875 7644
rect 9899 7642 9955 7644
rect 9659 7590 9705 7642
rect 9705 7590 9715 7642
rect 9739 7590 9769 7642
rect 9769 7590 9781 7642
rect 9781 7590 9795 7642
rect 9819 7590 9833 7642
rect 9833 7590 9845 7642
rect 9845 7590 9875 7642
rect 9899 7590 9909 7642
rect 9909 7590 9955 7642
rect 9659 7588 9715 7590
rect 9739 7588 9795 7590
rect 9819 7588 9875 7590
rect 9899 7588 9955 7590
rect 11242 9424 11298 9480
rect 9659 6554 9715 6556
rect 9739 6554 9795 6556
rect 9819 6554 9875 6556
rect 9899 6554 9955 6556
rect 9659 6502 9705 6554
rect 9705 6502 9715 6554
rect 9739 6502 9769 6554
rect 9769 6502 9781 6554
rect 9781 6502 9795 6554
rect 9819 6502 9833 6554
rect 9833 6502 9845 6554
rect 9845 6502 9875 6554
rect 9899 6502 9909 6554
rect 9909 6502 9955 6554
rect 9659 6500 9715 6502
rect 9739 6500 9795 6502
rect 9819 6500 9875 6502
rect 9899 6500 9955 6502
rect 9659 5466 9715 5468
rect 9739 5466 9795 5468
rect 9819 5466 9875 5468
rect 9899 5466 9955 5468
rect 9659 5414 9705 5466
rect 9705 5414 9715 5466
rect 9739 5414 9769 5466
rect 9769 5414 9781 5466
rect 9781 5414 9795 5466
rect 9819 5414 9833 5466
rect 9833 5414 9845 5466
rect 9845 5414 9875 5466
rect 9899 5414 9909 5466
rect 9909 5414 9955 5466
rect 9659 5412 9715 5414
rect 9739 5412 9795 5414
rect 9819 5412 9875 5414
rect 9899 5412 9955 5414
rect 7808 4922 7864 4924
rect 7888 4922 7944 4924
rect 7968 4922 8024 4924
rect 8048 4922 8104 4924
rect 7808 4870 7854 4922
rect 7854 4870 7864 4922
rect 7888 4870 7918 4922
rect 7918 4870 7930 4922
rect 7930 4870 7944 4922
rect 7968 4870 7982 4922
rect 7982 4870 7994 4922
rect 7994 4870 8024 4922
rect 8048 4870 8058 4922
rect 8058 4870 8104 4922
rect 7808 4868 7864 4870
rect 7888 4868 7944 4870
rect 7968 4868 8024 4870
rect 8048 4868 8104 4870
rect 7808 3834 7864 3836
rect 7888 3834 7944 3836
rect 7968 3834 8024 3836
rect 8048 3834 8104 3836
rect 7808 3782 7854 3834
rect 7854 3782 7864 3834
rect 7888 3782 7918 3834
rect 7918 3782 7930 3834
rect 7930 3782 7944 3834
rect 7968 3782 7982 3834
rect 7982 3782 7994 3834
rect 7994 3782 8024 3834
rect 8048 3782 8058 3834
rect 8058 3782 8104 3834
rect 7808 3780 7864 3782
rect 7888 3780 7944 3782
rect 7968 3780 8024 3782
rect 8048 3780 8104 3782
rect 5957 3290 6013 3292
rect 6037 3290 6093 3292
rect 6117 3290 6173 3292
rect 6197 3290 6253 3292
rect 5957 3238 6003 3290
rect 6003 3238 6013 3290
rect 6037 3238 6067 3290
rect 6067 3238 6079 3290
rect 6079 3238 6093 3290
rect 6117 3238 6131 3290
rect 6131 3238 6143 3290
rect 6143 3238 6173 3290
rect 6197 3238 6207 3290
rect 6207 3238 6253 3290
rect 5957 3236 6013 3238
rect 6037 3236 6093 3238
rect 6117 3236 6173 3238
rect 6197 3236 6253 3238
rect 9659 4378 9715 4380
rect 9739 4378 9795 4380
rect 9819 4378 9875 4380
rect 9899 4378 9955 4380
rect 9659 4326 9705 4378
rect 9705 4326 9715 4378
rect 9739 4326 9769 4378
rect 9769 4326 9781 4378
rect 9781 4326 9795 4378
rect 9819 4326 9833 4378
rect 9833 4326 9845 4378
rect 9845 4326 9875 4378
rect 9899 4326 9909 4378
rect 9909 4326 9955 4378
rect 9659 4324 9715 4326
rect 9739 4324 9795 4326
rect 9819 4324 9875 4326
rect 9899 4324 9955 4326
rect 10414 4528 10470 4584
rect 12346 13812 12348 13832
rect 12348 13812 12400 13832
rect 12400 13812 12402 13832
rect 11510 13626 11566 13628
rect 11590 13626 11646 13628
rect 11670 13626 11726 13628
rect 11750 13626 11806 13628
rect 11510 13574 11556 13626
rect 11556 13574 11566 13626
rect 11590 13574 11620 13626
rect 11620 13574 11632 13626
rect 11632 13574 11646 13626
rect 11670 13574 11684 13626
rect 11684 13574 11696 13626
rect 11696 13574 11726 13626
rect 11750 13574 11760 13626
rect 11760 13574 11806 13626
rect 11510 13572 11566 13574
rect 11590 13572 11646 13574
rect 11670 13572 11726 13574
rect 11750 13572 11806 13574
rect 11510 12538 11566 12540
rect 11590 12538 11646 12540
rect 11670 12538 11726 12540
rect 11750 12538 11806 12540
rect 11510 12486 11556 12538
rect 11556 12486 11566 12538
rect 11590 12486 11620 12538
rect 11620 12486 11632 12538
rect 11632 12486 11646 12538
rect 11670 12486 11684 12538
rect 11684 12486 11696 12538
rect 11696 12486 11726 12538
rect 11750 12486 11760 12538
rect 11760 12486 11806 12538
rect 11510 12484 11566 12486
rect 11590 12484 11646 12486
rect 11670 12484 11726 12486
rect 11750 12484 11806 12486
rect 11510 11450 11566 11452
rect 11590 11450 11646 11452
rect 11670 11450 11726 11452
rect 11750 11450 11806 11452
rect 11510 11398 11556 11450
rect 11556 11398 11566 11450
rect 11590 11398 11620 11450
rect 11620 11398 11632 11450
rect 11632 11398 11646 11450
rect 11670 11398 11684 11450
rect 11684 11398 11696 11450
rect 11696 11398 11726 11450
rect 11750 11398 11760 11450
rect 11760 11398 11806 11450
rect 11510 11396 11566 11398
rect 11590 11396 11646 11398
rect 11670 11396 11726 11398
rect 11750 11396 11806 11398
rect 11510 10362 11566 10364
rect 11590 10362 11646 10364
rect 11670 10362 11726 10364
rect 11750 10362 11806 10364
rect 11510 10310 11556 10362
rect 11556 10310 11566 10362
rect 11590 10310 11620 10362
rect 11620 10310 11632 10362
rect 11632 10310 11646 10362
rect 11670 10310 11684 10362
rect 11684 10310 11696 10362
rect 11696 10310 11726 10362
rect 11750 10310 11760 10362
rect 11760 10310 11806 10362
rect 11510 10308 11566 10310
rect 11590 10308 11646 10310
rect 11670 10308 11726 10310
rect 11750 10308 11806 10310
rect 12346 13776 12402 13812
rect 13361 14170 13417 14172
rect 13441 14170 13497 14172
rect 13521 14170 13577 14172
rect 13601 14170 13657 14172
rect 13361 14118 13407 14170
rect 13407 14118 13417 14170
rect 13441 14118 13471 14170
rect 13471 14118 13483 14170
rect 13483 14118 13497 14170
rect 13521 14118 13535 14170
rect 13535 14118 13547 14170
rect 13547 14118 13577 14170
rect 13601 14118 13611 14170
rect 13611 14118 13657 14170
rect 13361 14116 13417 14118
rect 13441 14116 13497 14118
rect 13521 14116 13577 14118
rect 13601 14116 13657 14118
rect 11510 9274 11566 9276
rect 11590 9274 11646 9276
rect 11670 9274 11726 9276
rect 11750 9274 11806 9276
rect 11510 9222 11556 9274
rect 11556 9222 11566 9274
rect 11590 9222 11620 9274
rect 11620 9222 11632 9274
rect 11632 9222 11646 9274
rect 11670 9222 11684 9274
rect 11684 9222 11696 9274
rect 11696 9222 11726 9274
rect 11750 9222 11760 9274
rect 11760 9222 11806 9274
rect 11510 9220 11566 9222
rect 11590 9220 11646 9222
rect 11670 9220 11726 9222
rect 11750 9220 11806 9222
rect 12898 10104 12954 10160
rect 12806 9988 12862 10024
rect 12806 9968 12808 9988
rect 12808 9968 12860 9988
rect 12860 9968 12862 9988
rect 11510 8186 11566 8188
rect 11590 8186 11646 8188
rect 11670 8186 11726 8188
rect 11750 8186 11806 8188
rect 11510 8134 11556 8186
rect 11556 8134 11566 8186
rect 11590 8134 11620 8186
rect 11620 8134 11632 8186
rect 11632 8134 11646 8186
rect 11670 8134 11684 8186
rect 11684 8134 11696 8186
rect 11696 8134 11726 8186
rect 11750 8134 11760 8186
rect 11760 8134 11806 8186
rect 11510 8132 11566 8134
rect 11590 8132 11646 8134
rect 11670 8132 11726 8134
rect 11750 8132 11806 8134
rect 11510 7098 11566 7100
rect 11590 7098 11646 7100
rect 11670 7098 11726 7100
rect 11750 7098 11806 7100
rect 11510 7046 11556 7098
rect 11556 7046 11566 7098
rect 11590 7046 11620 7098
rect 11620 7046 11632 7098
rect 11632 7046 11646 7098
rect 11670 7046 11684 7098
rect 11684 7046 11696 7098
rect 11696 7046 11726 7098
rect 11750 7046 11760 7098
rect 11760 7046 11806 7098
rect 11510 7044 11566 7046
rect 11590 7044 11646 7046
rect 11670 7044 11726 7046
rect 11750 7044 11806 7046
rect 13361 13082 13417 13084
rect 13441 13082 13497 13084
rect 13521 13082 13577 13084
rect 13601 13082 13657 13084
rect 13361 13030 13407 13082
rect 13407 13030 13417 13082
rect 13441 13030 13471 13082
rect 13471 13030 13483 13082
rect 13483 13030 13497 13082
rect 13521 13030 13535 13082
rect 13535 13030 13547 13082
rect 13547 13030 13577 13082
rect 13601 13030 13611 13082
rect 13611 13030 13657 13082
rect 13361 13028 13417 13030
rect 13441 13028 13497 13030
rect 13521 13028 13577 13030
rect 13601 13028 13657 13030
rect 14462 13812 14464 13832
rect 14464 13812 14516 13832
rect 14516 13812 14518 13832
rect 14462 13776 14518 13812
rect 13361 11994 13417 11996
rect 13441 11994 13497 11996
rect 13521 11994 13577 11996
rect 13601 11994 13657 11996
rect 13361 11942 13407 11994
rect 13407 11942 13417 11994
rect 13441 11942 13471 11994
rect 13471 11942 13483 11994
rect 13483 11942 13497 11994
rect 13521 11942 13535 11994
rect 13535 11942 13547 11994
rect 13547 11942 13577 11994
rect 13601 11942 13611 11994
rect 13611 11942 13657 11994
rect 13361 11940 13417 11942
rect 13441 11940 13497 11942
rect 13521 11940 13577 11942
rect 13601 11940 13657 11942
rect 13361 10906 13417 10908
rect 13441 10906 13497 10908
rect 13521 10906 13577 10908
rect 13601 10906 13657 10908
rect 13361 10854 13407 10906
rect 13407 10854 13417 10906
rect 13441 10854 13471 10906
rect 13471 10854 13483 10906
rect 13483 10854 13497 10906
rect 13521 10854 13535 10906
rect 13535 10854 13547 10906
rect 13547 10854 13577 10906
rect 13601 10854 13611 10906
rect 13611 10854 13657 10906
rect 13361 10852 13417 10854
rect 13441 10852 13497 10854
rect 13521 10852 13577 10854
rect 13601 10852 13657 10854
rect 13174 9460 13176 9480
rect 13176 9460 13228 9480
rect 13228 9460 13230 9480
rect 13174 9424 13230 9460
rect 13450 9968 13506 10024
rect 13361 9818 13417 9820
rect 13441 9818 13497 9820
rect 13521 9818 13577 9820
rect 13601 9818 13657 9820
rect 13361 9766 13407 9818
rect 13407 9766 13417 9818
rect 13441 9766 13471 9818
rect 13471 9766 13483 9818
rect 13483 9766 13497 9818
rect 13521 9766 13535 9818
rect 13535 9766 13547 9818
rect 13547 9766 13577 9818
rect 13601 9766 13611 9818
rect 13611 9766 13657 9818
rect 13361 9764 13417 9766
rect 13441 9764 13497 9766
rect 13521 9764 13577 9766
rect 13601 9764 13657 9766
rect 13361 8730 13417 8732
rect 13441 8730 13497 8732
rect 13521 8730 13577 8732
rect 13601 8730 13657 8732
rect 13361 8678 13407 8730
rect 13407 8678 13417 8730
rect 13441 8678 13471 8730
rect 13471 8678 13483 8730
rect 13483 8678 13497 8730
rect 13521 8678 13535 8730
rect 13535 8678 13547 8730
rect 13547 8678 13577 8730
rect 13601 8678 13611 8730
rect 13611 8678 13657 8730
rect 13361 8676 13417 8678
rect 13441 8676 13497 8678
rect 13521 8676 13577 8678
rect 13601 8676 13657 8678
rect 13361 7642 13417 7644
rect 13441 7642 13497 7644
rect 13521 7642 13577 7644
rect 13601 7642 13657 7644
rect 13361 7590 13407 7642
rect 13407 7590 13417 7642
rect 13441 7590 13471 7642
rect 13471 7590 13483 7642
rect 13483 7590 13497 7642
rect 13521 7590 13535 7642
rect 13535 7590 13547 7642
rect 13547 7590 13577 7642
rect 13601 7590 13611 7642
rect 13611 7590 13657 7642
rect 13361 7588 13417 7590
rect 13441 7588 13497 7590
rect 13521 7588 13577 7590
rect 13601 7588 13657 7590
rect 11510 6010 11566 6012
rect 11590 6010 11646 6012
rect 11670 6010 11726 6012
rect 11750 6010 11806 6012
rect 11510 5958 11556 6010
rect 11556 5958 11566 6010
rect 11590 5958 11620 6010
rect 11620 5958 11632 6010
rect 11632 5958 11646 6010
rect 11670 5958 11684 6010
rect 11684 5958 11696 6010
rect 11696 5958 11726 6010
rect 11750 5958 11760 6010
rect 11760 5958 11806 6010
rect 11510 5956 11566 5958
rect 11590 5956 11646 5958
rect 11670 5956 11726 5958
rect 11750 5956 11806 5958
rect 10874 5072 10930 5128
rect 11886 5108 11888 5128
rect 11888 5108 11940 5128
rect 11940 5108 11942 5128
rect 11886 5072 11942 5108
rect 11510 4922 11566 4924
rect 11590 4922 11646 4924
rect 11670 4922 11726 4924
rect 11750 4922 11806 4924
rect 11510 4870 11556 4922
rect 11556 4870 11566 4922
rect 11590 4870 11620 4922
rect 11620 4870 11632 4922
rect 11632 4870 11646 4922
rect 11670 4870 11684 4922
rect 11684 4870 11696 4922
rect 11696 4870 11726 4922
rect 11750 4870 11760 4922
rect 11760 4870 11806 4922
rect 11510 4868 11566 4870
rect 11590 4868 11646 4870
rect 11670 4868 11726 4870
rect 11750 4868 11806 4870
rect 11518 4548 11574 4584
rect 11518 4528 11520 4548
rect 11520 4528 11572 4548
rect 11572 4528 11574 4548
rect 9659 3290 9715 3292
rect 9739 3290 9795 3292
rect 9819 3290 9875 3292
rect 9899 3290 9955 3292
rect 9659 3238 9705 3290
rect 9705 3238 9715 3290
rect 9739 3238 9769 3290
rect 9769 3238 9781 3290
rect 9781 3238 9795 3290
rect 9819 3238 9833 3290
rect 9833 3238 9845 3290
rect 9845 3238 9875 3290
rect 9899 3238 9909 3290
rect 9909 3238 9955 3290
rect 9659 3236 9715 3238
rect 9739 3236 9795 3238
rect 9819 3236 9875 3238
rect 9899 3236 9955 3238
rect 7808 2746 7864 2748
rect 7888 2746 7944 2748
rect 7968 2746 8024 2748
rect 8048 2746 8104 2748
rect 7808 2694 7854 2746
rect 7854 2694 7864 2746
rect 7888 2694 7918 2746
rect 7918 2694 7930 2746
rect 7930 2694 7944 2746
rect 7968 2694 7982 2746
rect 7982 2694 7994 2746
rect 7994 2694 8024 2746
rect 8048 2694 8058 2746
rect 8058 2694 8104 2746
rect 7808 2692 7864 2694
rect 7888 2692 7944 2694
rect 7968 2692 8024 2694
rect 8048 2692 8104 2694
rect 11510 3834 11566 3836
rect 11590 3834 11646 3836
rect 11670 3834 11726 3836
rect 11750 3834 11806 3836
rect 11510 3782 11556 3834
rect 11556 3782 11566 3834
rect 11590 3782 11620 3834
rect 11620 3782 11632 3834
rect 11632 3782 11646 3834
rect 11670 3782 11684 3834
rect 11684 3782 11696 3834
rect 11696 3782 11726 3834
rect 11750 3782 11760 3834
rect 11760 3782 11806 3834
rect 11510 3780 11566 3782
rect 11590 3780 11646 3782
rect 11670 3780 11726 3782
rect 11750 3780 11806 3782
rect 13361 6554 13417 6556
rect 13441 6554 13497 6556
rect 13521 6554 13577 6556
rect 13601 6554 13657 6556
rect 13361 6502 13407 6554
rect 13407 6502 13417 6554
rect 13441 6502 13471 6554
rect 13471 6502 13483 6554
rect 13483 6502 13497 6554
rect 13521 6502 13535 6554
rect 13535 6502 13547 6554
rect 13547 6502 13577 6554
rect 13601 6502 13611 6554
rect 13611 6502 13657 6554
rect 13361 6500 13417 6502
rect 13441 6500 13497 6502
rect 13521 6500 13577 6502
rect 13601 6500 13657 6502
rect 15212 14714 15268 14716
rect 15292 14714 15348 14716
rect 15372 14714 15428 14716
rect 15452 14714 15508 14716
rect 15212 14662 15258 14714
rect 15258 14662 15268 14714
rect 15292 14662 15322 14714
rect 15322 14662 15334 14714
rect 15334 14662 15348 14714
rect 15372 14662 15386 14714
rect 15386 14662 15398 14714
rect 15398 14662 15428 14714
rect 15452 14662 15462 14714
rect 15462 14662 15508 14714
rect 15212 14660 15268 14662
rect 15292 14660 15348 14662
rect 15372 14660 15428 14662
rect 15452 14660 15508 14662
rect 15106 14456 15162 14512
rect 15212 13626 15268 13628
rect 15292 13626 15348 13628
rect 15372 13626 15428 13628
rect 15452 13626 15508 13628
rect 15212 13574 15258 13626
rect 15258 13574 15268 13626
rect 15292 13574 15322 13626
rect 15322 13574 15334 13626
rect 15334 13574 15348 13626
rect 15372 13574 15386 13626
rect 15386 13574 15398 13626
rect 15398 13574 15428 13626
rect 15452 13574 15462 13626
rect 15462 13574 15508 13626
rect 15212 13572 15268 13574
rect 15292 13572 15348 13574
rect 15372 13572 15428 13574
rect 15452 13572 15508 13574
rect 15212 12538 15268 12540
rect 15292 12538 15348 12540
rect 15372 12538 15428 12540
rect 15452 12538 15508 12540
rect 15212 12486 15258 12538
rect 15258 12486 15268 12538
rect 15292 12486 15322 12538
rect 15322 12486 15334 12538
rect 15334 12486 15348 12538
rect 15372 12486 15386 12538
rect 15386 12486 15398 12538
rect 15398 12486 15428 12538
rect 15452 12486 15462 12538
rect 15462 12486 15508 12538
rect 15212 12484 15268 12486
rect 15292 12484 15348 12486
rect 15372 12484 15428 12486
rect 15452 12484 15508 12486
rect 15106 12316 15108 12336
rect 15108 12316 15160 12336
rect 15160 12316 15162 12336
rect 15106 12280 15162 12316
rect 15212 11450 15268 11452
rect 15292 11450 15348 11452
rect 15372 11450 15428 11452
rect 15452 11450 15508 11452
rect 15212 11398 15258 11450
rect 15258 11398 15268 11450
rect 15292 11398 15322 11450
rect 15322 11398 15334 11450
rect 15334 11398 15348 11450
rect 15372 11398 15386 11450
rect 15386 11398 15398 11450
rect 15398 11398 15428 11450
rect 15452 11398 15462 11450
rect 15462 11398 15508 11450
rect 15212 11396 15268 11398
rect 15292 11396 15348 11398
rect 15372 11396 15428 11398
rect 15452 11396 15508 11398
rect 15106 10648 15162 10704
rect 15212 10362 15268 10364
rect 15292 10362 15348 10364
rect 15372 10362 15428 10364
rect 15452 10362 15508 10364
rect 15212 10310 15258 10362
rect 15258 10310 15268 10362
rect 15292 10310 15322 10362
rect 15322 10310 15334 10362
rect 15334 10310 15348 10362
rect 15372 10310 15386 10362
rect 15386 10310 15398 10362
rect 15398 10310 15428 10362
rect 15452 10310 15462 10362
rect 15462 10310 15508 10362
rect 15212 10308 15268 10310
rect 15292 10308 15348 10310
rect 15372 10308 15428 10310
rect 15452 10308 15508 10310
rect 15106 10104 15162 10160
rect 15212 9274 15268 9276
rect 15292 9274 15348 9276
rect 15372 9274 15428 9276
rect 15452 9274 15508 9276
rect 15212 9222 15258 9274
rect 15258 9222 15268 9274
rect 15292 9222 15322 9274
rect 15322 9222 15334 9274
rect 15334 9222 15348 9274
rect 15372 9222 15386 9274
rect 15386 9222 15398 9274
rect 15398 9222 15428 9274
rect 15452 9222 15462 9274
rect 15462 9222 15508 9274
rect 15212 9220 15268 9222
rect 15292 9220 15348 9222
rect 15372 9220 15428 9222
rect 15452 9220 15508 9222
rect 15106 8744 15162 8800
rect 15212 8186 15268 8188
rect 15292 8186 15348 8188
rect 15372 8186 15428 8188
rect 15452 8186 15508 8188
rect 15212 8134 15258 8186
rect 15258 8134 15268 8186
rect 15292 8134 15322 8186
rect 15322 8134 15334 8186
rect 15334 8134 15348 8186
rect 15372 8134 15386 8186
rect 15386 8134 15398 8186
rect 15398 8134 15428 8186
rect 15452 8134 15462 8186
rect 15462 8134 15508 8186
rect 15212 8132 15268 8134
rect 15292 8132 15348 8134
rect 15372 8132 15428 8134
rect 15452 8132 15508 8134
rect 15014 6840 15070 6896
rect 13361 5466 13417 5468
rect 13441 5466 13497 5468
rect 13521 5466 13577 5468
rect 13601 5466 13657 5468
rect 13361 5414 13407 5466
rect 13407 5414 13417 5466
rect 13441 5414 13471 5466
rect 13471 5414 13483 5466
rect 13483 5414 13497 5466
rect 13521 5414 13535 5466
rect 13535 5414 13547 5466
rect 13547 5414 13577 5466
rect 13601 5414 13611 5466
rect 13611 5414 13657 5466
rect 13361 5412 13417 5414
rect 13441 5412 13497 5414
rect 13521 5412 13577 5414
rect 13601 5412 13657 5414
rect 13361 4378 13417 4380
rect 13441 4378 13497 4380
rect 13521 4378 13577 4380
rect 13601 4378 13657 4380
rect 13361 4326 13407 4378
rect 13407 4326 13417 4378
rect 13441 4326 13471 4378
rect 13471 4326 13483 4378
rect 13483 4326 13497 4378
rect 13521 4326 13535 4378
rect 13535 4326 13547 4378
rect 13547 4326 13577 4378
rect 13601 4326 13611 4378
rect 13611 4326 13657 4378
rect 13361 4324 13417 4326
rect 13441 4324 13497 4326
rect 13521 4324 13577 4326
rect 13601 4324 13657 4326
rect 13361 3290 13417 3292
rect 13441 3290 13497 3292
rect 13521 3290 13577 3292
rect 13601 3290 13657 3292
rect 13361 3238 13407 3290
rect 13407 3238 13417 3290
rect 13441 3238 13471 3290
rect 13471 3238 13483 3290
rect 13483 3238 13497 3290
rect 13521 3238 13535 3290
rect 13535 3238 13547 3290
rect 13547 3238 13577 3290
rect 13601 3238 13611 3290
rect 13611 3238 13657 3290
rect 13361 3236 13417 3238
rect 13441 3236 13497 3238
rect 13521 3236 13577 3238
rect 13601 3236 13657 3238
rect 14462 3032 14518 3088
rect 11510 2746 11566 2748
rect 11590 2746 11646 2748
rect 11670 2746 11726 2748
rect 11750 2746 11806 2748
rect 11510 2694 11556 2746
rect 11556 2694 11566 2746
rect 11590 2694 11620 2746
rect 11620 2694 11632 2746
rect 11632 2694 11646 2746
rect 11670 2694 11684 2746
rect 11684 2694 11696 2746
rect 11696 2694 11726 2746
rect 11750 2694 11760 2746
rect 11760 2694 11806 2746
rect 11510 2692 11566 2694
rect 11590 2692 11646 2694
rect 11670 2692 11726 2694
rect 11750 2692 11806 2694
rect 2255 2202 2311 2204
rect 2335 2202 2391 2204
rect 2415 2202 2471 2204
rect 2495 2202 2551 2204
rect 2255 2150 2301 2202
rect 2301 2150 2311 2202
rect 2335 2150 2365 2202
rect 2365 2150 2377 2202
rect 2377 2150 2391 2202
rect 2415 2150 2429 2202
rect 2429 2150 2441 2202
rect 2441 2150 2471 2202
rect 2495 2150 2505 2202
rect 2505 2150 2551 2202
rect 2255 2148 2311 2150
rect 2335 2148 2391 2150
rect 2415 2148 2471 2150
rect 2495 2148 2551 2150
rect 5957 2202 6013 2204
rect 6037 2202 6093 2204
rect 6117 2202 6173 2204
rect 6197 2202 6253 2204
rect 5957 2150 6003 2202
rect 6003 2150 6013 2202
rect 6037 2150 6067 2202
rect 6067 2150 6079 2202
rect 6079 2150 6093 2202
rect 6117 2150 6131 2202
rect 6131 2150 6143 2202
rect 6143 2150 6173 2202
rect 6197 2150 6207 2202
rect 6207 2150 6253 2202
rect 5957 2148 6013 2150
rect 6037 2148 6093 2150
rect 6117 2148 6173 2150
rect 6197 2148 6253 2150
rect 9659 2202 9715 2204
rect 9739 2202 9795 2204
rect 9819 2202 9875 2204
rect 9899 2202 9955 2204
rect 9659 2150 9705 2202
rect 9705 2150 9715 2202
rect 9739 2150 9769 2202
rect 9769 2150 9781 2202
rect 9781 2150 9795 2202
rect 9819 2150 9833 2202
rect 9833 2150 9845 2202
rect 9845 2150 9875 2202
rect 9899 2150 9909 2202
rect 9909 2150 9955 2202
rect 9659 2148 9715 2150
rect 9739 2148 9795 2150
rect 9819 2148 9875 2150
rect 9899 2148 9955 2150
rect 13361 2202 13417 2204
rect 13441 2202 13497 2204
rect 13521 2202 13577 2204
rect 13601 2202 13657 2204
rect 13361 2150 13407 2202
rect 13407 2150 13417 2202
rect 13441 2150 13471 2202
rect 13471 2150 13483 2202
rect 13483 2150 13497 2202
rect 13521 2150 13535 2202
rect 13535 2150 13547 2202
rect 13547 2150 13577 2202
rect 13601 2150 13611 2202
rect 13611 2150 13657 2202
rect 13361 2148 13417 2150
rect 13441 2148 13497 2150
rect 13521 2148 13577 2150
rect 13601 2148 13657 2150
rect 4106 1658 4162 1660
rect 4186 1658 4242 1660
rect 4266 1658 4322 1660
rect 4346 1658 4402 1660
rect 4106 1606 4152 1658
rect 4152 1606 4162 1658
rect 4186 1606 4216 1658
rect 4216 1606 4228 1658
rect 4228 1606 4242 1658
rect 4266 1606 4280 1658
rect 4280 1606 4292 1658
rect 4292 1606 4322 1658
rect 4346 1606 4356 1658
rect 4356 1606 4402 1658
rect 4106 1604 4162 1606
rect 4186 1604 4242 1606
rect 4266 1604 4322 1606
rect 4346 1604 4402 1606
rect 7808 1658 7864 1660
rect 7888 1658 7944 1660
rect 7968 1658 8024 1660
rect 8048 1658 8104 1660
rect 7808 1606 7854 1658
rect 7854 1606 7864 1658
rect 7888 1606 7918 1658
rect 7918 1606 7930 1658
rect 7930 1606 7944 1658
rect 7968 1606 7982 1658
rect 7982 1606 7994 1658
rect 7994 1606 8024 1658
rect 8048 1606 8058 1658
rect 8058 1606 8104 1658
rect 7808 1604 7864 1606
rect 7888 1604 7944 1606
rect 7968 1604 8024 1606
rect 8048 1604 8104 1606
rect 11510 1658 11566 1660
rect 11590 1658 11646 1660
rect 11670 1658 11726 1660
rect 11750 1658 11806 1660
rect 11510 1606 11556 1658
rect 11556 1606 11566 1658
rect 11590 1606 11620 1658
rect 11620 1606 11632 1658
rect 11632 1606 11646 1658
rect 11670 1606 11684 1658
rect 11684 1606 11696 1658
rect 11696 1606 11726 1658
rect 11750 1606 11760 1658
rect 11760 1606 11806 1658
rect 11510 1604 11566 1606
rect 11590 1604 11646 1606
rect 11670 1604 11726 1606
rect 11750 1604 11806 1606
rect 15212 7098 15268 7100
rect 15292 7098 15348 7100
rect 15372 7098 15428 7100
rect 15452 7098 15508 7100
rect 15212 7046 15258 7098
rect 15258 7046 15268 7098
rect 15292 7046 15322 7098
rect 15322 7046 15334 7098
rect 15334 7046 15348 7098
rect 15372 7046 15386 7098
rect 15386 7046 15398 7098
rect 15398 7046 15428 7098
rect 15452 7046 15462 7098
rect 15462 7046 15508 7098
rect 15212 7044 15268 7046
rect 15292 7044 15348 7046
rect 15372 7044 15428 7046
rect 15452 7044 15508 7046
rect 15212 6010 15268 6012
rect 15292 6010 15348 6012
rect 15372 6010 15428 6012
rect 15452 6010 15508 6012
rect 15212 5958 15258 6010
rect 15258 5958 15268 6010
rect 15292 5958 15322 6010
rect 15322 5958 15334 6010
rect 15334 5958 15348 6010
rect 15372 5958 15386 6010
rect 15386 5958 15398 6010
rect 15398 5958 15428 6010
rect 15452 5958 15462 6010
rect 15462 5958 15508 6010
rect 15212 5956 15268 5958
rect 15292 5956 15348 5958
rect 15372 5956 15428 5958
rect 15452 5956 15508 5958
rect 15106 5480 15162 5536
rect 15212 4922 15268 4924
rect 15292 4922 15348 4924
rect 15372 4922 15428 4924
rect 15452 4922 15508 4924
rect 15212 4870 15258 4922
rect 15258 4870 15268 4922
rect 15292 4870 15322 4922
rect 15322 4870 15334 4922
rect 15334 4870 15348 4922
rect 15372 4870 15386 4922
rect 15386 4870 15398 4922
rect 15398 4870 15428 4922
rect 15452 4870 15462 4922
rect 15462 4870 15508 4922
rect 15212 4868 15268 4870
rect 15292 4868 15348 4870
rect 15372 4868 15428 4870
rect 15452 4868 15508 4870
rect 15212 3834 15268 3836
rect 15292 3834 15348 3836
rect 15372 3834 15428 3836
rect 15452 3834 15508 3836
rect 15212 3782 15258 3834
rect 15258 3782 15268 3834
rect 15292 3782 15322 3834
rect 15322 3782 15334 3834
rect 15334 3782 15348 3834
rect 15372 3782 15386 3834
rect 15386 3782 15398 3834
rect 15398 3782 15428 3834
rect 15452 3782 15462 3834
rect 15462 3782 15508 3834
rect 15212 3780 15268 3782
rect 15292 3780 15348 3782
rect 15372 3780 15428 3782
rect 15452 3780 15508 3782
rect 15212 2746 15268 2748
rect 15292 2746 15348 2748
rect 15372 2746 15428 2748
rect 15452 2746 15508 2748
rect 15212 2694 15258 2746
rect 15258 2694 15268 2746
rect 15292 2694 15322 2746
rect 15322 2694 15334 2746
rect 15334 2694 15348 2746
rect 15372 2694 15386 2746
rect 15386 2694 15398 2746
rect 15398 2694 15428 2746
rect 15452 2694 15462 2746
rect 15462 2694 15508 2746
rect 15212 2692 15268 2694
rect 15292 2692 15348 2694
rect 15372 2692 15428 2694
rect 15452 2692 15508 2694
rect 15212 1658 15268 1660
rect 15292 1658 15348 1660
rect 15372 1658 15428 1660
rect 15452 1658 15508 1660
rect 15212 1606 15258 1658
rect 15258 1606 15268 1658
rect 15292 1606 15322 1658
rect 15322 1606 15334 1658
rect 15334 1606 15348 1658
rect 15372 1606 15386 1658
rect 15386 1606 15398 1658
rect 15398 1606 15428 1658
rect 15452 1606 15462 1658
rect 15462 1606 15508 1658
rect 15212 1604 15268 1606
rect 15292 1604 15348 1606
rect 15372 1604 15428 1606
rect 15452 1604 15508 1606
rect 15014 1128 15070 1184
rect 2255 1114 2311 1116
rect 2335 1114 2391 1116
rect 2415 1114 2471 1116
rect 2495 1114 2551 1116
rect 2255 1062 2301 1114
rect 2301 1062 2311 1114
rect 2335 1062 2365 1114
rect 2365 1062 2377 1114
rect 2377 1062 2391 1114
rect 2415 1062 2429 1114
rect 2429 1062 2441 1114
rect 2441 1062 2471 1114
rect 2495 1062 2505 1114
rect 2505 1062 2551 1114
rect 2255 1060 2311 1062
rect 2335 1060 2391 1062
rect 2415 1060 2471 1062
rect 2495 1060 2551 1062
rect 5957 1114 6013 1116
rect 6037 1114 6093 1116
rect 6117 1114 6173 1116
rect 6197 1114 6253 1116
rect 5957 1062 6003 1114
rect 6003 1062 6013 1114
rect 6037 1062 6067 1114
rect 6067 1062 6079 1114
rect 6079 1062 6093 1114
rect 6117 1062 6131 1114
rect 6131 1062 6143 1114
rect 6143 1062 6173 1114
rect 6197 1062 6207 1114
rect 6207 1062 6253 1114
rect 5957 1060 6013 1062
rect 6037 1060 6093 1062
rect 6117 1060 6173 1062
rect 6197 1060 6253 1062
rect 9659 1114 9715 1116
rect 9739 1114 9795 1116
rect 9819 1114 9875 1116
rect 9899 1114 9955 1116
rect 9659 1062 9705 1114
rect 9705 1062 9715 1114
rect 9739 1062 9769 1114
rect 9769 1062 9781 1114
rect 9781 1062 9795 1114
rect 9819 1062 9833 1114
rect 9833 1062 9845 1114
rect 9845 1062 9875 1114
rect 9899 1062 9909 1114
rect 9909 1062 9955 1114
rect 9659 1060 9715 1062
rect 9739 1060 9795 1062
rect 9819 1060 9875 1062
rect 9899 1060 9955 1062
rect 13361 1114 13417 1116
rect 13441 1114 13497 1116
rect 13521 1114 13577 1116
rect 13601 1114 13657 1116
rect 13361 1062 13407 1114
rect 13407 1062 13417 1114
rect 13441 1062 13471 1114
rect 13471 1062 13483 1114
rect 13483 1062 13497 1114
rect 13521 1062 13535 1114
rect 13535 1062 13547 1114
rect 13547 1062 13577 1114
rect 13601 1062 13611 1114
rect 13611 1062 13657 1114
rect 13361 1060 13417 1062
rect 13441 1060 13497 1062
rect 13521 1060 13577 1062
rect 13601 1060 13657 1062
rect 4106 570 4162 572
rect 4186 570 4242 572
rect 4266 570 4322 572
rect 4346 570 4402 572
rect 4106 518 4152 570
rect 4152 518 4162 570
rect 4186 518 4216 570
rect 4216 518 4228 570
rect 4228 518 4242 570
rect 4266 518 4280 570
rect 4280 518 4292 570
rect 4292 518 4322 570
rect 4346 518 4356 570
rect 4356 518 4402 570
rect 4106 516 4162 518
rect 4186 516 4242 518
rect 4266 516 4322 518
rect 4346 516 4402 518
rect 7808 570 7864 572
rect 7888 570 7944 572
rect 7968 570 8024 572
rect 8048 570 8104 572
rect 7808 518 7854 570
rect 7854 518 7864 570
rect 7888 518 7918 570
rect 7918 518 7930 570
rect 7930 518 7944 570
rect 7968 518 7982 570
rect 7982 518 7994 570
rect 7994 518 8024 570
rect 8048 518 8058 570
rect 8058 518 8104 570
rect 7808 516 7864 518
rect 7888 516 7944 518
rect 7968 516 8024 518
rect 8048 516 8104 518
rect 11510 570 11566 572
rect 11590 570 11646 572
rect 11670 570 11726 572
rect 11750 570 11806 572
rect 11510 518 11556 570
rect 11556 518 11566 570
rect 11590 518 11620 570
rect 11620 518 11632 570
rect 11632 518 11646 570
rect 11670 518 11684 570
rect 11684 518 11696 570
rect 11696 518 11726 570
rect 11750 518 11760 570
rect 11760 518 11806 570
rect 11510 516 11566 518
rect 11590 516 11646 518
rect 11670 516 11726 518
rect 11750 516 11806 518
rect 15212 570 15268 572
rect 15292 570 15348 572
rect 15372 570 15428 572
rect 15452 570 15508 572
rect 15212 518 15258 570
rect 15258 518 15268 570
rect 15292 518 15322 570
rect 15322 518 15334 570
rect 15334 518 15348 570
rect 15372 518 15386 570
rect 15386 518 15398 570
rect 15398 518 15428 570
rect 15452 518 15462 570
rect 15462 518 15508 570
rect 15212 516 15268 518
rect 15292 516 15348 518
rect 15372 516 15428 518
rect 15452 516 15508 518
<< metal3 >>
rect 2245 15264 2561 15265
rect 2245 15200 2251 15264
rect 2315 15200 2331 15264
rect 2395 15200 2411 15264
rect 2475 15200 2491 15264
rect 2555 15200 2561 15264
rect 2245 15199 2561 15200
rect 5947 15264 6263 15265
rect 5947 15200 5953 15264
rect 6017 15200 6033 15264
rect 6097 15200 6113 15264
rect 6177 15200 6193 15264
rect 6257 15200 6263 15264
rect 5947 15199 6263 15200
rect 9649 15264 9965 15265
rect 9649 15200 9655 15264
rect 9719 15200 9735 15264
rect 9799 15200 9815 15264
rect 9879 15200 9895 15264
rect 9959 15200 9965 15264
rect 9649 15199 9965 15200
rect 13351 15264 13667 15265
rect 13351 15200 13357 15264
rect 13421 15200 13437 15264
rect 13501 15200 13517 15264
rect 13581 15200 13597 15264
rect 13661 15200 13667 15264
rect 13351 15199 13667 15200
rect 4096 14720 4412 14721
rect 4096 14656 4102 14720
rect 4166 14656 4182 14720
rect 4246 14656 4262 14720
rect 4326 14656 4342 14720
rect 4406 14656 4412 14720
rect 4096 14655 4412 14656
rect 7798 14720 8114 14721
rect 7798 14656 7804 14720
rect 7868 14656 7884 14720
rect 7948 14656 7964 14720
rect 8028 14656 8044 14720
rect 8108 14656 8114 14720
rect 7798 14655 8114 14656
rect 11500 14720 11816 14721
rect 11500 14656 11506 14720
rect 11570 14656 11586 14720
rect 11650 14656 11666 14720
rect 11730 14656 11746 14720
rect 11810 14656 11816 14720
rect 11500 14655 11816 14656
rect 15202 14720 15518 14721
rect 15202 14656 15208 14720
rect 15272 14656 15288 14720
rect 15352 14656 15368 14720
rect 15432 14656 15448 14720
rect 15512 14656 15518 14720
rect 15202 14655 15518 14656
rect 15101 14514 15167 14517
rect 15600 14514 16000 14544
rect 15101 14512 16000 14514
rect 15101 14456 15106 14512
rect 15162 14456 16000 14512
rect 15101 14454 16000 14456
rect 15101 14451 15167 14454
rect 15600 14424 16000 14454
rect 2245 14176 2561 14177
rect 2245 14112 2251 14176
rect 2315 14112 2331 14176
rect 2395 14112 2411 14176
rect 2475 14112 2491 14176
rect 2555 14112 2561 14176
rect 2245 14111 2561 14112
rect 5947 14176 6263 14177
rect 5947 14112 5953 14176
rect 6017 14112 6033 14176
rect 6097 14112 6113 14176
rect 6177 14112 6193 14176
rect 6257 14112 6263 14176
rect 5947 14111 6263 14112
rect 9649 14176 9965 14177
rect 9649 14112 9655 14176
rect 9719 14112 9735 14176
rect 9799 14112 9815 14176
rect 9879 14112 9895 14176
rect 9959 14112 9965 14176
rect 9649 14111 9965 14112
rect 13351 14176 13667 14177
rect 13351 14112 13357 14176
rect 13421 14112 13437 14176
rect 13501 14112 13517 14176
rect 13581 14112 13597 14176
rect 13661 14112 13667 14176
rect 13351 14111 13667 14112
rect 12341 13834 12407 13837
rect 14457 13834 14523 13837
rect 12341 13832 14523 13834
rect 12341 13776 12346 13832
rect 12402 13776 14462 13832
rect 14518 13776 14523 13832
rect 12341 13774 14523 13776
rect 12341 13771 12407 13774
rect 14457 13771 14523 13774
rect 4096 13632 4412 13633
rect 4096 13568 4102 13632
rect 4166 13568 4182 13632
rect 4246 13568 4262 13632
rect 4326 13568 4342 13632
rect 4406 13568 4412 13632
rect 4096 13567 4412 13568
rect 7798 13632 8114 13633
rect 7798 13568 7804 13632
rect 7868 13568 7884 13632
rect 7948 13568 7964 13632
rect 8028 13568 8044 13632
rect 8108 13568 8114 13632
rect 7798 13567 8114 13568
rect 11500 13632 11816 13633
rect 11500 13568 11506 13632
rect 11570 13568 11586 13632
rect 11650 13568 11666 13632
rect 11730 13568 11746 13632
rect 11810 13568 11816 13632
rect 11500 13567 11816 13568
rect 15202 13632 15518 13633
rect 15202 13568 15208 13632
rect 15272 13568 15288 13632
rect 15352 13568 15368 13632
rect 15432 13568 15448 13632
rect 15512 13568 15518 13632
rect 15202 13567 15518 13568
rect 2245 13088 2561 13089
rect 2245 13024 2251 13088
rect 2315 13024 2331 13088
rect 2395 13024 2411 13088
rect 2475 13024 2491 13088
rect 2555 13024 2561 13088
rect 2245 13023 2561 13024
rect 5947 13088 6263 13089
rect 5947 13024 5953 13088
rect 6017 13024 6033 13088
rect 6097 13024 6113 13088
rect 6177 13024 6193 13088
rect 6257 13024 6263 13088
rect 5947 13023 6263 13024
rect 9649 13088 9965 13089
rect 9649 13024 9655 13088
rect 9719 13024 9735 13088
rect 9799 13024 9815 13088
rect 9879 13024 9895 13088
rect 9959 13024 9965 13088
rect 9649 13023 9965 13024
rect 13351 13088 13667 13089
rect 13351 13024 13357 13088
rect 13421 13024 13437 13088
rect 13501 13024 13517 13088
rect 13581 13024 13597 13088
rect 13661 13024 13667 13088
rect 13351 13023 13667 13024
rect 4096 12544 4412 12545
rect 4096 12480 4102 12544
rect 4166 12480 4182 12544
rect 4246 12480 4262 12544
rect 4326 12480 4342 12544
rect 4406 12480 4412 12544
rect 4096 12479 4412 12480
rect 7798 12544 8114 12545
rect 7798 12480 7804 12544
rect 7868 12480 7884 12544
rect 7948 12480 7964 12544
rect 8028 12480 8044 12544
rect 8108 12480 8114 12544
rect 7798 12479 8114 12480
rect 11500 12544 11816 12545
rect 11500 12480 11506 12544
rect 11570 12480 11586 12544
rect 11650 12480 11666 12544
rect 11730 12480 11746 12544
rect 11810 12480 11816 12544
rect 11500 12479 11816 12480
rect 15202 12544 15518 12545
rect 15202 12480 15208 12544
rect 15272 12480 15288 12544
rect 15352 12480 15368 12544
rect 15432 12480 15448 12544
rect 15512 12480 15518 12544
rect 15600 12520 16000 12640
rect 15202 12479 15518 12480
rect 15101 12338 15167 12341
rect 15702 12338 15762 12520
rect 15101 12336 15762 12338
rect 15101 12280 15106 12336
rect 15162 12280 15762 12336
rect 15101 12278 15762 12280
rect 15101 12275 15167 12278
rect 2245 12000 2561 12001
rect 2245 11936 2251 12000
rect 2315 11936 2331 12000
rect 2395 11936 2411 12000
rect 2475 11936 2491 12000
rect 2555 11936 2561 12000
rect 2245 11935 2561 11936
rect 5947 12000 6263 12001
rect 5947 11936 5953 12000
rect 6017 11936 6033 12000
rect 6097 11936 6113 12000
rect 6177 11936 6193 12000
rect 6257 11936 6263 12000
rect 5947 11935 6263 11936
rect 9649 12000 9965 12001
rect 9649 11936 9655 12000
rect 9719 11936 9735 12000
rect 9799 11936 9815 12000
rect 9879 11936 9895 12000
rect 9959 11936 9965 12000
rect 9649 11935 9965 11936
rect 13351 12000 13667 12001
rect 13351 11936 13357 12000
rect 13421 11936 13437 12000
rect 13501 11936 13517 12000
rect 13581 11936 13597 12000
rect 13661 11936 13667 12000
rect 13351 11935 13667 11936
rect 4096 11456 4412 11457
rect 4096 11392 4102 11456
rect 4166 11392 4182 11456
rect 4246 11392 4262 11456
rect 4326 11392 4342 11456
rect 4406 11392 4412 11456
rect 4096 11391 4412 11392
rect 7798 11456 8114 11457
rect 7798 11392 7804 11456
rect 7868 11392 7884 11456
rect 7948 11392 7964 11456
rect 8028 11392 8044 11456
rect 8108 11392 8114 11456
rect 7798 11391 8114 11392
rect 11500 11456 11816 11457
rect 11500 11392 11506 11456
rect 11570 11392 11586 11456
rect 11650 11392 11666 11456
rect 11730 11392 11746 11456
rect 11810 11392 11816 11456
rect 11500 11391 11816 11392
rect 15202 11456 15518 11457
rect 15202 11392 15208 11456
rect 15272 11392 15288 11456
rect 15352 11392 15368 11456
rect 15432 11392 15448 11456
rect 15512 11392 15518 11456
rect 15202 11391 15518 11392
rect 2245 10912 2561 10913
rect 2245 10848 2251 10912
rect 2315 10848 2331 10912
rect 2395 10848 2411 10912
rect 2475 10848 2491 10912
rect 2555 10848 2561 10912
rect 2245 10847 2561 10848
rect 5947 10912 6263 10913
rect 5947 10848 5953 10912
rect 6017 10848 6033 10912
rect 6097 10848 6113 10912
rect 6177 10848 6193 10912
rect 6257 10848 6263 10912
rect 5947 10847 6263 10848
rect 9649 10912 9965 10913
rect 9649 10848 9655 10912
rect 9719 10848 9735 10912
rect 9799 10848 9815 10912
rect 9879 10848 9895 10912
rect 9959 10848 9965 10912
rect 9649 10847 9965 10848
rect 13351 10912 13667 10913
rect 13351 10848 13357 10912
rect 13421 10848 13437 10912
rect 13501 10848 13517 10912
rect 13581 10848 13597 10912
rect 13661 10848 13667 10912
rect 13351 10847 13667 10848
rect 15101 10706 15167 10709
rect 15600 10706 16000 10736
rect 15101 10704 16000 10706
rect 15101 10648 15106 10704
rect 15162 10648 16000 10704
rect 15101 10646 16000 10648
rect 15101 10643 15167 10646
rect 15600 10616 16000 10646
rect 4096 10368 4412 10369
rect 4096 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4342 10368
rect 4406 10304 4412 10368
rect 4096 10303 4412 10304
rect 7798 10368 8114 10369
rect 7798 10304 7804 10368
rect 7868 10304 7884 10368
rect 7948 10304 7964 10368
rect 8028 10304 8044 10368
rect 8108 10304 8114 10368
rect 7798 10303 8114 10304
rect 11500 10368 11816 10369
rect 11500 10304 11506 10368
rect 11570 10304 11586 10368
rect 11650 10304 11666 10368
rect 11730 10304 11746 10368
rect 11810 10304 11816 10368
rect 11500 10303 11816 10304
rect 15202 10368 15518 10369
rect 15202 10304 15208 10368
rect 15272 10304 15288 10368
rect 15352 10304 15368 10368
rect 15432 10304 15448 10368
rect 15512 10304 15518 10368
rect 15202 10303 15518 10304
rect 12893 10162 12959 10165
rect 15101 10162 15167 10165
rect 12893 10160 15167 10162
rect 12893 10104 12898 10160
rect 12954 10104 15106 10160
rect 15162 10104 15167 10160
rect 12893 10102 15167 10104
rect 12893 10099 12959 10102
rect 15101 10099 15167 10102
rect 12801 10026 12867 10029
rect 13445 10026 13511 10029
rect 12801 10024 13511 10026
rect 12801 9968 12806 10024
rect 12862 9968 13450 10024
rect 13506 9968 13511 10024
rect 12801 9966 13511 9968
rect 12801 9963 12867 9966
rect 13445 9963 13511 9966
rect 2245 9824 2561 9825
rect 2245 9760 2251 9824
rect 2315 9760 2331 9824
rect 2395 9760 2411 9824
rect 2475 9760 2491 9824
rect 2555 9760 2561 9824
rect 2245 9759 2561 9760
rect 5947 9824 6263 9825
rect 5947 9760 5953 9824
rect 6017 9760 6033 9824
rect 6097 9760 6113 9824
rect 6177 9760 6193 9824
rect 6257 9760 6263 9824
rect 5947 9759 6263 9760
rect 9649 9824 9965 9825
rect 9649 9760 9655 9824
rect 9719 9760 9735 9824
rect 9799 9760 9815 9824
rect 9879 9760 9895 9824
rect 9959 9760 9965 9824
rect 9649 9759 9965 9760
rect 13351 9824 13667 9825
rect 13351 9760 13357 9824
rect 13421 9760 13437 9824
rect 13501 9760 13517 9824
rect 13581 9760 13597 9824
rect 13661 9760 13667 9824
rect 13351 9759 13667 9760
rect 11237 9482 11303 9485
rect 13169 9482 13235 9485
rect 11237 9480 13235 9482
rect 11237 9424 11242 9480
rect 11298 9424 13174 9480
rect 13230 9424 13235 9480
rect 11237 9422 13235 9424
rect 11237 9419 11303 9422
rect 13169 9419 13235 9422
rect 4096 9280 4412 9281
rect 4096 9216 4102 9280
rect 4166 9216 4182 9280
rect 4246 9216 4262 9280
rect 4326 9216 4342 9280
rect 4406 9216 4412 9280
rect 4096 9215 4412 9216
rect 7798 9280 8114 9281
rect 7798 9216 7804 9280
rect 7868 9216 7884 9280
rect 7948 9216 7964 9280
rect 8028 9216 8044 9280
rect 8108 9216 8114 9280
rect 7798 9215 8114 9216
rect 11500 9280 11816 9281
rect 11500 9216 11506 9280
rect 11570 9216 11586 9280
rect 11650 9216 11666 9280
rect 11730 9216 11746 9280
rect 11810 9216 11816 9280
rect 11500 9215 11816 9216
rect 15202 9280 15518 9281
rect 15202 9216 15208 9280
rect 15272 9216 15288 9280
rect 15352 9216 15368 9280
rect 15432 9216 15448 9280
rect 15512 9216 15518 9280
rect 15202 9215 15518 9216
rect 15101 8802 15167 8805
rect 15600 8802 16000 8832
rect 15101 8800 16000 8802
rect 15101 8744 15106 8800
rect 15162 8744 16000 8800
rect 15101 8742 16000 8744
rect 15101 8739 15167 8742
rect 2245 8736 2561 8737
rect 2245 8672 2251 8736
rect 2315 8672 2331 8736
rect 2395 8672 2411 8736
rect 2475 8672 2491 8736
rect 2555 8672 2561 8736
rect 2245 8671 2561 8672
rect 5947 8736 6263 8737
rect 5947 8672 5953 8736
rect 6017 8672 6033 8736
rect 6097 8672 6113 8736
rect 6177 8672 6193 8736
rect 6257 8672 6263 8736
rect 5947 8671 6263 8672
rect 9649 8736 9965 8737
rect 9649 8672 9655 8736
rect 9719 8672 9735 8736
rect 9799 8672 9815 8736
rect 9879 8672 9895 8736
rect 9959 8672 9965 8736
rect 9649 8671 9965 8672
rect 13351 8736 13667 8737
rect 13351 8672 13357 8736
rect 13421 8672 13437 8736
rect 13501 8672 13517 8736
rect 13581 8672 13597 8736
rect 13661 8672 13667 8736
rect 15600 8712 16000 8742
rect 13351 8671 13667 8672
rect 4096 8192 4412 8193
rect 4096 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4342 8192
rect 4406 8128 4412 8192
rect 4096 8127 4412 8128
rect 7798 8192 8114 8193
rect 7798 8128 7804 8192
rect 7868 8128 7884 8192
rect 7948 8128 7964 8192
rect 8028 8128 8044 8192
rect 8108 8128 8114 8192
rect 7798 8127 8114 8128
rect 11500 8192 11816 8193
rect 11500 8128 11506 8192
rect 11570 8128 11586 8192
rect 11650 8128 11666 8192
rect 11730 8128 11746 8192
rect 11810 8128 11816 8192
rect 11500 8127 11816 8128
rect 15202 8192 15518 8193
rect 15202 8128 15208 8192
rect 15272 8128 15288 8192
rect 15352 8128 15368 8192
rect 15432 8128 15448 8192
rect 15512 8128 15518 8192
rect 15202 8127 15518 8128
rect 2245 7648 2561 7649
rect 2245 7584 2251 7648
rect 2315 7584 2331 7648
rect 2395 7584 2411 7648
rect 2475 7584 2491 7648
rect 2555 7584 2561 7648
rect 2245 7583 2561 7584
rect 5947 7648 6263 7649
rect 5947 7584 5953 7648
rect 6017 7584 6033 7648
rect 6097 7584 6113 7648
rect 6177 7584 6193 7648
rect 6257 7584 6263 7648
rect 5947 7583 6263 7584
rect 9649 7648 9965 7649
rect 9649 7584 9655 7648
rect 9719 7584 9735 7648
rect 9799 7584 9815 7648
rect 9879 7584 9895 7648
rect 9959 7584 9965 7648
rect 9649 7583 9965 7584
rect 13351 7648 13667 7649
rect 13351 7584 13357 7648
rect 13421 7584 13437 7648
rect 13501 7584 13517 7648
rect 13581 7584 13597 7648
rect 13661 7584 13667 7648
rect 13351 7583 13667 7584
rect 4096 7104 4412 7105
rect 4096 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4342 7104
rect 4406 7040 4412 7104
rect 4096 7039 4412 7040
rect 7798 7104 8114 7105
rect 7798 7040 7804 7104
rect 7868 7040 7884 7104
rect 7948 7040 7964 7104
rect 8028 7040 8044 7104
rect 8108 7040 8114 7104
rect 7798 7039 8114 7040
rect 11500 7104 11816 7105
rect 11500 7040 11506 7104
rect 11570 7040 11586 7104
rect 11650 7040 11666 7104
rect 11730 7040 11746 7104
rect 11810 7040 11816 7104
rect 11500 7039 11816 7040
rect 15202 7104 15518 7105
rect 15202 7040 15208 7104
rect 15272 7040 15288 7104
rect 15352 7040 15368 7104
rect 15432 7040 15448 7104
rect 15512 7040 15518 7104
rect 15202 7039 15518 7040
rect 15009 6898 15075 6901
rect 15600 6898 16000 6928
rect 15009 6896 16000 6898
rect 15009 6840 15014 6896
rect 15070 6840 16000 6896
rect 15009 6838 16000 6840
rect 15009 6835 15075 6838
rect 15600 6808 16000 6838
rect 2245 6560 2561 6561
rect 2245 6496 2251 6560
rect 2315 6496 2331 6560
rect 2395 6496 2411 6560
rect 2475 6496 2491 6560
rect 2555 6496 2561 6560
rect 2245 6495 2561 6496
rect 5947 6560 6263 6561
rect 5947 6496 5953 6560
rect 6017 6496 6033 6560
rect 6097 6496 6113 6560
rect 6177 6496 6193 6560
rect 6257 6496 6263 6560
rect 5947 6495 6263 6496
rect 9649 6560 9965 6561
rect 9649 6496 9655 6560
rect 9719 6496 9735 6560
rect 9799 6496 9815 6560
rect 9879 6496 9895 6560
rect 9959 6496 9965 6560
rect 9649 6495 9965 6496
rect 13351 6560 13667 6561
rect 13351 6496 13357 6560
rect 13421 6496 13437 6560
rect 13501 6496 13517 6560
rect 13581 6496 13597 6560
rect 13661 6496 13667 6560
rect 13351 6495 13667 6496
rect 7465 6218 7531 6221
rect 7741 6218 7807 6221
rect 7465 6216 7807 6218
rect 7465 6160 7470 6216
rect 7526 6160 7746 6216
rect 7802 6160 7807 6216
rect 7465 6158 7807 6160
rect 7465 6155 7531 6158
rect 7741 6155 7807 6158
rect 4096 6016 4412 6017
rect 4096 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4342 6016
rect 4406 5952 4412 6016
rect 4096 5951 4412 5952
rect 7798 6016 8114 6017
rect 7798 5952 7804 6016
rect 7868 5952 7884 6016
rect 7948 5952 7964 6016
rect 8028 5952 8044 6016
rect 8108 5952 8114 6016
rect 7798 5951 8114 5952
rect 11500 6016 11816 6017
rect 11500 5952 11506 6016
rect 11570 5952 11586 6016
rect 11650 5952 11666 6016
rect 11730 5952 11746 6016
rect 11810 5952 11816 6016
rect 11500 5951 11816 5952
rect 15202 6016 15518 6017
rect 15202 5952 15208 6016
rect 15272 5952 15288 6016
rect 15352 5952 15368 6016
rect 15432 5952 15448 6016
rect 15512 5952 15518 6016
rect 15202 5951 15518 5952
rect 15101 5538 15167 5541
rect 15101 5536 15762 5538
rect 15101 5480 15106 5536
rect 15162 5480 15762 5536
rect 15101 5478 15762 5480
rect 15101 5475 15167 5478
rect 2245 5472 2561 5473
rect 2245 5408 2251 5472
rect 2315 5408 2331 5472
rect 2395 5408 2411 5472
rect 2475 5408 2491 5472
rect 2555 5408 2561 5472
rect 2245 5407 2561 5408
rect 5947 5472 6263 5473
rect 5947 5408 5953 5472
rect 6017 5408 6033 5472
rect 6097 5408 6113 5472
rect 6177 5408 6193 5472
rect 6257 5408 6263 5472
rect 5947 5407 6263 5408
rect 9649 5472 9965 5473
rect 9649 5408 9655 5472
rect 9719 5408 9735 5472
rect 9799 5408 9815 5472
rect 9879 5408 9895 5472
rect 9959 5408 9965 5472
rect 9649 5407 9965 5408
rect 13351 5472 13667 5473
rect 13351 5408 13357 5472
rect 13421 5408 13437 5472
rect 13501 5408 13517 5472
rect 13581 5408 13597 5472
rect 13661 5408 13667 5472
rect 13351 5407 13667 5408
rect 10869 5130 10935 5133
rect 11881 5130 11947 5133
rect 10869 5128 11947 5130
rect 10869 5072 10874 5128
rect 10930 5072 11886 5128
rect 11942 5072 11947 5128
rect 10869 5070 11947 5072
rect 10869 5067 10935 5070
rect 11881 5067 11947 5070
rect 15702 5024 15762 5478
rect 4096 4928 4412 4929
rect 4096 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4342 4928
rect 4406 4864 4412 4928
rect 4096 4863 4412 4864
rect 7798 4928 8114 4929
rect 7798 4864 7804 4928
rect 7868 4864 7884 4928
rect 7948 4864 7964 4928
rect 8028 4864 8044 4928
rect 8108 4864 8114 4928
rect 7798 4863 8114 4864
rect 11500 4928 11816 4929
rect 11500 4864 11506 4928
rect 11570 4864 11586 4928
rect 11650 4864 11666 4928
rect 11730 4864 11746 4928
rect 11810 4864 11816 4928
rect 11500 4863 11816 4864
rect 15202 4928 15518 4929
rect 15202 4864 15208 4928
rect 15272 4864 15288 4928
rect 15352 4864 15368 4928
rect 15432 4864 15448 4928
rect 15512 4864 15518 4928
rect 15600 4904 16000 5024
rect 15202 4863 15518 4864
rect 10409 4586 10475 4589
rect 11513 4586 11579 4589
rect 10409 4584 11579 4586
rect 10409 4528 10414 4584
rect 10470 4528 11518 4584
rect 11574 4528 11579 4584
rect 10409 4526 11579 4528
rect 10409 4523 10475 4526
rect 11513 4523 11579 4526
rect 2245 4384 2561 4385
rect 2245 4320 2251 4384
rect 2315 4320 2331 4384
rect 2395 4320 2411 4384
rect 2475 4320 2491 4384
rect 2555 4320 2561 4384
rect 2245 4319 2561 4320
rect 5947 4384 6263 4385
rect 5947 4320 5953 4384
rect 6017 4320 6033 4384
rect 6097 4320 6113 4384
rect 6177 4320 6193 4384
rect 6257 4320 6263 4384
rect 5947 4319 6263 4320
rect 9649 4384 9965 4385
rect 9649 4320 9655 4384
rect 9719 4320 9735 4384
rect 9799 4320 9815 4384
rect 9879 4320 9895 4384
rect 9959 4320 9965 4384
rect 9649 4319 9965 4320
rect 13351 4384 13667 4385
rect 13351 4320 13357 4384
rect 13421 4320 13437 4384
rect 13501 4320 13517 4384
rect 13581 4320 13597 4384
rect 13661 4320 13667 4384
rect 13351 4319 13667 4320
rect 4096 3840 4412 3841
rect 4096 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4342 3840
rect 4406 3776 4412 3840
rect 4096 3775 4412 3776
rect 7798 3840 8114 3841
rect 7798 3776 7804 3840
rect 7868 3776 7884 3840
rect 7948 3776 7964 3840
rect 8028 3776 8044 3840
rect 8108 3776 8114 3840
rect 7798 3775 8114 3776
rect 11500 3840 11816 3841
rect 11500 3776 11506 3840
rect 11570 3776 11586 3840
rect 11650 3776 11666 3840
rect 11730 3776 11746 3840
rect 11810 3776 11816 3840
rect 11500 3775 11816 3776
rect 15202 3840 15518 3841
rect 15202 3776 15208 3840
rect 15272 3776 15288 3840
rect 15352 3776 15368 3840
rect 15432 3776 15448 3840
rect 15512 3776 15518 3840
rect 15202 3775 15518 3776
rect 2245 3296 2561 3297
rect 2245 3232 2251 3296
rect 2315 3232 2331 3296
rect 2395 3232 2411 3296
rect 2475 3232 2491 3296
rect 2555 3232 2561 3296
rect 2245 3231 2561 3232
rect 5947 3296 6263 3297
rect 5947 3232 5953 3296
rect 6017 3232 6033 3296
rect 6097 3232 6113 3296
rect 6177 3232 6193 3296
rect 6257 3232 6263 3296
rect 5947 3231 6263 3232
rect 9649 3296 9965 3297
rect 9649 3232 9655 3296
rect 9719 3232 9735 3296
rect 9799 3232 9815 3296
rect 9879 3232 9895 3296
rect 9959 3232 9965 3296
rect 9649 3231 9965 3232
rect 13351 3296 13667 3297
rect 13351 3232 13357 3296
rect 13421 3232 13437 3296
rect 13501 3232 13517 3296
rect 13581 3232 13597 3296
rect 13661 3232 13667 3296
rect 13351 3231 13667 3232
rect 14457 3090 14523 3093
rect 15600 3090 16000 3120
rect 14457 3088 16000 3090
rect 14457 3032 14462 3088
rect 14518 3032 16000 3088
rect 14457 3030 16000 3032
rect 14457 3027 14523 3030
rect 15600 3000 16000 3030
rect 4096 2752 4412 2753
rect 4096 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4342 2752
rect 4406 2688 4412 2752
rect 4096 2687 4412 2688
rect 7798 2752 8114 2753
rect 7798 2688 7804 2752
rect 7868 2688 7884 2752
rect 7948 2688 7964 2752
rect 8028 2688 8044 2752
rect 8108 2688 8114 2752
rect 7798 2687 8114 2688
rect 11500 2752 11816 2753
rect 11500 2688 11506 2752
rect 11570 2688 11586 2752
rect 11650 2688 11666 2752
rect 11730 2688 11746 2752
rect 11810 2688 11816 2752
rect 11500 2687 11816 2688
rect 15202 2752 15518 2753
rect 15202 2688 15208 2752
rect 15272 2688 15288 2752
rect 15352 2688 15368 2752
rect 15432 2688 15448 2752
rect 15512 2688 15518 2752
rect 15202 2687 15518 2688
rect 2245 2208 2561 2209
rect 2245 2144 2251 2208
rect 2315 2144 2331 2208
rect 2395 2144 2411 2208
rect 2475 2144 2491 2208
rect 2555 2144 2561 2208
rect 2245 2143 2561 2144
rect 5947 2208 6263 2209
rect 5947 2144 5953 2208
rect 6017 2144 6033 2208
rect 6097 2144 6113 2208
rect 6177 2144 6193 2208
rect 6257 2144 6263 2208
rect 5947 2143 6263 2144
rect 9649 2208 9965 2209
rect 9649 2144 9655 2208
rect 9719 2144 9735 2208
rect 9799 2144 9815 2208
rect 9879 2144 9895 2208
rect 9959 2144 9965 2208
rect 9649 2143 9965 2144
rect 13351 2208 13667 2209
rect 13351 2144 13357 2208
rect 13421 2144 13437 2208
rect 13501 2144 13517 2208
rect 13581 2144 13597 2208
rect 13661 2144 13667 2208
rect 13351 2143 13667 2144
rect 4096 1664 4412 1665
rect 4096 1600 4102 1664
rect 4166 1600 4182 1664
rect 4246 1600 4262 1664
rect 4326 1600 4342 1664
rect 4406 1600 4412 1664
rect 4096 1599 4412 1600
rect 7798 1664 8114 1665
rect 7798 1600 7804 1664
rect 7868 1600 7884 1664
rect 7948 1600 7964 1664
rect 8028 1600 8044 1664
rect 8108 1600 8114 1664
rect 7798 1599 8114 1600
rect 11500 1664 11816 1665
rect 11500 1600 11506 1664
rect 11570 1600 11586 1664
rect 11650 1600 11666 1664
rect 11730 1600 11746 1664
rect 11810 1600 11816 1664
rect 11500 1599 11816 1600
rect 15202 1664 15518 1665
rect 15202 1600 15208 1664
rect 15272 1600 15288 1664
rect 15352 1600 15368 1664
rect 15432 1600 15448 1664
rect 15512 1600 15518 1664
rect 15202 1599 15518 1600
rect 15009 1186 15075 1189
rect 15600 1186 16000 1216
rect 15009 1184 16000 1186
rect 15009 1128 15014 1184
rect 15070 1128 16000 1184
rect 15009 1126 16000 1128
rect 15009 1123 15075 1126
rect 2245 1120 2561 1121
rect 2245 1056 2251 1120
rect 2315 1056 2331 1120
rect 2395 1056 2411 1120
rect 2475 1056 2491 1120
rect 2555 1056 2561 1120
rect 2245 1055 2561 1056
rect 5947 1120 6263 1121
rect 5947 1056 5953 1120
rect 6017 1056 6033 1120
rect 6097 1056 6113 1120
rect 6177 1056 6193 1120
rect 6257 1056 6263 1120
rect 5947 1055 6263 1056
rect 9649 1120 9965 1121
rect 9649 1056 9655 1120
rect 9719 1056 9735 1120
rect 9799 1056 9815 1120
rect 9879 1056 9895 1120
rect 9959 1056 9965 1120
rect 9649 1055 9965 1056
rect 13351 1120 13667 1121
rect 13351 1056 13357 1120
rect 13421 1056 13437 1120
rect 13501 1056 13517 1120
rect 13581 1056 13597 1120
rect 13661 1056 13667 1120
rect 15600 1096 16000 1126
rect 13351 1055 13667 1056
rect 4096 576 4412 577
rect 4096 512 4102 576
rect 4166 512 4182 576
rect 4246 512 4262 576
rect 4326 512 4342 576
rect 4406 512 4412 576
rect 4096 511 4412 512
rect 7798 576 8114 577
rect 7798 512 7804 576
rect 7868 512 7884 576
rect 7948 512 7964 576
rect 8028 512 8044 576
rect 8108 512 8114 576
rect 7798 511 8114 512
rect 11500 576 11816 577
rect 11500 512 11506 576
rect 11570 512 11586 576
rect 11650 512 11666 576
rect 11730 512 11746 576
rect 11810 512 11816 576
rect 11500 511 11816 512
rect 15202 576 15518 577
rect 15202 512 15208 576
rect 15272 512 15288 576
rect 15352 512 15368 576
rect 15432 512 15448 576
rect 15512 512 15518 576
rect 15202 511 15518 512
<< via3 >>
rect 2251 15260 2315 15264
rect 2251 15204 2255 15260
rect 2255 15204 2311 15260
rect 2311 15204 2315 15260
rect 2251 15200 2315 15204
rect 2331 15260 2395 15264
rect 2331 15204 2335 15260
rect 2335 15204 2391 15260
rect 2391 15204 2395 15260
rect 2331 15200 2395 15204
rect 2411 15260 2475 15264
rect 2411 15204 2415 15260
rect 2415 15204 2471 15260
rect 2471 15204 2475 15260
rect 2411 15200 2475 15204
rect 2491 15260 2555 15264
rect 2491 15204 2495 15260
rect 2495 15204 2551 15260
rect 2551 15204 2555 15260
rect 2491 15200 2555 15204
rect 5953 15260 6017 15264
rect 5953 15204 5957 15260
rect 5957 15204 6013 15260
rect 6013 15204 6017 15260
rect 5953 15200 6017 15204
rect 6033 15260 6097 15264
rect 6033 15204 6037 15260
rect 6037 15204 6093 15260
rect 6093 15204 6097 15260
rect 6033 15200 6097 15204
rect 6113 15260 6177 15264
rect 6113 15204 6117 15260
rect 6117 15204 6173 15260
rect 6173 15204 6177 15260
rect 6113 15200 6177 15204
rect 6193 15260 6257 15264
rect 6193 15204 6197 15260
rect 6197 15204 6253 15260
rect 6253 15204 6257 15260
rect 6193 15200 6257 15204
rect 9655 15260 9719 15264
rect 9655 15204 9659 15260
rect 9659 15204 9715 15260
rect 9715 15204 9719 15260
rect 9655 15200 9719 15204
rect 9735 15260 9799 15264
rect 9735 15204 9739 15260
rect 9739 15204 9795 15260
rect 9795 15204 9799 15260
rect 9735 15200 9799 15204
rect 9815 15260 9879 15264
rect 9815 15204 9819 15260
rect 9819 15204 9875 15260
rect 9875 15204 9879 15260
rect 9815 15200 9879 15204
rect 9895 15260 9959 15264
rect 9895 15204 9899 15260
rect 9899 15204 9955 15260
rect 9955 15204 9959 15260
rect 9895 15200 9959 15204
rect 13357 15260 13421 15264
rect 13357 15204 13361 15260
rect 13361 15204 13417 15260
rect 13417 15204 13421 15260
rect 13357 15200 13421 15204
rect 13437 15260 13501 15264
rect 13437 15204 13441 15260
rect 13441 15204 13497 15260
rect 13497 15204 13501 15260
rect 13437 15200 13501 15204
rect 13517 15260 13581 15264
rect 13517 15204 13521 15260
rect 13521 15204 13577 15260
rect 13577 15204 13581 15260
rect 13517 15200 13581 15204
rect 13597 15260 13661 15264
rect 13597 15204 13601 15260
rect 13601 15204 13657 15260
rect 13657 15204 13661 15260
rect 13597 15200 13661 15204
rect 4102 14716 4166 14720
rect 4102 14660 4106 14716
rect 4106 14660 4162 14716
rect 4162 14660 4166 14716
rect 4102 14656 4166 14660
rect 4182 14716 4246 14720
rect 4182 14660 4186 14716
rect 4186 14660 4242 14716
rect 4242 14660 4246 14716
rect 4182 14656 4246 14660
rect 4262 14716 4326 14720
rect 4262 14660 4266 14716
rect 4266 14660 4322 14716
rect 4322 14660 4326 14716
rect 4262 14656 4326 14660
rect 4342 14716 4406 14720
rect 4342 14660 4346 14716
rect 4346 14660 4402 14716
rect 4402 14660 4406 14716
rect 4342 14656 4406 14660
rect 7804 14716 7868 14720
rect 7804 14660 7808 14716
rect 7808 14660 7864 14716
rect 7864 14660 7868 14716
rect 7804 14656 7868 14660
rect 7884 14716 7948 14720
rect 7884 14660 7888 14716
rect 7888 14660 7944 14716
rect 7944 14660 7948 14716
rect 7884 14656 7948 14660
rect 7964 14716 8028 14720
rect 7964 14660 7968 14716
rect 7968 14660 8024 14716
rect 8024 14660 8028 14716
rect 7964 14656 8028 14660
rect 8044 14716 8108 14720
rect 8044 14660 8048 14716
rect 8048 14660 8104 14716
rect 8104 14660 8108 14716
rect 8044 14656 8108 14660
rect 11506 14716 11570 14720
rect 11506 14660 11510 14716
rect 11510 14660 11566 14716
rect 11566 14660 11570 14716
rect 11506 14656 11570 14660
rect 11586 14716 11650 14720
rect 11586 14660 11590 14716
rect 11590 14660 11646 14716
rect 11646 14660 11650 14716
rect 11586 14656 11650 14660
rect 11666 14716 11730 14720
rect 11666 14660 11670 14716
rect 11670 14660 11726 14716
rect 11726 14660 11730 14716
rect 11666 14656 11730 14660
rect 11746 14716 11810 14720
rect 11746 14660 11750 14716
rect 11750 14660 11806 14716
rect 11806 14660 11810 14716
rect 11746 14656 11810 14660
rect 15208 14716 15272 14720
rect 15208 14660 15212 14716
rect 15212 14660 15268 14716
rect 15268 14660 15272 14716
rect 15208 14656 15272 14660
rect 15288 14716 15352 14720
rect 15288 14660 15292 14716
rect 15292 14660 15348 14716
rect 15348 14660 15352 14716
rect 15288 14656 15352 14660
rect 15368 14716 15432 14720
rect 15368 14660 15372 14716
rect 15372 14660 15428 14716
rect 15428 14660 15432 14716
rect 15368 14656 15432 14660
rect 15448 14716 15512 14720
rect 15448 14660 15452 14716
rect 15452 14660 15508 14716
rect 15508 14660 15512 14716
rect 15448 14656 15512 14660
rect 2251 14172 2315 14176
rect 2251 14116 2255 14172
rect 2255 14116 2311 14172
rect 2311 14116 2315 14172
rect 2251 14112 2315 14116
rect 2331 14172 2395 14176
rect 2331 14116 2335 14172
rect 2335 14116 2391 14172
rect 2391 14116 2395 14172
rect 2331 14112 2395 14116
rect 2411 14172 2475 14176
rect 2411 14116 2415 14172
rect 2415 14116 2471 14172
rect 2471 14116 2475 14172
rect 2411 14112 2475 14116
rect 2491 14172 2555 14176
rect 2491 14116 2495 14172
rect 2495 14116 2551 14172
rect 2551 14116 2555 14172
rect 2491 14112 2555 14116
rect 5953 14172 6017 14176
rect 5953 14116 5957 14172
rect 5957 14116 6013 14172
rect 6013 14116 6017 14172
rect 5953 14112 6017 14116
rect 6033 14172 6097 14176
rect 6033 14116 6037 14172
rect 6037 14116 6093 14172
rect 6093 14116 6097 14172
rect 6033 14112 6097 14116
rect 6113 14172 6177 14176
rect 6113 14116 6117 14172
rect 6117 14116 6173 14172
rect 6173 14116 6177 14172
rect 6113 14112 6177 14116
rect 6193 14172 6257 14176
rect 6193 14116 6197 14172
rect 6197 14116 6253 14172
rect 6253 14116 6257 14172
rect 6193 14112 6257 14116
rect 9655 14172 9719 14176
rect 9655 14116 9659 14172
rect 9659 14116 9715 14172
rect 9715 14116 9719 14172
rect 9655 14112 9719 14116
rect 9735 14172 9799 14176
rect 9735 14116 9739 14172
rect 9739 14116 9795 14172
rect 9795 14116 9799 14172
rect 9735 14112 9799 14116
rect 9815 14172 9879 14176
rect 9815 14116 9819 14172
rect 9819 14116 9875 14172
rect 9875 14116 9879 14172
rect 9815 14112 9879 14116
rect 9895 14172 9959 14176
rect 9895 14116 9899 14172
rect 9899 14116 9955 14172
rect 9955 14116 9959 14172
rect 9895 14112 9959 14116
rect 13357 14172 13421 14176
rect 13357 14116 13361 14172
rect 13361 14116 13417 14172
rect 13417 14116 13421 14172
rect 13357 14112 13421 14116
rect 13437 14172 13501 14176
rect 13437 14116 13441 14172
rect 13441 14116 13497 14172
rect 13497 14116 13501 14172
rect 13437 14112 13501 14116
rect 13517 14172 13581 14176
rect 13517 14116 13521 14172
rect 13521 14116 13577 14172
rect 13577 14116 13581 14172
rect 13517 14112 13581 14116
rect 13597 14172 13661 14176
rect 13597 14116 13601 14172
rect 13601 14116 13657 14172
rect 13657 14116 13661 14172
rect 13597 14112 13661 14116
rect 4102 13628 4166 13632
rect 4102 13572 4106 13628
rect 4106 13572 4162 13628
rect 4162 13572 4166 13628
rect 4102 13568 4166 13572
rect 4182 13628 4246 13632
rect 4182 13572 4186 13628
rect 4186 13572 4242 13628
rect 4242 13572 4246 13628
rect 4182 13568 4246 13572
rect 4262 13628 4326 13632
rect 4262 13572 4266 13628
rect 4266 13572 4322 13628
rect 4322 13572 4326 13628
rect 4262 13568 4326 13572
rect 4342 13628 4406 13632
rect 4342 13572 4346 13628
rect 4346 13572 4402 13628
rect 4402 13572 4406 13628
rect 4342 13568 4406 13572
rect 7804 13628 7868 13632
rect 7804 13572 7808 13628
rect 7808 13572 7864 13628
rect 7864 13572 7868 13628
rect 7804 13568 7868 13572
rect 7884 13628 7948 13632
rect 7884 13572 7888 13628
rect 7888 13572 7944 13628
rect 7944 13572 7948 13628
rect 7884 13568 7948 13572
rect 7964 13628 8028 13632
rect 7964 13572 7968 13628
rect 7968 13572 8024 13628
rect 8024 13572 8028 13628
rect 7964 13568 8028 13572
rect 8044 13628 8108 13632
rect 8044 13572 8048 13628
rect 8048 13572 8104 13628
rect 8104 13572 8108 13628
rect 8044 13568 8108 13572
rect 11506 13628 11570 13632
rect 11506 13572 11510 13628
rect 11510 13572 11566 13628
rect 11566 13572 11570 13628
rect 11506 13568 11570 13572
rect 11586 13628 11650 13632
rect 11586 13572 11590 13628
rect 11590 13572 11646 13628
rect 11646 13572 11650 13628
rect 11586 13568 11650 13572
rect 11666 13628 11730 13632
rect 11666 13572 11670 13628
rect 11670 13572 11726 13628
rect 11726 13572 11730 13628
rect 11666 13568 11730 13572
rect 11746 13628 11810 13632
rect 11746 13572 11750 13628
rect 11750 13572 11806 13628
rect 11806 13572 11810 13628
rect 11746 13568 11810 13572
rect 15208 13628 15272 13632
rect 15208 13572 15212 13628
rect 15212 13572 15268 13628
rect 15268 13572 15272 13628
rect 15208 13568 15272 13572
rect 15288 13628 15352 13632
rect 15288 13572 15292 13628
rect 15292 13572 15348 13628
rect 15348 13572 15352 13628
rect 15288 13568 15352 13572
rect 15368 13628 15432 13632
rect 15368 13572 15372 13628
rect 15372 13572 15428 13628
rect 15428 13572 15432 13628
rect 15368 13568 15432 13572
rect 15448 13628 15512 13632
rect 15448 13572 15452 13628
rect 15452 13572 15508 13628
rect 15508 13572 15512 13628
rect 15448 13568 15512 13572
rect 2251 13084 2315 13088
rect 2251 13028 2255 13084
rect 2255 13028 2311 13084
rect 2311 13028 2315 13084
rect 2251 13024 2315 13028
rect 2331 13084 2395 13088
rect 2331 13028 2335 13084
rect 2335 13028 2391 13084
rect 2391 13028 2395 13084
rect 2331 13024 2395 13028
rect 2411 13084 2475 13088
rect 2411 13028 2415 13084
rect 2415 13028 2471 13084
rect 2471 13028 2475 13084
rect 2411 13024 2475 13028
rect 2491 13084 2555 13088
rect 2491 13028 2495 13084
rect 2495 13028 2551 13084
rect 2551 13028 2555 13084
rect 2491 13024 2555 13028
rect 5953 13084 6017 13088
rect 5953 13028 5957 13084
rect 5957 13028 6013 13084
rect 6013 13028 6017 13084
rect 5953 13024 6017 13028
rect 6033 13084 6097 13088
rect 6033 13028 6037 13084
rect 6037 13028 6093 13084
rect 6093 13028 6097 13084
rect 6033 13024 6097 13028
rect 6113 13084 6177 13088
rect 6113 13028 6117 13084
rect 6117 13028 6173 13084
rect 6173 13028 6177 13084
rect 6113 13024 6177 13028
rect 6193 13084 6257 13088
rect 6193 13028 6197 13084
rect 6197 13028 6253 13084
rect 6253 13028 6257 13084
rect 6193 13024 6257 13028
rect 9655 13084 9719 13088
rect 9655 13028 9659 13084
rect 9659 13028 9715 13084
rect 9715 13028 9719 13084
rect 9655 13024 9719 13028
rect 9735 13084 9799 13088
rect 9735 13028 9739 13084
rect 9739 13028 9795 13084
rect 9795 13028 9799 13084
rect 9735 13024 9799 13028
rect 9815 13084 9879 13088
rect 9815 13028 9819 13084
rect 9819 13028 9875 13084
rect 9875 13028 9879 13084
rect 9815 13024 9879 13028
rect 9895 13084 9959 13088
rect 9895 13028 9899 13084
rect 9899 13028 9955 13084
rect 9955 13028 9959 13084
rect 9895 13024 9959 13028
rect 13357 13084 13421 13088
rect 13357 13028 13361 13084
rect 13361 13028 13417 13084
rect 13417 13028 13421 13084
rect 13357 13024 13421 13028
rect 13437 13084 13501 13088
rect 13437 13028 13441 13084
rect 13441 13028 13497 13084
rect 13497 13028 13501 13084
rect 13437 13024 13501 13028
rect 13517 13084 13581 13088
rect 13517 13028 13521 13084
rect 13521 13028 13577 13084
rect 13577 13028 13581 13084
rect 13517 13024 13581 13028
rect 13597 13084 13661 13088
rect 13597 13028 13601 13084
rect 13601 13028 13657 13084
rect 13657 13028 13661 13084
rect 13597 13024 13661 13028
rect 4102 12540 4166 12544
rect 4102 12484 4106 12540
rect 4106 12484 4162 12540
rect 4162 12484 4166 12540
rect 4102 12480 4166 12484
rect 4182 12540 4246 12544
rect 4182 12484 4186 12540
rect 4186 12484 4242 12540
rect 4242 12484 4246 12540
rect 4182 12480 4246 12484
rect 4262 12540 4326 12544
rect 4262 12484 4266 12540
rect 4266 12484 4322 12540
rect 4322 12484 4326 12540
rect 4262 12480 4326 12484
rect 4342 12540 4406 12544
rect 4342 12484 4346 12540
rect 4346 12484 4402 12540
rect 4402 12484 4406 12540
rect 4342 12480 4406 12484
rect 7804 12540 7868 12544
rect 7804 12484 7808 12540
rect 7808 12484 7864 12540
rect 7864 12484 7868 12540
rect 7804 12480 7868 12484
rect 7884 12540 7948 12544
rect 7884 12484 7888 12540
rect 7888 12484 7944 12540
rect 7944 12484 7948 12540
rect 7884 12480 7948 12484
rect 7964 12540 8028 12544
rect 7964 12484 7968 12540
rect 7968 12484 8024 12540
rect 8024 12484 8028 12540
rect 7964 12480 8028 12484
rect 8044 12540 8108 12544
rect 8044 12484 8048 12540
rect 8048 12484 8104 12540
rect 8104 12484 8108 12540
rect 8044 12480 8108 12484
rect 11506 12540 11570 12544
rect 11506 12484 11510 12540
rect 11510 12484 11566 12540
rect 11566 12484 11570 12540
rect 11506 12480 11570 12484
rect 11586 12540 11650 12544
rect 11586 12484 11590 12540
rect 11590 12484 11646 12540
rect 11646 12484 11650 12540
rect 11586 12480 11650 12484
rect 11666 12540 11730 12544
rect 11666 12484 11670 12540
rect 11670 12484 11726 12540
rect 11726 12484 11730 12540
rect 11666 12480 11730 12484
rect 11746 12540 11810 12544
rect 11746 12484 11750 12540
rect 11750 12484 11806 12540
rect 11806 12484 11810 12540
rect 11746 12480 11810 12484
rect 15208 12540 15272 12544
rect 15208 12484 15212 12540
rect 15212 12484 15268 12540
rect 15268 12484 15272 12540
rect 15208 12480 15272 12484
rect 15288 12540 15352 12544
rect 15288 12484 15292 12540
rect 15292 12484 15348 12540
rect 15348 12484 15352 12540
rect 15288 12480 15352 12484
rect 15368 12540 15432 12544
rect 15368 12484 15372 12540
rect 15372 12484 15428 12540
rect 15428 12484 15432 12540
rect 15368 12480 15432 12484
rect 15448 12540 15512 12544
rect 15448 12484 15452 12540
rect 15452 12484 15508 12540
rect 15508 12484 15512 12540
rect 15448 12480 15512 12484
rect 2251 11996 2315 12000
rect 2251 11940 2255 11996
rect 2255 11940 2311 11996
rect 2311 11940 2315 11996
rect 2251 11936 2315 11940
rect 2331 11996 2395 12000
rect 2331 11940 2335 11996
rect 2335 11940 2391 11996
rect 2391 11940 2395 11996
rect 2331 11936 2395 11940
rect 2411 11996 2475 12000
rect 2411 11940 2415 11996
rect 2415 11940 2471 11996
rect 2471 11940 2475 11996
rect 2411 11936 2475 11940
rect 2491 11996 2555 12000
rect 2491 11940 2495 11996
rect 2495 11940 2551 11996
rect 2551 11940 2555 11996
rect 2491 11936 2555 11940
rect 5953 11996 6017 12000
rect 5953 11940 5957 11996
rect 5957 11940 6013 11996
rect 6013 11940 6017 11996
rect 5953 11936 6017 11940
rect 6033 11996 6097 12000
rect 6033 11940 6037 11996
rect 6037 11940 6093 11996
rect 6093 11940 6097 11996
rect 6033 11936 6097 11940
rect 6113 11996 6177 12000
rect 6113 11940 6117 11996
rect 6117 11940 6173 11996
rect 6173 11940 6177 11996
rect 6113 11936 6177 11940
rect 6193 11996 6257 12000
rect 6193 11940 6197 11996
rect 6197 11940 6253 11996
rect 6253 11940 6257 11996
rect 6193 11936 6257 11940
rect 9655 11996 9719 12000
rect 9655 11940 9659 11996
rect 9659 11940 9715 11996
rect 9715 11940 9719 11996
rect 9655 11936 9719 11940
rect 9735 11996 9799 12000
rect 9735 11940 9739 11996
rect 9739 11940 9795 11996
rect 9795 11940 9799 11996
rect 9735 11936 9799 11940
rect 9815 11996 9879 12000
rect 9815 11940 9819 11996
rect 9819 11940 9875 11996
rect 9875 11940 9879 11996
rect 9815 11936 9879 11940
rect 9895 11996 9959 12000
rect 9895 11940 9899 11996
rect 9899 11940 9955 11996
rect 9955 11940 9959 11996
rect 9895 11936 9959 11940
rect 13357 11996 13421 12000
rect 13357 11940 13361 11996
rect 13361 11940 13417 11996
rect 13417 11940 13421 11996
rect 13357 11936 13421 11940
rect 13437 11996 13501 12000
rect 13437 11940 13441 11996
rect 13441 11940 13497 11996
rect 13497 11940 13501 11996
rect 13437 11936 13501 11940
rect 13517 11996 13581 12000
rect 13517 11940 13521 11996
rect 13521 11940 13577 11996
rect 13577 11940 13581 11996
rect 13517 11936 13581 11940
rect 13597 11996 13661 12000
rect 13597 11940 13601 11996
rect 13601 11940 13657 11996
rect 13657 11940 13661 11996
rect 13597 11936 13661 11940
rect 4102 11452 4166 11456
rect 4102 11396 4106 11452
rect 4106 11396 4162 11452
rect 4162 11396 4166 11452
rect 4102 11392 4166 11396
rect 4182 11452 4246 11456
rect 4182 11396 4186 11452
rect 4186 11396 4242 11452
rect 4242 11396 4246 11452
rect 4182 11392 4246 11396
rect 4262 11452 4326 11456
rect 4262 11396 4266 11452
rect 4266 11396 4322 11452
rect 4322 11396 4326 11452
rect 4262 11392 4326 11396
rect 4342 11452 4406 11456
rect 4342 11396 4346 11452
rect 4346 11396 4402 11452
rect 4402 11396 4406 11452
rect 4342 11392 4406 11396
rect 7804 11452 7868 11456
rect 7804 11396 7808 11452
rect 7808 11396 7864 11452
rect 7864 11396 7868 11452
rect 7804 11392 7868 11396
rect 7884 11452 7948 11456
rect 7884 11396 7888 11452
rect 7888 11396 7944 11452
rect 7944 11396 7948 11452
rect 7884 11392 7948 11396
rect 7964 11452 8028 11456
rect 7964 11396 7968 11452
rect 7968 11396 8024 11452
rect 8024 11396 8028 11452
rect 7964 11392 8028 11396
rect 8044 11452 8108 11456
rect 8044 11396 8048 11452
rect 8048 11396 8104 11452
rect 8104 11396 8108 11452
rect 8044 11392 8108 11396
rect 11506 11452 11570 11456
rect 11506 11396 11510 11452
rect 11510 11396 11566 11452
rect 11566 11396 11570 11452
rect 11506 11392 11570 11396
rect 11586 11452 11650 11456
rect 11586 11396 11590 11452
rect 11590 11396 11646 11452
rect 11646 11396 11650 11452
rect 11586 11392 11650 11396
rect 11666 11452 11730 11456
rect 11666 11396 11670 11452
rect 11670 11396 11726 11452
rect 11726 11396 11730 11452
rect 11666 11392 11730 11396
rect 11746 11452 11810 11456
rect 11746 11396 11750 11452
rect 11750 11396 11806 11452
rect 11806 11396 11810 11452
rect 11746 11392 11810 11396
rect 15208 11452 15272 11456
rect 15208 11396 15212 11452
rect 15212 11396 15268 11452
rect 15268 11396 15272 11452
rect 15208 11392 15272 11396
rect 15288 11452 15352 11456
rect 15288 11396 15292 11452
rect 15292 11396 15348 11452
rect 15348 11396 15352 11452
rect 15288 11392 15352 11396
rect 15368 11452 15432 11456
rect 15368 11396 15372 11452
rect 15372 11396 15428 11452
rect 15428 11396 15432 11452
rect 15368 11392 15432 11396
rect 15448 11452 15512 11456
rect 15448 11396 15452 11452
rect 15452 11396 15508 11452
rect 15508 11396 15512 11452
rect 15448 11392 15512 11396
rect 2251 10908 2315 10912
rect 2251 10852 2255 10908
rect 2255 10852 2311 10908
rect 2311 10852 2315 10908
rect 2251 10848 2315 10852
rect 2331 10908 2395 10912
rect 2331 10852 2335 10908
rect 2335 10852 2391 10908
rect 2391 10852 2395 10908
rect 2331 10848 2395 10852
rect 2411 10908 2475 10912
rect 2411 10852 2415 10908
rect 2415 10852 2471 10908
rect 2471 10852 2475 10908
rect 2411 10848 2475 10852
rect 2491 10908 2555 10912
rect 2491 10852 2495 10908
rect 2495 10852 2551 10908
rect 2551 10852 2555 10908
rect 2491 10848 2555 10852
rect 5953 10908 6017 10912
rect 5953 10852 5957 10908
rect 5957 10852 6013 10908
rect 6013 10852 6017 10908
rect 5953 10848 6017 10852
rect 6033 10908 6097 10912
rect 6033 10852 6037 10908
rect 6037 10852 6093 10908
rect 6093 10852 6097 10908
rect 6033 10848 6097 10852
rect 6113 10908 6177 10912
rect 6113 10852 6117 10908
rect 6117 10852 6173 10908
rect 6173 10852 6177 10908
rect 6113 10848 6177 10852
rect 6193 10908 6257 10912
rect 6193 10852 6197 10908
rect 6197 10852 6253 10908
rect 6253 10852 6257 10908
rect 6193 10848 6257 10852
rect 9655 10908 9719 10912
rect 9655 10852 9659 10908
rect 9659 10852 9715 10908
rect 9715 10852 9719 10908
rect 9655 10848 9719 10852
rect 9735 10908 9799 10912
rect 9735 10852 9739 10908
rect 9739 10852 9795 10908
rect 9795 10852 9799 10908
rect 9735 10848 9799 10852
rect 9815 10908 9879 10912
rect 9815 10852 9819 10908
rect 9819 10852 9875 10908
rect 9875 10852 9879 10908
rect 9815 10848 9879 10852
rect 9895 10908 9959 10912
rect 9895 10852 9899 10908
rect 9899 10852 9955 10908
rect 9955 10852 9959 10908
rect 9895 10848 9959 10852
rect 13357 10908 13421 10912
rect 13357 10852 13361 10908
rect 13361 10852 13417 10908
rect 13417 10852 13421 10908
rect 13357 10848 13421 10852
rect 13437 10908 13501 10912
rect 13437 10852 13441 10908
rect 13441 10852 13497 10908
rect 13497 10852 13501 10908
rect 13437 10848 13501 10852
rect 13517 10908 13581 10912
rect 13517 10852 13521 10908
rect 13521 10852 13577 10908
rect 13577 10852 13581 10908
rect 13517 10848 13581 10852
rect 13597 10908 13661 10912
rect 13597 10852 13601 10908
rect 13601 10852 13657 10908
rect 13657 10852 13661 10908
rect 13597 10848 13661 10852
rect 4102 10364 4166 10368
rect 4102 10308 4106 10364
rect 4106 10308 4162 10364
rect 4162 10308 4166 10364
rect 4102 10304 4166 10308
rect 4182 10364 4246 10368
rect 4182 10308 4186 10364
rect 4186 10308 4242 10364
rect 4242 10308 4246 10364
rect 4182 10304 4246 10308
rect 4262 10364 4326 10368
rect 4262 10308 4266 10364
rect 4266 10308 4322 10364
rect 4322 10308 4326 10364
rect 4262 10304 4326 10308
rect 4342 10364 4406 10368
rect 4342 10308 4346 10364
rect 4346 10308 4402 10364
rect 4402 10308 4406 10364
rect 4342 10304 4406 10308
rect 7804 10364 7868 10368
rect 7804 10308 7808 10364
rect 7808 10308 7864 10364
rect 7864 10308 7868 10364
rect 7804 10304 7868 10308
rect 7884 10364 7948 10368
rect 7884 10308 7888 10364
rect 7888 10308 7944 10364
rect 7944 10308 7948 10364
rect 7884 10304 7948 10308
rect 7964 10364 8028 10368
rect 7964 10308 7968 10364
rect 7968 10308 8024 10364
rect 8024 10308 8028 10364
rect 7964 10304 8028 10308
rect 8044 10364 8108 10368
rect 8044 10308 8048 10364
rect 8048 10308 8104 10364
rect 8104 10308 8108 10364
rect 8044 10304 8108 10308
rect 11506 10364 11570 10368
rect 11506 10308 11510 10364
rect 11510 10308 11566 10364
rect 11566 10308 11570 10364
rect 11506 10304 11570 10308
rect 11586 10364 11650 10368
rect 11586 10308 11590 10364
rect 11590 10308 11646 10364
rect 11646 10308 11650 10364
rect 11586 10304 11650 10308
rect 11666 10364 11730 10368
rect 11666 10308 11670 10364
rect 11670 10308 11726 10364
rect 11726 10308 11730 10364
rect 11666 10304 11730 10308
rect 11746 10364 11810 10368
rect 11746 10308 11750 10364
rect 11750 10308 11806 10364
rect 11806 10308 11810 10364
rect 11746 10304 11810 10308
rect 15208 10364 15272 10368
rect 15208 10308 15212 10364
rect 15212 10308 15268 10364
rect 15268 10308 15272 10364
rect 15208 10304 15272 10308
rect 15288 10364 15352 10368
rect 15288 10308 15292 10364
rect 15292 10308 15348 10364
rect 15348 10308 15352 10364
rect 15288 10304 15352 10308
rect 15368 10364 15432 10368
rect 15368 10308 15372 10364
rect 15372 10308 15428 10364
rect 15428 10308 15432 10364
rect 15368 10304 15432 10308
rect 15448 10364 15512 10368
rect 15448 10308 15452 10364
rect 15452 10308 15508 10364
rect 15508 10308 15512 10364
rect 15448 10304 15512 10308
rect 2251 9820 2315 9824
rect 2251 9764 2255 9820
rect 2255 9764 2311 9820
rect 2311 9764 2315 9820
rect 2251 9760 2315 9764
rect 2331 9820 2395 9824
rect 2331 9764 2335 9820
rect 2335 9764 2391 9820
rect 2391 9764 2395 9820
rect 2331 9760 2395 9764
rect 2411 9820 2475 9824
rect 2411 9764 2415 9820
rect 2415 9764 2471 9820
rect 2471 9764 2475 9820
rect 2411 9760 2475 9764
rect 2491 9820 2555 9824
rect 2491 9764 2495 9820
rect 2495 9764 2551 9820
rect 2551 9764 2555 9820
rect 2491 9760 2555 9764
rect 5953 9820 6017 9824
rect 5953 9764 5957 9820
rect 5957 9764 6013 9820
rect 6013 9764 6017 9820
rect 5953 9760 6017 9764
rect 6033 9820 6097 9824
rect 6033 9764 6037 9820
rect 6037 9764 6093 9820
rect 6093 9764 6097 9820
rect 6033 9760 6097 9764
rect 6113 9820 6177 9824
rect 6113 9764 6117 9820
rect 6117 9764 6173 9820
rect 6173 9764 6177 9820
rect 6113 9760 6177 9764
rect 6193 9820 6257 9824
rect 6193 9764 6197 9820
rect 6197 9764 6253 9820
rect 6253 9764 6257 9820
rect 6193 9760 6257 9764
rect 9655 9820 9719 9824
rect 9655 9764 9659 9820
rect 9659 9764 9715 9820
rect 9715 9764 9719 9820
rect 9655 9760 9719 9764
rect 9735 9820 9799 9824
rect 9735 9764 9739 9820
rect 9739 9764 9795 9820
rect 9795 9764 9799 9820
rect 9735 9760 9799 9764
rect 9815 9820 9879 9824
rect 9815 9764 9819 9820
rect 9819 9764 9875 9820
rect 9875 9764 9879 9820
rect 9815 9760 9879 9764
rect 9895 9820 9959 9824
rect 9895 9764 9899 9820
rect 9899 9764 9955 9820
rect 9955 9764 9959 9820
rect 9895 9760 9959 9764
rect 13357 9820 13421 9824
rect 13357 9764 13361 9820
rect 13361 9764 13417 9820
rect 13417 9764 13421 9820
rect 13357 9760 13421 9764
rect 13437 9820 13501 9824
rect 13437 9764 13441 9820
rect 13441 9764 13497 9820
rect 13497 9764 13501 9820
rect 13437 9760 13501 9764
rect 13517 9820 13581 9824
rect 13517 9764 13521 9820
rect 13521 9764 13577 9820
rect 13577 9764 13581 9820
rect 13517 9760 13581 9764
rect 13597 9820 13661 9824
rect 13597 9764 13601 9820
rect 13601 9764 13657 9820
rect 13657 9764 13661 9820
rect 13597 9760 13661 9764
rect 4102 9276 4166 9280
rect 4102 9220 4106 9276
rect 4106 9220 4162 9276
rect 4162 9220 4166 9276
rect 4102 9216 4166 9220
rect 4182 9276 4246 9280
rect 4182 9220 4186 9276
rect 4186 9220 4242 9276
rect 4242 9220 4246 9276
rect 4182 9216 4246 9220
rect 4262 9276 4326 9280
rect 4262 9220 4266 9276
rect 4266 9220 4322 9276
rect 4322 9220 4326 9276
rect 4262 9216 4326 9220
rect 4342 9276 4406 9280
rect 4342 9220 4346 9276
rect 4346 9220 4402 9276
rect 4402 9220 4406 9276
rect 4342 9216 4406 9220
rect 7804 9276 7868 9280
rect 7804 9220 7808 9276
rect 7808 9220 7864 9276
rect 7864 9220 7868 9276
rect 7804 9216 7868 9220
rect 7884 9276 7948 9280
rect 7884 9220 7888 9276
rect 7888 9220 7944 9276
rect 7944 9220 7948 9276
rect 7884 9216 7948 9220
rect 7964 9276 8028 9280
rect 7964 9220 7968 9276
rect 7968 9220 8024 9276
rect 8024 9220 8028 9276
rect 7964 9216 8028 9220
rect 8044 9276 8108 9280
rect 8044 9220 8048 9276
rect 8048 9220 8104 9276
rect 8104 9220 8108 9276
rect 8044 9216 8108 9220
rect 11506 9276 11570 9280
rect 11506 9220 11510 9276
rect 11510 9220 11566 9276
rect 11566 9220 11570 9276
rect 11506 9216 11570 9220
rect 11586 9276 11650 9280
rect 11586 9220 11590 9276
rect 11590 9220 11646 9276
rect 11646 9220 11650 9276
rect 11586 9216 11650 9220
rect 11666 9276 11730 9280
rect 11666 9220 11670 9276
rect 11670 9220 11726 9276
rect 11726 9220 11730 9276
rect 11666 9216 11730 9220
rect 11746 9276 11810 9280
rect 11746 9220 11750 9276
rect 11750 9220 11806 9276
rect 11806 9220 11810 9276
rect 11746 9216 11810 9220
rect 15208 9276 15272 9280
rect 15208 9220 15212 9276
rect 15212 9220 15268 9276
rect 15268 9220 15272 9276
rect 15208 9216 15272 9220
rect 15288 9276 15352 9280
rect 15288 9220 15292 9276
rect 15292 9220 15348 9276
rect 15348 9220 15352 9276
rect 15288 9216 15352 9220
rect 15368 9276 15432 9280
rect 15368 9220 15372 9276
rect 15372 9220 15428 9276
rect 15428 9220 15432 9276
rect 15368 9216 15432 9220
rect 15448 9276 15512 9280
rect 15448 9220 15452 9276
rect 15452 9220 15508 9276
rect 15508 9220 15512 9276
rect 15448 9216 15512 9220
rect 2251 8732 2315 8736
rect 2251 8676 2255 8732
rect 2255 8676 2311 8732
rect 2311 8676 2315 8732
rect 2251 8672 2315 8676
rect 2331 8732 2395 8736
rect 2331 8676 2335 8732
rect 2335 8676 2391 8732
rect 2391 8676 2395 8732
rect 2331 8672 2395 8676
rect 2411 8732 2475 8736
rect 2411 8676 2415 8732
rect 2415 8676 2471 8732
rect 2471 8676 2475 8732
rect 2411 8672 2475 8676
rect 2491 8732 2555 8736
rect 2491 8676 2495 8732
rect 2495 8676 2551 8732
rect 2551 8676 2555 8732
rect 2491 8672 2555 8676
rect 5953 8732 6017 8736
rect 5953 8676 5957 8732
rect 5957 8676 6013 8732
rect 6013 8676 6017 8732
rect 5953 8672 6017 8676
rect 6033 8732 6097 8736
rect 6033 8676 6037 8732
rect 6037 8676 6093 8732
rect 6093 8676 6097 8732
rect 6033 8672 6097 8676
rect 6113 8732 6177 8736
rect 6113 8676 6117 8732
rect 6117 8676 6173 8732
rect 6173 8676 6177 8732
rect 6113 8672 6177 8676
rect 6193 8732 6257 8736
rect 6193 8676 6197 8732
rect 6197 8676 6253 8732
rect 6253 8676 6257 8732
rect 6193 8672 6257 8676
rect 9655 8732 9719 8736
rect 9655 8676 9659 8732
rect 9659 8676 9715 8732
rect 9715 8676 9719 8732
rect 9655 8672 9719 8676
rect 9735 8732 9799 8736
rect 9735 8676 9739 8732
rect 9739 8676 9795 8732
rect 9795 8676 9799 8732
rect 9735 8672 9799 8676
rect 9815 8732 9879 8736
rect 9815 8676 9819 8732
rect 9819 8676 9875 8732
rect 9875 8676 9879 8732
rect 9815 8672 9879 8676
rect 9895 8732 9959 8736
rect 9895 8676 9899 8732
rect 9899 8676 9955 8732
rect 9955 8676 9959 8732
rect 9895 8672 9959 8676
rect 13357 8732 13421 8736
rect 13357 8676 13361 8732
rect 13361 8676 13417 8732
rect 13417 8676 13421 8732
rect 13357 8672 13421 8676
rect 13437 8732 13501 8736
rect 13437 8676 13441 8732
rect 13441 8676 13497 8732
rect 13497 8676 13501 8732
rect 13437 8672 13501 8676
rect 13517 8732 13581 8736
rect 13517 8676 13521 8732
rect 13521 8676 13577 8732
rect 13577 8676 13581 8732
rect 13517 8672 13581 8676
rect 13597 8732 13661 8736
rect 13597 8676 13601 8732
rect 13601 8676 13657 8732
rect 13657 8676 13661 8732
rect 13597 8672 13661 8676
rect 4102 8188 4166 8192
rect 4102 8132 4106 8188
rect 4106 8132 4162 8188
rect 4162 8132 4166 8188
rect 4102 8128 4166 8132
rect 4182 8188 4246 8192
rect 4182 8132 4186 8188
rect 4186 8132 4242 8188
rect 4242 8132 4246 8188
rect 4182 8128 4246 8132
rect 4262 8188 4326 8192
rect 4262 8132 4266 8188
rect 4266 8132 4322 8188
rect 4322 8132 4326 8188
rect 4262 8128 4326 8132
rect 4342 8188 4406 8192
rect 4342 8132 4346 8188
rect 4346 8132 4402 8188
rect 4402 8132 4406 8188
rect 4342 8128 4406 8132
rect 7804 8188 7868 8192
rect 7804 8132 7808 8188
rect 7808 8132 7864 8188
rect 7864 8132 7868 8188
rect 7804 8128 7868 8132
rect 7884 8188 7948 8192
rect 7884 8132 7888 8188
rect 7888 8132 7944 8188
rect 7944 8132 7948 8188
rect 7884 8128 7948 8132
rect 7964 8188 8028 8192
rect 7964 8132 7968 8188
rect 7968 8132 8024 8188
rect 8024 8132 8028 8188
rect 7964 8128 8028 8132
rect 8044 8188 8108 8192
rect 8044 8132 8048 8188
rect 8048 8132 8104 8188
rect 8104 8132 8108 8188
rect 8044 8128 8108 8132
rect 11506 8188 11570 8192
rect 11506 8132 11510 8188
rect 11510 8132 11566 8188
rect 11566 8132 11570 8188
rect 11506 8128 11570 8132
rect 11586 8188 11650 8192
rect 11586 8132 11590 8188
rect 11590 8132 11646 8188
rect 11646 8132 11650 8188
rect 11586 8128 11650 8132
rect 11666 8188 11730 8192
rect 11666 8132 11670 8188
rect 11670 8132 11726 8188
rect 11726 8132 11730 8188
rect 11666 8128 11730 8132
rect 11746 8188 11810 8192
rect 11746 8132 11750 8188
rect 11750 8132 11806 8188
rect 11806 8132 11810 8188
rect 11746 8128 11810 8132
rect 15208 8188 15272 8192
rect 15208 8132 15212 8188
rect 15212 8132 15268 8188
rect 15268 8132 15272 8188
rect 15208 8128 15272 8132
rect 15288 8188 15352 8192
rect 15288 8132 15292 8188
rect 15292 8132 15348 8188
rect 15348 8132 15352 8188
rect 15288 8128 15352 8132
rect 15368 8188 15432 8192
rect 15368 8132 15372 8188
rect 15372 8132 15428 8188
rect 15428 8132 15432 8188
rect 15368 8128 15432 8132
rect 15448 8188 15512 8192
rect 15448 8132 15452 8188
rect 15452 8132 15508 8188
rect 15508 8132 15512 8188
rect 15448 8128 15512 8132
rect 2251 7644 2315 7648
rect 2251 7588 2255 7644
rect 2255 7588 2311 7644
rect 2311 7588 2315 7644
rect 2251 7584 2315 7588
rect 2331 7644 2395 7648
rect 2331 7588 2335 7644
rect 2335 7588 2391 7644
rect 2391 7588 2395 7644
rect 2331 7584 2395 7588
rect 2411 7644 2475 7648
rect 2411 7588 2415 7644
rect 2415 7588 2471 7644
rect 2471 7588 2475 7644
rect 2411 7584 2475 7588
rect 2491 7644 2555 7648
rect 2491 7588 2495 7644
rect 2495 7588 2551 7644
rect 2551 7588 2555 7644
rect 2491 7584 2555 7588
rect 5953 7644 6017 7648
rect 5953 7588 5957 7644
rect 5957 7588 6013 7644
rect 6013 7588 6017 7644
rect 5953 7584 6017 7588
rect 6033 7644 6097 7648
rect 6033 7588 6037 7644
rect 6037 7588 6093 7644
rect 6093 7588 6097 7644
rect 6033 7584 6097 7588
rect 6113 7644 6177 7648
rect 6113 7588 6117 7644
rect 6117 7588 6173 7644
rect 6173 7588 6177 7644
rect 6113 7584 6177 7588
rect 6193 7644 6257 7648
rect 6193 7588 6197 7644
rect 6197 7588 6253 7644
rect 6253 7588 6257 7644
rect 6193 7584 6257 7588
rect 9655 7644 9719 7648
rect 9655 7588 9659 7644
rect 9659 7588 9715 7644
rect 9715 7588 9719 7644
rect 9655 7584 9719 7588
rect 9735 7644 9799 7648
rect 9735 7588 9739 7644
rect 9739 7588 9795 7644
rect 9795 7588 9799 7644
rect 9735 7584 9799 7588
rect 9815 7644 9879 7648
rect 9815 7588 9819 7644
rect 9819 7588 9875 7644
rect 9875 7588 9879 7644
rect 9815 7584 9879 7588
rect 9895 7644 9959 7648
rect 9895 7588 9899 7644
rect 9899 7588 9955 7644
rect 9955 7588 9959 7644
rect 9895 7584 9959 7588
rect 13357 7644 13421 7648
rect 13357 7588 13361 7644
rect 13361 7588 13417 7644
rect 13417 7588 13421 7644
rect 13357 7584 13421 7588
rect 13437 7644 13501 7648
rect 13437 7588 13441 7644
rect 13441 7588 13497 7644
rect 13497 7588 13501 7644
rect 13437 7584 13501 7588
rect 13517 7644 13581 7648
rect 13517 7588 13521 7644
rect 13521 7588 13577 7644
rect 13577 7588 13581 7644
rect 13517 7584 13581 7588
rect 13597 7644 13661 7648
rect 13597 7588 13601 7644
rect 13601 7588 13657 7644
rect 13657 7588 13661 7644
rect 13597 7584 13661 7588
rect 4102 7100 4166 7104
rect 4102 7044 4106 7100
rect 4106 7044 4162 7100
rect 4162 7044 4166 7100
rect 4102 7040 4166 7044
rect 4182 7100 4246 7104
rect 4182 7044 4186 7100
rect 4186 7044 4242 7100
rect 4242 7044 4246 7100
rect 4182 7040 4246 7044
rect 4262 7100 4326 7104
rect 4262 7044 4266 7100
rect 4266 7044 4322 7100
rect 4322 7044 4326 7100
rect 4262 7040 4326 7044
rect 4342 7100 4406 7104
rect 4342 7044 4346 7100
rect 4346 7044 4402 7100
rect 4402 7044 4406 7100
rect 4342 7040 4406 7044
rect 7804 7100 7868 7104
rect 7804 7044 7808 7100
rect 7808 7044 7864 7100
rect 7864 7044 7868 7100
rect 7804 7040 7868 7044
rect 7884 7100 7948 7104
rect 7884 7044 7888 7100
rect 7888 7044 7944 7100
rect 7944 7044 7948 7100
rect 7884 7040 7948 7044
rect 7964 7100 8028 7104
rect 7964 7044 7968 7100
rect 7968 7044 8024 7100
rect 8024 7044 8028 7100
rect 7964 7040 8028 7044
rect 8044 7100 8108 7104
rect 8044 7044 8048 7100
rect 8048 7044 8104 7100
rect 8104 7044 8108 7100
rect 8044 7040 8108 7044
rect 11506 7100 11570 7104
rect 11506 7044 11510 7100
rect 11510 7044 11566 7100
rect 11566 7044 11570 7100
rect 11506 7040 11570 7044
rect 11586 7100 11650 7104
rect 11586 7044 11590 7100
rect 11590 7044 11646 7100
rect 11646 7044 11650 7100
rect 11586 7040 11650 7044
rect 11666 7100 11730 7104
rect 11666 7044 11670 7100
rect 11670 7044 11726 7100
rect 11726 7044 11730 7100
rect 11666 7040 11730 7044
rect 11746 7100 11810 7104
rect 11746 7044 11750 7100
rect 11750 7044 11806 7100
rect 11806 7044 11810 7100
rect 11746 7040 11810 7044
rect 15208 7100 15272 7104
rect 15208 7044 15212 7100
rect 15212 7044 15268 7100
rect 15268 7044 15272 7100
rect 15208 7040 15272 7044
rect 15288 7100 15352 7104
rect 15288 7044 15292 7100
rect 15292 7044 15348 7100
rect 15348 7044 15352 7100
rect 15288 7040 15352 7044
rect 15368 7100 15432 7104
rect 15368 7044 15372 7100
rect 15372 7044 15428 7100
rect 15428 7044 15432 7100
rect 15368 7040 15432 7044
rect 15448 7100 15512 7104
rect 15448 7044 15452 7100
rect 15452 7044 15508 7100
rect 15508 7044 15512 7100
rect 15448 7040 15512 7044
rect 2251 6556 2315 6560
rect 2251 6500 2255 6556
rect 2255 6500 2311 6556
rect 2311 6500 2315 6556
rect 2251 6496 2315 6500
rect 2331 6556 2395 6560
rect 2331 6500 2335 6556
rect 2335 6500 2391 6556
rect 2391 6500 2395 6556
rect 2331 6496 2395 6500
rect 2411 6556 2475 6560
rect 2411 6500 2415 6556
rect 2415 6500 2471 6556
rect 2471 6500 2475 6556
rect 2411 6496 2475 6500
rect 2491 6556 2555 6560
rect 2491 6500 2495 6556
rect 2495 6500 2551 6556
rect 2551 6500 2555 6556
rect 2491 6496 2555 6500
rect 5953 6556 6017 6560
rect 5953 6500 5957 6556
rect 5957 6500 6013 6556
rect 6013 6500 6017 6556
rect 5953 6496 6017 6500
rect 6033 6556 6097 6560
rect 6033 6500 6037 6556
rect 6037 6500 6093 6556
rect 6093 6500 6097 6556
rect 6033 6496 6097 6500
rect 6113 6556 6177 6560
rect 6113 6500 6117 6556
rect 6117 6500 6173 6556
rect 6173 6500 6177 6556
rect 6113 6496 6177 6500
rect 6193 6556 6257 6560
rect 6193 6500 6197 6556
rect 6197 6500 6253 6556
rect 6253 6500 6257 6556
rect 6193 6496 6257 6500
rect 9655 6556 9719 6560
rect 9655 6500 9659 6556
rect 9659 6500 9715 6556
rect 9715 6500 9719 6556
rect 9655 6496 9719 6500
rect 9735 6556 9799 6560
rect 9735 6500 9739 6556
rect 9739 6500 9795 6556
rect 9795 6500 9799 6556
rect 9735 6496 9799 6500
rect 9815 6556 9879 6560
rect 9815 6500 9819 6556
rect 9819 6500 9875 6556
rect 9875 6500 9879 6556
rect 9815 6496 9879 6500
rect 9895 6556 9959 6560
rect 9895 6500 9899 6556
rect 9899 6500 9955 6556
rect 9955 6500 9959 6556
rect 9895 6496 9959 6500
rect 13357 6556 13421 6560
rect 13357 6500 13361 6556
rect 13361 6500 13417 6556
rect 13417 6500 13421 6556
rect 13357 6496 13421 6500
rect 13437 6556 13501 6560
rect 13437 6500 13441 6556
rect 13441 6500 13497 6556
rect 13497 6500 13501 6556
rect 13437 6496 13501 6500
rect 13517 6556 13581 6560
rect 13517 6500 13521 6556
rect 13521 6500 13577 6556
rect 13577 6500 13581 6556
rect 13517 6496 13581 6500
rect 13597 6556 13661 6560
rect 13597 6500 13601 6556
rect 13601 6500 13657 6556
rect 13657 6500 13661 6556
rect 13597 6496 13661 6500
rect 4102 6012 4166 6016
rect 4102 5956 4106 6012
rect 4106 5956 4162 6012
rect 4162 5956 4166 6012
rect 4102 5952 4166 5956
rect 4182 6012 4246 6016
rect 4182 5956 4186 6012
rect 4186 5956 4242 6012
rect 4242 5956 4246 6012
rect 4182 5952 4246 5956
rect 4262 6012 4326 6016
rect 4262 5956 4266 6012
rect 4266 5956 4322 6012
rect 4322 5956 4326 6012
rect 4262 5952 4326 5956
rect 4342 6012 4406 6016
rect 4342 5956 4346 6012
rect 4346 5956 4402 6012
rect 4402 5956 4406 6012
rect 4342 5952 4406 5956
rect 7804 6012 7868 6016
rect 7804 5956 7808 6012
rect 7808 5956 7864 6012
rect 7864 5956 7868 6012
rect 7804 5952 7868 5956
rect 7884 6012 7948 6016
rect 7884 5956 7888 6012
rect 7888 5956 7944 6012
rect 7944 5956 7948 6012
rect 7884 5952 7948 5956
rect 7964 6012 8028 6016
rect 7964 5956 7968 6012
rect 7968 5956 8024 6012
rect 8024 5956 8028 6012
rect 7964 5952 8028 5956
rect 8044 6012 8108 6016
rect 8044 5956 8048 6012
rect 8048 5956 8104 6012
rect 8104 5956 8108 6012
rect 8044 5952 8108 5956
rect 11506 6012 11570 6016
rect 11506 5956 11510 6012
rect 11510 5956 11566 6012
rect 11566 5956 11570 6012
rect 11506 5952 11570 5956
rect 11586 6012 11650 6016
rect 11586 5956 11590 6012
rect 11590 5956 11646 6012
rect 11646 5956 11650 6012
rect 11586 5952 11650 5956
rect 11666 6012 11730 6016
rect 11666 5956 11670 6012
rect 11670 5956 11726 6012
rect 11726 5956 11730 6012
rect 11666 5952 11730 5956
rect 11746 6012 11810 6016
rect 11746 5956 11750 6012
rect 11750 5956 11806 6012
rect 11806 5956 11810 6012
rect 11746 5952 11810 5956
rect 15208 6012 15272 6016
rect 15208 5956 15212 6012
rect 15212 5956 15268 6012
rect 15268 5956 15272 6012
rect 15208 5952 15272 5956
rect 15288 6012 15352 6016
rect 15288 5956 15292 6012
rect 15292 5956 15348 6012
rect 15348 5956 15352 6012
rect 15288 5952 15352 5956
rect 15368 6012 15432 6016
rect 15368 5956 15372 6012
rect 15372 5956 15428 6012
rect 15428 5956 15432 6012
rect 15368 5952 15432 5956
rect 15448 6012 15512 6016
rect 15448 5956 15452 6012
rect 15452 5956 15508 6012
rect 15508 5956 15512 6012
rect 15448 5952 15512 5956
rect 2251 5468 2315 5472
rect 2251 5412 2255 5468
rect 2255 5412 2311 5468
rect 2311 5412 2315 5468
rect 2251 5408 2315 5412
rect 2331 5468 2395 5472
rect 2331 5412 2335 5468
rect 2335 5412 2391 5468
rect 2391 5412 2395 5468
rect 2331 5408 2395 5412
rect 2411 5468 2475 5472
rect 2411 5412 2415 5468
rect 2415 5412 2471 5468
rect 2471 5412 2475 5468
rect 2411 5408 2475 5412
rect 2491 5468 2555 5472
rect 2491 5412 2495 5468
rect 2495 5412 2551 5468
rect 2551 5412 2555 5468
rect 2491 5408 2555 5412
rect 5953 5468 6017 5472
rect 5953 5412 5957 5468
rect 5957 5412 6013 5468
rect 6013 5412 6017 5468
rect 5953 5408 6017 5412
rect 6033 5468 6097 5472
rect 6033 5412 6037 5468
rect 6037 5412 6093 5468
rect 6093 5412 6097 5468
rect 6033 5408 6097 5412
rect 6113 5468 6177 5472
rect 6113 5412 6117 5468
rect 6117 5412 6173 5468
rect 6173 5412 6177 5468
rect 6113 5408 6177 5412
rect 6193 5468 6257 5472
rect 6193 5412 6197 5468
rect 6197 5412 6253 5468
rect 6253 5412 6257 5468
rect 6193 5408 6257 5412
rect 9655 5468 9719 5472
rect 9655 5412 9659 5468
rect 9659 5412 9715 5468
rect 9715 5412 9719 5468
rect 9655 5408 9719 5412
rect 9735 5468 9799 5472
rect 9735 5412 9739 5468
rect 9739 5412 9795 5468
rect 9795 5412 9799 5468
rect 9735 5408 9799 5412
rect 9815 5468 9879 5472
rect 9815 5412 9819 5468
rect 9819 5412 9875 5468
rect 9875 5412 9879 5468
rect 9815 5408 9879 5412
rect 9895 5468 9959 5472
rect 9895 5412 9899 5468
rect 9899 5412 9955 5468
rect 9955 5412 9959 5468
rect 9895 5408 9959 5412
rect 13357 5468 13421 5472
rect 13357 5412 13361 5468
rect 13361 5412 13417 5468
rect 13417 5412 13421 5468
rect 13357 5408 13421 5412
rect 13437 5468 13501 5472
rect 13437 5412 13441 5468
rect 13441 5412 13497 5468
rect 13497 5412 13501 5468
rect 13437 5408 13501 5412
rect 13517 5468 13581 5472
rect 13517 5412 13521 5468
rect 13521 5412 13577 5468
rect 13577 5412 13581 5468
rect 13517 5408 13581 5412
rect 13597 5468 13661 5472
rect 13597 5412 13601 5468
rect 13601 5412 13657 5468
rect 13657 5412 13661 5468
rect 13597 5408 13661 5412
rect 4102 4924 4166 4928
rect 4102 4868 4106 4924
rect 4106 4868 4162 4924
rect 4162 4868 4166 4924
rect 4102 4864 4166 4868
rect 4182 4924 4246 4928
rect 4182 4868 4186 4924
rect 4186 4868 4242 4924
rect 4242 4868 4246 4924
rect 4182 4864 4246 4868
rect 4262 4924 4326 4928
rect 4262 4868 4266 4924
rect 4266 4868 4322 4924
rect 4322 4868 4326 4924
rect 4262 4864 4326 4868
rect 4342 4924 4406 4928
rect 4342 4868 4346 4924
rect 4346 4868 4402 4924
rect 4402 4868 4406 4924
rect 4342 4864 4406 4868
rect 7804 4924 7868 4928
rect 7804 4868 7808 4924
rect 7808 4868 7864 4924
rect 7864 4868 7868 4924
rect 7804 4864 7868 4868
rect 7884 4924 7948 4928
rect 7884 4868 7888 4924
rect 7888 4868 7944 4924
rect 7944 4868 7948 4924
rect 7884 4864 7948 4868
rect 7964 4924 8028 4928
rect 7964 4868 7968 4924
rect 7968 4868 8024 4924
rect 8024 4868 8028 4924
rect 7964 4864 8028 4868
rect 8044 4924 8108 4928
rect 8044 4868 8048 4924
rect 8048 4868 8104 4924
rect 8104 4868 8108 4924
rect 8044 4864 8108 4868
rect 11506 4924 11570 4928
rect 11506 4868 11510 4924
rect 11510 4868 11566 4924
rect 11566 4868 11570 4924
rect 11506 4864 11570 4868
rect 11586 4924 11650 4928
rect 11586 4868 11590 4924
rect 11590 4868 11646 4924
rect 11646 4868 11650 4924
rect 11586 4864 11650 4868
rect 11666 4924 11730 4928
rect 11666 4868 11670 4924
rect 11670 4868 11726 4924
rect 11726 4868 11730 4924
rect 11666 4864 11730 4868
rect 11746 4924 11810 4928
rect 11746 4868 11750 4924
rect 11750 4868 11806 4924
rect 11806 4868 11810 4924
rect 11746 4864 11810 4868
rect 15208 4924 15272 4928
rect 15208 4868 15212 4924
rect 15212 4868 15268 4924
rect 15268 4868 15272 4924
rect 15208 4864 15272 4868
rect 15288 4924 15352 4928
rect 15288 4868 15292 4924
rect 15292 4868 15348 4924
rect 15348 4868 15352 4924
rect 15288 4864 15352 4868
rect 15368 4924 15432 4928
rect 15368 4868 15372 4924
rect 15372 4868 15428 4924
rect 15428 4868 15432 4924
rect 15368 4864 15432 4868
rect 15448 4924 15512 4928
rect 15448 4868 15452 4924
rect 15452 4868 15508 4924
rect 15508 4868 15512 4924
rect 15448 4864 15512 4868
rect 2251 4380 2315 4384
rect 2251 4324 2255 4380
rect 2255 4324 2311 4380
rect 2311 4324 2315 4380
rect 2251 4320 2315 4324
rect 2331 4380 2395 4384
rect 2331 4324 2335 4380
rect 2335 4324 2391 4380
rect 2391 4324 2395 4380
rect 2331 4320 2395 4324
rect 2411 4380 2475 4384
rect 2411 4324 2415 4380
rect 2415 4324 2471 4380
rect 2471 4324 2475 4380
rect 2411 4320 2475 4324
rect 2491 4380 2555 4384
rect 2491 4324 2495 4380
rect 2495 4324 2551 4380
rect 2551 4324 2555 4380
rect 2491 4320 2555 4324
rect 5953 4380 6017 4384
rect 5953 4324 5957 4380
rect 5957 4324 6013 4380
rect 6013 4324 6017 4380
rect 5953 4320 6017 4324
rect 6033 4380 6097 4384
rect 6033 4324 6037 4380
rect 6037 4324 6093 4380
rect 6093 4324 6097 4380
rect 6033 4320 6097 4324
rect 6113 4380 6177 4384
rect 6113 4324 6117 4380
rect 6117 4324 6173 4380
rect 6173 4324 6177 4380
rect 6113 4320 6177 4324
rect 6193 4380 6257 4384
rect 6193 4324 6197 4380
rect 6197 4324 6253 4380
rect 6253 4324 6257 4380
rect 6193 4320 6257 4324
rect 9655 4380 9719 4384
rect 9655 4324 9659 4380
rect 9659 4324 9715 4380
rect 9715 4324 9719 4380
rect 9655 4320 9719 4324
rect 9735 4380 9799 4384
rect 9735 4324 9739 4380
rect 9739 4324 9795 4380
rect 9795 4324 9799 4380
rect 9735 4320 9799 4324
rect 9815 4380 9879 4384
rect 9815 4324 9819 4380
rect 9819 4324 9875 4380
rect 9875 4324 9879 4380
rect 9815 4320 9879 4324
rect 9895 4380 9959 4384
rect 9895 4324 9899 4380
rect 9899 4324 9955 4380
rect 9955 4324 9959 4380
rect 9895 4320 9959 4324
rect 13357 4380 13421 4384
rect 13357 4324 13361 4380
rect 13361 4324 13417 4380
rect 13417 4324 13421 4380
rect 13357 4320 13421 4324
rect 13437 4380 13501 4384
rect 13437 4324 13441 4380
rect 13441 4324 13497 4380
rect 13497 4324 13501 4380
rect 13437 4320 13501 4324
rect 13517 4380 13581 4384
rect 13517 4324 13521 4380
rect 13521 4324 13577 4380
rect 13577 4324 13581 4380
rect 13517 4320 13581 4324
rect 13597 4380 13661 4384
rect 13597 4324 13601 4380
rect 13601 4324 13657 4380
rect 13657 4324 13661 4380
rect 13597 4320 13661 4324
rect 4102 3836 4166 3840
rect 4102 3780 4106 3836
rect 4106 3780 4162 3836
rect 4162 3780 4166 3836
rect 4102 3776 4166 3780
rect 4182 3836 4246 3840
rect 4182 3780 4186 3836
rect 4186 3780 4242 3836
rect 4242 3780 4246 3836
rect 4182 3776 4246 3780
rect 4262 3836 4326 3840
rect 4262 3780 4266 3836
rect 4266 3780 4322 3836
rect 4322 3780 4326 3836
rect 4262 3776 4326 3780
rect 4342 3836 4406 3840
rect 4342 3780 4346 3836
rect 4346 3780 4402 3836
rect 4402 3780 4406 3836
rect 4342 3776 4406 3780
rect 7804 3836 7868 3840
rect 7804 3780 7808 3836
rect 7808 3780 7864 3836
rect 7864 3780 7868 3836
rect 7804 3776 7868 3780
rect 7884 3836 7948 3840
rect 7884 3780 7888 3836
rect 7888 3780 7944 3836
rect 7944 3780 7948 3836
rect 7884 3776 7948 3780
rect 7964 3836 8028 3840
rect 7964 3780 7968 3836
rect 7968 3780 8024 3836
rect 8024 3780 8028 3836
rect 7964 3776 8028 3780
rect 8044 3836 8108 3840
rect 8044 3780 8048 3836
rect 8048 3780 8104 3836
rect 8104 3780 8108 3836
rect 8044 3776 8108 3780
rect 11506 3836 11570 3840
rect 11506 3780 11510 3836
rect 11510 3780 11566 3836
rect 11566 3780 11570 3836
rect 11506 3776 11570 3780
rect 11586 3836 11650 3840
rect 11586 3780 11590 3836
rect 11590 3780 11646 3836
rect 11646 3780 11650 3836
rect 11586 3776 11650 3780
rect 11666 3836 11730 3840
rect 11666 3780 11670 3836
rect 11670 3780 11726 3836
rect 11726 3780 11730 3836
rect 11666 3776 11730 3780
rect 11746 3836 11810 3840
rect 11746 3780 11750 3836
rect 11750 3780 11806 3836
rect 11806 3780 11810 3836
rect 11746 3776 11810 3780
rect 15208 3836 15272 3840
rect 15208 3780 15212 3836
rect 15212 3780 15268 3836
rect 15268 3780 15272 3836
rect 15208 3776 15272 3780
rect 15288 3836 15352 3840
rect 15288 3780 15292 3836
rect 15292 3780 15348 3836
rect 15348 3780 15352 3836
rect 15288 3776 15352 3780
rect 15368 3836 15432 3840
rect 15368 3780 15372 3836
rect 15372 3780 15428 3836
rect 15428 3780 15432 3836
rect 15368 3776 15432 3780
rect 15448 3836 15512 3840
rect 15448 3780 15452 3836
rect 15452 3780 15508 3836
rect 15508 3780 15512 3836
rect 15448 3776 15512 3780
rect 2251 3292 2315 3296
rect 2251 3236 2255 3292
rect 2255 3236 2311 3292
rect 2311 3236 2315 3292
rect 2251 3232 2315 3236
rect 2331 3292 2395 3296
rect 2331 3236 2335 3292
rect 2335 3236 2391 3292
rect 2391 3236 2395 3292
rect 2331 3232 2395 3236
rect 2411 3292 2475 3296
rect 2411 3236 2415 3292
rect 2415 3236 2471 3292
rect 2471 3236 2475 3292
rect 2411 3232 2475 3236
rect 2491 3292 2555 3296
rect 2491 3236 2495 3292
rect 2495 3236 2551 3292
rect 2551 3236 2555 3292
rect 2491 3232 2555 3236
rect 5953 3292 6017 3296
rect 5953 3236 5957 3292
rect 5957 3236 6013 3292
rect 6013 3236 6017 3292
rect 5953 3232 6017 3236
rect 6033 3292 6097 3296
rect 6033 3236 6037 3292
rect 6037 3236 6093 3292
rect 6093 3236 6097 3292
rect 6033 3232 6097 3236
rect 6113 3292 6177 3296
rect 6113 3236 6117 3292
rect 6117 3236 6173 3292
rect 6173 3236 6177 3292
rect 6113 3232 6177 3236
rect 6193 3292 6257 3296
rect 6193 3236 6197 3292
rect 6197 3236 6253 3292
rect 6253 3236 6257 3292
rect 6193 3232 6257 3236
rect 9655 3292 9719 3296
rect 9655 3236 9659 3292
rect 9659 3236 9715 3292
rect 9715 3236 9719 3292
rect 9655 3232 9719 3236
rect 9735 3292 9799 3296
rect 9735 3236 9739 3292
rect 9739 3236 9795 3292
rect 9795 3236 9799 3292
rect 9735 3232 9799 3236
rect 9815 3292 9879 3296
rect 9815 3236 9819 3292
rect 9819 3236 9875 3292
rect 9875 3236 9879 3292
rect 9815 3232 9879 3236
rect 9895 3292 9959 3296
rect 9895 3236 9899 3292
rect 9899 3236 9955 3292
rect 9955 3236 9959 3292
rect 9895 3232 9959 3236
rect 13357 3292 13421 3296
rect 13357 3236 13361 3292
rect 13361 3236 13417 3292
rect 13417 3236 13421 3292
rect 13357 3232 13421 3236
rect 13437 3292 13501 3296
rect 13437 3236 13441 3292
rect 13441 3236 13497 3292
rect 13497 3236 13501 3292
rect 13437 3232 13501 3236
rect 13517 3292 13581 3296
rect 13517 3236 13521 3292
rect 13521 3236 13577 3292
rect 13577 3236 13581 3292
rect 13517 3232 13581 3236
rect 13597 3292 13661 3296
rect 13597 3236 13601 3292
rect 13601 3236 13657 3292
rect 13657 3236 13661 3292
rect 13597 3232 13661 3236
rect 4102 2748 4166 2752
rect 4102 2692 4106 2748
rect 4106 2692 4162 2748
rect 4162 2692 4166 2748
rect 4102 2688 4166 2692
rect 4182 2748 4246 2752
rect 4182 2692 4186 2748
rect 4186 2692 4242 2748
rect 4242 2692 4246 2748
rect 4182 2688 4246 2692
rect 4262 2748 4326 2752
rect 4262 2692 4266 2748
rect 4266 2692 4322 2748
rect 4322 2692 4326 2748
rect 4262 2688 4326 2692
rect 4342 2748 4406 2752
rect 4342 2692 4346 2748
rect 4346 2692 4402 2748
rect 4402 2692 4406 2748
rect 4342 2688 4406 2692
rect 7804 2748 7868 2752
rect 7804 2692 7808 2748
rect 7808 2692 7864 2748
rect 7864 2692 7868 2748
rect 7804 2688 7868 2692
rect 7884 2748 7948 2752
rect 7884 2692 7888 2748
rect 7888 2692 7944 2748
rect 7944 2692 7948 2748
rect 7884 2688 7948 2692
rect 7964 2748 8028 2752
rect 7964 2692 7968 2748
rect 7968 2692 8024 2748
rect 8024 2692 8028 2748
rect 7964 2688 8028 2692
rect 8044 2748 8108 2752
rect 8044 2692 8048 2748
rect 8048 2692 8104 2748
rect 8104 2692 8108 2748
rect 8044 2688 8108 2692
rect 11506 2748 11570 2752
rect 11506 2692 11510 2748
rect 11510 2692 11566 2748
rect 11566 2692 11570 2748
rect 11506 2688 11570 2692
rect 11586 2748 11650 2752
rect 11586 2692 11590 2748
rect 11590 2692 11646 2748
rect 11646 2692 11650 2748
rect 11586 2688 11650 2692
rect 11666 2748 11730 2752
rect 11666 2692 11670 2748
rect 11670 2692 11726 2748
rect 11726 2692 11730 2748
rect 11666 2688 11730 2692
rect 11746 2748 11810 2752
rect 11746 2692 11750 2748
rect 11750 2692 11806 2748
rect 11806 2692 11810 2748
rect 11746 2688 11810 2692
rect 15208 2748 15272 2752
rect 15208 2692 15212 2748
rect 15212 2692 15268 2748
rect 15268 2692 15272 2748
rect 15208 2688 15272 2692
rect 15288 2748 15352 2752
rect 15288 2692 15292 2748
rect 15292 2692 15348 2748
rect 15348 2692 15352 2748
rect 15288 2688 15352 2692
rect 15368 2748 15432 2752
rect 15368 2692 15372 2748
rect 15372 2692 15428 2748
rect 15428 2692 15432 2748
rect 15368 2688 15432 2692
rect 15448 2748 15512 2752
rect 15448 2692 15452 2748
rect 15452 2692 15508 2748
rect 15508 2692 15512 2748
rect 15448 2688 15512 2692
rect 2251 2204 2315 2208
rect 2251 2148 2255 2204
rect 2255 2148 2311 2204
rect 2311 2148 2315 2204
rect 2251 2144 2315 2148
rect 2331 2204 2395 2208
rect 2331 2148 2335 2204
rect 2335 2148 2391 2204
rect 2391 2148 2395 2204
rect 2331 2144 2395 2148
rect 2411 2204 2475 2208
rect 2411 2148 2415 2204
rect 2415 2148 2471 2204
rect 2471 2148 2475 2204
rect 2411 2144 2475 2148
rect 2491 2204 2555 2208
rect 2491 2148 2495 2204
rect 2495 2148 2551 2204
rect 2551 2148 2555 2204
rect 2491 2144 2555 2148
rect 5953 2204 6017 2208
rect 5953 2148 5957 2204
rect 5957 2148 6013 2204
rect 6013 2148 6017 2204
rect 5953 2144 6017 2148
rect 6033 2204 6097 2208
rect 6033 2148 6037 2204
rect 6037 2148 6093 2204
rect 6093 2148 6097 2204
rect 6033 2144 6097 2148
rect 6113 2204 6177 2208
rect 6113 2148 6117 2204
rect 6117 2148 6173 2204
rect 6173 2148 6177 2204
rect 6113 2144 6177 2148
rect 6193 2204 6257 2208
rect 6193 2148 6197 2204
rect 6197 2148 6253 2204
rect 6253 2148 6257 2204
rect 6193 2144 6257 2148
rect 9655 2204 9719 2208
rect 9655 2148 9659 2204
rect 9659 2148 9715 2204
rect 9715 2148 9719 2204
rect 9655 2144 9719 2148
rect 9735 2204 9799 2208
rect 9735 2148 9739 2204
rect 9739 2148 9795 2204
rect 9795 2148 9799 2204
rect 9735 2144 9799 2148
rect 9815 2204 9879 2208
rect 9815 2148 9819 2204
rect 9819 2148 9875 2204
rect 9875 2148 9879 2204
rect 9815 2144 9879 2148
rect 9895 2204 9959 2208
rect 9895 2148 9899 2204
rect 9899 2148 9955 2204
rect 9955 2148 9959 2204
rect 9895 2144 9959 2148
rect 13357 2204 13421 2208
rect 13357 2148 13361 2204
rect 13361 2148 13417 2204
rect 13417 2148 13421 2204
rect 13357 2144 13421 2148
rect 13437 2204 13501 2208
rect 13437 2148 13441 2204
rect 13441 2148 13497 2204
rect 13497 2148 13501 2204
rect 13437 2144 13501 2148
rect 13517 2204 13581 2208
rect 13517 2148 13521 2204
rect 13521 2148 13577 2204
rect 13577 2148 13581 2204
rect 13517 2144 13581 2148
rect 13597 2204 13661 2208
rect 13597 2148 13601 2204
rect 13601 2148 13657 2204
rect 13657 2148 13661 2204
rect 13597 2144 13661 2148
rect 4102 1660 4166 1664
rect 4102 1604 4106 1660
rect 4106 1604 4162 1660
rect 4162 1604 4166 1660
rect 4102 1600 4166 1604
rect 4182 1660 4246 1664
rect 4182 1604 4186 1660
rect 4186 1604 4242 1660
rect 4242 1604 4246 1660
rect 4182 1600 4246 1604
rect 4262 1660 4326 1664
rect 4262 1604 4266 1660
rect 4266 1604 4322 1660
rect 4322 1604 4326 1660
rect 4262 1600 4326 1604
rect 4342 1660 4406 1664
rect 4342 1604 4346 1660
rect 4346 1604 4402 1660
rect 4402 1604 4406 1660
rect 4342 1600 4406 1604
rect 7804 1660 7868 1664
rect 7804 1604 7808 1660
rect 7808 1604 7864 1660
rect 7864 1604 7868 1660
rect 7804 1600 7868 1604
rect 7884 1660 7948 1664
rect 7884 1604 7888 1660
rect 7888 1604 7944 1660
rect 7944 1604 7948 1660
rect 7884 1600 7948 1604
rect 7964 1660 8028 1664
rect 7964 1604 7968 1660
rect 7968 1604 8024 1660
rect 8024 1604 8028 1660
rect 7964 1600 8028 1604
rect 8044 1660 8108 1664
rect 8044 1604 8048 1660
rect 8048 1604 8104 1660
rect 8104 1604 8108 1660
rect 8044 1600 8108 1604
rect 11506 1660 11570 1664
rect 11506 1604 11510 1660
rect 11510 1604 11566 1660
rect 11566 1604 11570 1660
rect 11506 1600 11570 1604
rect 11586 1660 11650 1664
rect 11586 1604 11590 1660
rect 11590 1604 11646 1660
rect 11646 1604 11650 1660
rect 11586 1600 11650 1604
rect 11666 1660 11730 1664
rect 11666 1604 11670 1660
rect 11670 1604 11726 1660
rect 11726 1604 11730 1660
rect 11666 1600 11730 1604
rect 11746 1660 11810 1664
rect 11746 1604 11750 1660
rect 11750 1604 11806 1660
rect 11806 1604 11810 1660
rect 11746 1600 11810 1604
rect 15208 1660 15272 1664
rect 15208 1604 15212 1660
rect 15212 1604 15268 1660
rect 15268 1604 15272 1660
rect 15208 1600 15272 1604
rect 15288 1660 15352 1664
rect 15288 1604 15292 1660
rect 15292 1604 15348 1660
rect 15348 1604 15352 1660
rect 15288 1600 15352 1604
rect 15368 1660 15432 1664
rect 15368 1604 15372 1660
rect 15372 1604 15428 1660
rect 15428 1604 15432 1660
rect 15368 1600 15432 1604
rect 15448 1660 15512 1664
rect 15448 1604 15452 1660
rect 15452 1604 15508 1660
rect 15508 1604 15512 1660
rect 15448 1600 15512 1604
rect 2251 1116 2315 1120
rect 2251 1060 2255 1116
rect 2255 1060 2311 1116
rect 2311 1060 2315 1116
rect 2251 1056 2315 1060
rect 2331 1116 2395 1120
rect 2331 1060 2335 1116
rect 2335 1060 2391 1116
rect 2391 1060 2395 1116
rect 2331 1056 2395 1060
rect 2411 1116 2475 1120
rect 2411 1060 2415 1116
rect 2415 1060 2471 1116
rect 2471 1060 2475 1116
rect 2411 1056 2475 1060
rect 2491 1116 2555 1120
rect 2491 1060 2495 1116
rect 2495 1060 2551 1116
rect 2551 1060 2555 1116
rect 2491 1056 2555 1060
rect 5953 1116 6017 1120
rect 5953 1060 5957 1116
rect 5957 1060 6013 1116
rect 6013 1060 6017 1116
rect 5953 1056 6017 1060
rect 6033 1116 6097 1120
rect 6033 1060 6037 1116
rect 6037 1060 6093 1116
rect 6093 1060 6097 1116
rect 6033 1056 6097 1060
rect 6113 1116 6177 1120
rect 6113 1060 6117 1116
rect 6117 1060 6173 1116
rect 6173 1060 6177 1116
rect 6113 1056 6177 1060
rect 6193 1116 6257 1120
rect 6193 1060 6197 1116
rect 6197 1060 6253 1116
rect 6253 1060 6257 1116
rect 6193 1056 6257 1060
rect 9655 1116 9719 1120
rect 9655 1060 9659 1116
rect 9659 1060 9715 1116
rect 9715 1060 9719 1116
rect 9655 1056 9719 1060
rect 9735 1116 9799 1120
rect 9735 1060 9739 1116
rect 9739 1060 9795 1116
rect 9795 1060 9799 1116
rect 9735 1056 9799 1060
rect 9815 1116 9879 1120
rect 9815 1060 9819 1116
rect 9819 1060 9875 1116
rect 9875 1060 9879 1116
rect 9815 1056 9879 1060
rect 9895 1116 9959 1120
rect 9895 1060 9899 1116
rect 9899 1060 9955 1116
rect 9955 1060 9959 1116
rect 9895 1056 9959 1060
rect 13357 1116 13421 1120
rect 13357 1060 13361 1116
rect 13361 1060 13417 1116
rect 13417 1060 13421 1116
rect 13357 1056 13421 1060
rect 13437 1116 13501 1120
rect 13437 1060 13441 1116
rect 13441 1060 13497 1116
rect 13497 1060 13501 1116
rect 13437 1056 13501 1060
rect 13517 1116 13581 1120
rect 13517 1060 13521 1116
rect 13521 1060 13577 1116
rect 13577 1060 13581 1116
rect 13517 1056 13581 1060
rect 13597 1116 13661 1120
rect 13597 1060 13601 1116
rect 13601 1060 13657 1116
rect 13657 1060 13661 1116
rect 13597 1056 13661 1060
rect 4102 572 4166 576
rect 4102 516 4106 572
rect 4106 516 4162 572
rect 4162 516 4166 572
rect 4102 512 4166 516
rect 4182 572 4246 576
rect 4182 516 4186 572
rect 4186 516 4242 572
rect 4242 516 4246 572
rect 4182 512 4246 516
rect 4262 572 4326 576
rect 4262 516 4266 572
rect 4266 516 4322 572
rect 4322 516 4326 572
rect 4262 512 4326 516
rect 4342 572 4406 576
rect 4342 516 4346 572
rect 4346 516 4402 572
rect 4402 516 4406 572
rect 4342 512 4406 516
rect 7804 572 7868 576
rect 7804 516 7808 572
rect 7808 516 7864 572
rect 7864 516 7868 572
rect 7804 512 7868 516
rect 7884 572 7948 576
rect 7884 516 7888 572
rect 7888 516 7944 572
rect 7944 516 7948 572
rect 7884 512 7948 516
rect 7964 572 8028 576
rect 7964 516 7968 572
rect 7968 516 8024 572
rect 8024 516 8028 572
rect 7964 512 8028 516
rect 8044 572 8108 576
rect 8044 516 8048 572
rect 8048 516 8104 572
rect 8104 516 8108 572
rect 8044 512 8108 516
rect 11506 572 11570 576
rect 11506 516 11510 572
rect 11510 516 11566 572
rect 11566 516 11570 572
rect 11506 512 11570 516
rect 11586 572 11650 576
rect 11586 516 11590 572
rect 11590 516 11646 572
rect 11646 516 11650 572
rect 11586 512 11650 516
rect 11666 572 11730 576
rect 11666 516 11670 572
rect 11670 516 11726 572
rect 11726 516 11730 572
rect 11666 512 11730 516
rect 11746 572 11810 576
rect 11746 516 11750 572
rect 11750 516 11806 572
rect 11806 516 11810 572
rect 11746 512 11810 516
rect 15208 572 15272 576
rect 15208 516 15212 572
rect 15212 516 15268 572
rect 15268 516 15272 572
rect 15208 512 15272 516
rect 15288 572 15352 576
rect 15288 516 15292 572
rect 15292 516 15348 572
rect 15348 516 15352 572
rect 15288 512 15352 516
rect 15368 572 15432 576
rect 15368 516 15372 572
rect 15372 516 15428 572
rect 15428 516 15432 572
rect 15368 512 15432 516
rect 15448 572 15512 576
rect 15448 516 15452 572
rect 15452 516 15508 572
rect 15508 516 15512 572
rect 15448 512 15512 516
<< metal4 >>
rect 2243 15264 2563 15280
rect 2243 15200 2251 15264
rect 2315 15200 2331 15264
rect 2395 15200 2411 15264
rect 2475 15200 2491 15264
rect 2555 15200 2563 15264
rect 2243 14176 2563 15200
rect 2243 14112 2251 14176
rect 2315 14112 2331 14176
rect 2395 14112 2411 14176
rect 2475 14112 2491 14176
rect 2555 14112 2563 14176
rect 2243 13088 2563 14112
rect 2243 13024 2251 13088
rect 2315 13024 2331 13088
rect 2395 13024 2411 13088
rect 2475 13024 2491 13088
rect 2555 13024 2563 13088
rect 2243 12000 2563 13024
rect 2243 11936 2251 12000
rect 2315 11936 2331 12000
rect 2395 11936 2411 12000
rect 2475 11936 2491 12000
rect 2555 11936 2563 12000
rect 2243 10912 2563 11936
rect 2243 10848 2251 10912
rect 2315 10848 2331 10912
rect 2395 10848 2411 10912
rect 2475 10848 2491 10912
rect 2555 10848 2563 10912
rect 2243 9824 2563 10848
rect 2243 9760 2251 9824
rect 2315 9760 2331 9824
rect 2395 9760 2411 9824
rect 2475 9760 2491 9824
rect 2555 9760 2563 9824
rect 2243 8736 2563 9760
rect 2243 8672 2251 8736
rect 2315 8672 2331 8736
rect 2395 8672 2411 8736
rect 2475 8672 2491 8736
rect 2555 8672 2563 8736
rect 2243 7648 2563 8672
rect 2243 7584 2251 7648
rect 2315 7584 2331 7648
rect 2395 7584 2411 7648
rect 2475 7584 2491 7648
rect 2555 7584 2563 7648
rect 2243 6560 2563 7584
rect 2243 6496 2251 6560
rect 2315 6496 2331 6560
rect 2395 6496 2411 6560
rect 2475 6496 2491 6560
rect 2555 6496 2563 6560
rect 2243 5472 2563 6496
rect 2243 5408 2251 5472
rect 2315 5408 2331 5472
rect 2395 5408 2411 5472
rect 2475 5408 2491 5472
rect 2555 5408 2563 5472
rect 2243 4384 2563 5408
rect 2243 4320 2251 4384
rect 2315 4320 2331 4384
rect 2395 4320 2411 4384
rect 2475 4320 2491 4384
rect 2555 4320 2563 4384
rect 2243 3296 2563 4320
rect 2243 3232 2251 3296
rect 2315 3232 2331 3296
rect 2395 3232 2411 3296
rect 2475 3232 2491 3296
rect 2555 3232 2563 3296
rect 2243 2208 2563 3232
rect 2243 2144 2251 2208
rect 2315 2144 2331 2208
rect 2395 2144 2411 2208
rect 2475 2144 2491 2208
rect 2555 2144 2563 2208
rect 2243 1120 2563 2144
rect 2243 1056 2251 1120
rect 2315 1056 2331 1120
rect 2395 1056 2411 1120
rect 2475 1056 2491 1120
rect 2555 1056 2563 1120
rect 2243 496 2563 1056
rect 4094 14720 4414 15280
rect 4094 14656 4102 14720
rect 4166 14656 4182 14720
rect 4246 14656 4262 14720
rect 4326 14656 4342 14720
rect 4406 14656 4414 14720
rect 4094 13632 4414 14656
rect 4094 13568 4102 13632
rect 4166 13568 4182 13632
rect 4246 13568 4262 13632
rect 4326 13568 4342 13632
rect 4406 13568 4414 13632
rect 4094 12544 4414 13568
rect 4094 12480 4102 12544
rect 4166 12480 4182 12544
rect 4246 12480 4262 12544
rect 4326 12480 4342 12544
rect 4406 12480 4414 12544
rect 4094 11456 4414 12480
rect 4094 11392 4102 11456
rect 4166 11392 4182 11456
rect 4246 11392 4262 11456
rect 4326 11392 4342 11456
rect 4406 11392 4414 11456
rect 4094 10368 4414 11392
rect 4094 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4342 10368
rect 4406 10304 4414 10368
rect 4094 9280 4414 10304
rect 4094 9216 4102 9280
rect 4166 9216 4182 9280
rect 4246 9216 4262 9280
rect 4326 9216 4342 9280
rect 4406 9216 4414 9280
rect 4094 8192 4414 9216
rect 4094 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4342 8192
rect 4406 8128 4414 8192
rect 4094 7104 4414 8128
rect 4094 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4342 7104
rect 4406 7040 4414 7104
rect 4094 6016 4414 7040
rect 4094 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4342 6016
rect 4406 5952 4414 6016
rect 4094 4928 4414 5952
rect 4094 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4342 4928
rect 4406 4864 4414 4928
rect 4094 3840 4414 4864
rect 4094 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4342 3840
rect 4406 3776 4414 3840
rect 4094 2752 4414 3776
rect 4094 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4342 2752
rect 4406 2688 4414 2752
rect 4094 1664 4414 2688
rect 4094 1600 4102 1664
rect 4166 1600 4182 1664
rect 4246 1600 4262 1664
rect 4326 1600 4342 1664
rect 4406 1600 4414 1664
rect 4094 576 4414 1600
rect 4094 512 4102 576
rect 4166 512 4182 576
rect 4246 512 4262 576
rect 4326 512 4342 576
rect 4406 512 4414 576
rect 4094 496 4414 512
rect 5945 15264 6265 15280
rect 5945 15200 5953 15264
rect 6017 15200 6033 15264
rect 6097 15200 6113 15264
rect 6177 15200 6193 15264
rect 6257 15200 6265 15264
rect 5945 14176 6265 15200
rect 5945 14112 5953 14176
rect 6017 14112 6033 14176
rect 6097 14112 6113 14176
rect 6177 14112 6193 14176
rect 6257 14112 6265 14176
rect 5945 13088 6265 14112
rect 5945 13024 5953 13088
rect 6017 13024 6033 13088
rect 6097 13024 6113 13088
rect 6177 13024 6193 13088
rect 6257 13024 6265 13088
rect 5945 12000 6265 13024
rect 5945 11936 5953 12000
rect 6017 11936 6033 12000
rect 6097 11936 6113 12000
rect 6177 11936 6193 12000
rect 6257 11936 6265 12000
rect 5945 10912 6265 11936
rect 5945 10848 5953 10912
rect 6017 10848 6033 10912
rect 6097 10848 6113 10912
rect 6177 10848 6193 10912
rect 6257 10848 6265 10912
rect 5945 9824 6265 10848
rect 5945 9760 5953 9824
rect 6017 9760 6033 9824
rect 6097 9760 6113 9824
rect 6177 9760 6193 9824
rect 6257 9760 6265 9824
rect 5945 8736 6265 9760
rect 5945 8672 5953 8736
rect 6017 8672 6033 8736
rect 6097 8672 6113 8736
rect 6177 8672 6193 8736
rect 6257 8672 6265 8736
rect 5945 7648 6265 8672
rect 5945 7584 5953 7648
rect 6017 7584 6033 7648
rect 6097 7584 6113 7648
rect 6177 7584 6193 7648
rect 6257 7584 6265 7648
rect 5945 6560 6265 7584
rect 5945 6496 5953 6560
rect 6017 6496 6033 6560
rect 6097 6496 6113 6560
rect 6177 6496 6193 6560
rect 6257 6496 6265 6560
rect 5945 5472 6265 6496
rect 5945 5408 5953 5472
rect 6017 5408 6033 5472
rect 6097 5408 6113 5472
rect 6177 5408 6193 5472
rect 6257 5408 6265 5472
rect 5945 4384 6265 5408
rect 5945 4320 5953 4384
rect 6017 4320 6033 4384
rect 6097 4320 6113 4384
rect 6177 4320 6193 4384
rect 6257 4320 6265 4384
rect 5945 3296 6265 4320
rect 5945 3232 5953 3296
rect 6017 3232 6033 3296
rect 6097 3232 6113 3296
rect 6177 3232 6193 3296
rect 6257 3232 6265 3296
rect 5945 2208 6265 3232
rect 5945 2144 5953 2208
rect 6017 2144 6033 2208
rect 6097 2144 6113 2208
rect 6177 2144 6193 2208
rect 6257 2144 6265 2208
rect 5945 1120 6265 2144
rect 5945 1056 5953 1120
rect 6017 1056 6033 1120
rect 6097 1056 6113 1120
rect 6177 1056 6193 1120
rect 6257 1056 6265 1120
rect 5945 496 6265 1056
rect 7796 14720 8116 15280
rect 7796 14656 7804 14720
rect 7868 14656 7884 14720
rect 7948 14656 7964 14720
rect 8028 14656 8044 14720
rect 8108 14656 8116 14720
rect 7796 13632 8116 14656
rect 7796 13568 7804 13632
rect 7868 13568 7884 13632
rect 7948 13568 7964 13632
rect 8028 13568 8044 13632
rect 8108 13568 8116 13632
rect 7796 12544 8116 13568
rect 7796 12480 7804 12544
rect 7868 12480 7884 12544
rect 7948 12480 7964 12544
rect 8028 12480 8044 12544
rect 8108 12480 8116 12544
rect 7796 11456 8116 12480
rect 7796 11392 7804 11456
rect 7868 11392 7884 11456
rect 7948 11392 7964 11456
rect 8028 11392 8044 11456
rect 8108 11392 8116 11456
rect 7796 10368 8116 11392
rect 7796 10304 7804 10368
rect 7868 10304 7884 10368
rect 7948 10304 7964 10368
rect 8028 10304 8044 10368
rect 8108 10304 8116 10368
rect 7796 9280 8116 10304
rect 7796 9216 7804 9280
rect 7868 9216 7884 9280
rect 7948 9216 7964 9280
rect 8028 9216 8044 9280
rect 8108 9216 8116 9280
rect 7796 8192 8116 9216
rect 7796 8128 7804 8192
rect 7868 8128 7884 8192
rect 7948 8128 7964 8192
rect 8028 8128 8044 8192
rect 8108 8128 8116 8192
rect 7796 7104 8116 8128
rect 7796 7040 7804 7104
rect 7868 7040 7884 7104
rect 7948 7040 7964 7104
rect 8028 7040 8044 7104
rect 8108 7040 8116 7104
rect 7796 6016 8116 7040
rect 7796 5952 7804 6016
rect 7868 5952 7884 6016
rect 7948 5952 7964 6016
rect 8028 5952 8044 6016
rect 8108 5952 8116 6016
rect 7796 4928 8116 5952
rect 7796 4864 7804 4928
rect 7868 4864 7884 4928
rect 7948 4864 7964 4928
rect 8028 4864 8044 4928
rect 8108 4864 8116 4928
rect 7796 3840 8116 4864
rect 7796 3776 7804 3840
rect 7868 3776 7884 3840
rect 7948 3776 7964 3840
rect 8028 3776 8044 3840
rect 8108 3776 8116 3840
rect 7796 2752 8116 3776
rect 7796 2688 7804 2752
rect 7868 2688 7884 2752
rect 7948 2688 7964 2752
rect 8028 2688 8044 2752
rect 8108 2688 8116 2752
rect 7796 1664 8116 2688
rect 7796 1600 7804 1664
rect 7868 1600 7884 1664
rect 7948 1600 7964 1664
rect 8028 1600 8044 1664
rect 8108 1600 8116 1664
rect 7796 576 8116 1600
rect 7796 512 7804 576
rect 7868 512 7884 576
rect 7948 512 7964 576
rect 8028 512 8044 576
rect 8108 512 8116 576
rect 7796 496 8116 512
rect 9647 15264 9967 15280
rect 9647 15200 9655 15264
rect 9719 15200 9735 15264
rect 9799 15200 9815 15264
rect 9879 15200 9895 15264
rect 9959 15200 9967 15264
rect 9647 14176 9967 15200
rect 9647 14112 9655 14176
rect 9719 14112 9735 14176
rect 9799 14112 9815 14176
rect 9879 14112 9895 14176
rect 9959 14112 9967 14176
rect 9647 13088 9967 14112
rect 9647 13024 9655 13088
rect 9719 13024 9735 13088
rect 9799 13024 9815 13088
rect 9879 13024 9895 13088
rect 9959 13024 9967 13088
rect 9647 12000 9967 13024
rect 9647 11936 9655 12000
rect 9719 11936 9735 12000
rect 9799 11936 9815 12000
rect 9879 11936 9895 12000
rect 9959 11936 9967 12000
rect 9647 10912 9967 11936
rect 9647 10848 9655 10912
rect 9719 10848 9735 10912
rect 9799 10848 9815 10912
rect 9879 10848 9895 10912
rect 9959 10848 9967 10912
rect 9647 9824 9967 10848
rect 9647 9760 9655 9824
rect 9719 9760 9735 9824
rect 9799 9760 9815 9824
rect 9879 9760 9895 9824
rect 9959 9760 9967 9824
rect 9647 8736 9967 9760
rect 9647 8672 9655 8736
rect 9719 8672 9735 8736
rect 9799 8672 9815 8736
rect 9879 8672 9895 8736
rect 9959 8672 9967 8736
rect 9647 7648 9967 8672
rect 9647 7584 9655 7648
rect 9719 7584 9735 7648
rect 9799 7584 9815 7648
rect 9879 7584 9895 7648
rect 9959 7584 9967 7648
rect 9647 6560 9967 7584
rect 9647 6496 9655 6560
rect 9719 6496 9735 6560
rect 9799 6496 9815 6560
rect 9879 6496 9895 6560
rect 9959 6496 9967 6560
rect 9647 5472 9967 6496
rect 9647 5408 9655 5472
rect 9719 5408 9735 5472
rect 9799 5408 9815 5472
rect 9879 5408 9895 5472
rect 9959 5408 9967 5472
rect 9647 4384 9967 5408
rect 9647 4320 9655 4384
rect 9719 4320 9735 4384
rect 9799 4320 9815 4384
rect 9879 4320 9895 4384
rect 9959 4320 9967 4384
rect 9647 3296 9967 4320
rect 9647 3232 9655 3296
rect 9719 3232 9735 3296
rect 9799 3232 9815 3296
rect 9879 3232 9895 3296
rect 9959 3232 9967 3296
rect 9647 2208 9967 3232
rect 9647 2144 9655 2208
rect 9719 2144 9735 2208
rect 9799 2144 9815 2208
rect 9879 2144 9895 2208
rect 9959 2144 9967 2208
rect 9647 1120 9967 2144
rect 9647 1056 9655 1120
rect 9719 1056 9735 1120
rect 9799 1056 9815 1120
rect 9879 1056 9895 1120
rect 9959 1056 9967 1120
rect 9647 496 9967 1056
rect 11498 14720 11818 15280
rect 11498 14656 11506 14720
rect 11570 14656 11586 14720
rect 11650 14656 11666 14720
rect 11730 14656 11746 14720
rect 11810 14656 11818 14720
rect 11498 13632 11818 14656
rect 11498 13568 11506 13632
rect 11570 13568 11586 13632
rect 11650 13568 11666 13632
rect 11730 13568 11746 13632
rect 11810 13568 11818 13632
rect 11498 12544 11818 13568
rect 11498 12480 11506 12544
rect 11570 12480 11586 12544
rect 11650 12480 11666 12544
rect 11730 12480 11746 12544
rect 11810 12480 11818 12544
rect 11498 11456 11818 12480
rect 11498 11392 11506 11456
rect 11570 11392 11586 11456
rect 11650 11392 11666 11456
rect 11730 11392 11746 11456
rect 11810 11392 11818 11456
rect 11498 10368 11818 11392
rect 11498 10304 11506 10368
rect 11570 10304 11586 10368
rect 11650 10304 11666 10368
rect 11730 10304 11746 10368
rect 11810 10304 11818 10368
rect 11498 9280 11818 10304
rect 11498 9216 11506 9280
rect 11570 9216 11586 9280
rect 11650 9216 11666 9280
rect 11730 9216 11746 9280
rect 11810 9216 11818 9280
rect 11498 8192 11818 9216
rect 11498 8128 11506 8192
rect 11570 8128 11586 8192
rect 11650 8128 11666 8192
rect 11730 8128 11746 8192
rect 11810 8128 11818 8192
rect 11498 7104 11818 8128
rect 11498 7040 11506 7104
rect 11570 7040 11586 7104
rect 11650 7040 11666 7104
rect 11730 7040 11746 7104
rect 11810 7040 11818 7104
rect 11498 6016 11818 7040
rect 11498 5952 11506 6016
rect 11570 5952 11586 6016
rect 11650 5952 11666 6016
rect 11730 5952 11746 6016
rect 11810 5952 11818 6016
rect 11498 4928 11818 5952
rect 11498 4864 11506 4928
rect 11570 4864 11586 4928
rect 11650 4864 11666 4928
rect 11730 4864 11746 4928
rect 11810 4864 11818 4928
rect 11498 3840 11818 4864
rect 11498 3776 11506 3840
rect 11570 3776 11586 3840
rect 11650 3776 11666 3840
rect 11730 3776 11746 3840
rect 11810 3776 11818 3840
rect 11498 2752 11818 3776
rect 11498 2688 11506 2752
rect 11570 2688 11586 2752
rect 11650 2688 11666 2752
rect 11730 2688 11746 2752
rect 11810 2688 11818 2752
rect 11498 1664 11818 2688
rect 11498 1600 11506 1664
rect 11570 1600 11586 1664
rect 11650 1600 11666 1664
rect 11730 1600 11746 1664
rect 11810 1600 11818 1664
rect 11498 576 11818 1600
rect 11498 512 11506 576
rect 11570 512 11586 576
rect 11650 512 11666 576
rect 11730 512 11746 576
rect 11810 512 11818 576
rect 11498 496 11818 512
rect 13349 15264 13669 15280
rect 13349 15200 13357 15264
rect 13421 15200 13437 15264
rect 13501 15200 13517 15264
rect 13581 15200 13597 15264
rect 13661 15200 13669 15264
rect 13349 14176 13669 15200
rect 13349 14112 13357 14176
rect 13421 14112 13437 14176
rect 13501 14112 13517 14176
rect 13581 14112 13597 14176
rect 13661 14112 13669 14176
rect 13349 13088 13669 14112
rect 13349 13024 13357 13088
rect 13421 13024 13437 13088
rect 13501 13024 13517 13088
rect 13581 13024 13597 13088
rect 13661 13024 13669 13088
rect 13349 12000 13669 13024
rect 13349 11936 13357 12000
rect 13421 11936 13437 12000
rect 13501 11936 13517 12000
rect 13581 11936 13597 12000
rect 13661 11936 13669 12000
rect 13349 10912 13669 11936
rect 13349 10848 13357 10912
rect 13421 10848 13437 10912
rect 13501 10848 13517 10912
rect 13581 10848 13597 10912
rect 13661 10848 13669 10912
rect 13349 9824 13669 10848
rect 13349 9760 13357 9824
rect 13421 9760 13437 9824
rect 13501 9760 13517 9824
rect 13581 9760 13597 9824
rect 13661 9760 13669 9824
rect 13349 8736 13669 9760
rect 13349 8672 13357 8736
rect 13421 8672 13437 8736
rect 13501 8672 13517 8736
rect 13581 8672 13597 8736
rect 13661 8672 13669 8736
rect 13349 7648 13669 8672
rect 13349 7584 13357 7648
rect 13421 7584 13437 7648
rect 13501 7584 13517 7648
rect 13581 7584 13597 7648
rect 13661 7584 13669 7648
rect 13349 6560 13669 7584
rect 13349 6496 13357 6560
rect 13421 6496 13437 6560
rect 13501 6496 13517 6560
rect 13581 6496 13597 6560
rect 13661 6496 13669 6560
rect 13349 5472 13669 6496
rect 13349 5408 13357 5472
rect 13421 5408 13437 5472
rect 13501 5408 13517 5472
rect 13581 5408 13597 5472
rect 13661 5408 13669 5472
rect 13349 4384 13669 5408
rect 13349 4320 13357 4384
rect 13421 4320 13437 4384
rect 13501 4320 13517 4384
rect 13581 4320 13597 4384
rect 13661 4320 13669 4384
rect 13349 3296 13669 4320
rect 13349 3232 13357 3296
rect 13421 3232 13437 3296
rect 13501 3232 13517 3296
rect 13581 3232 13597 3296
rect 13661 3232 13669 3296
rect 13349 2208 13669 3232
rect 13349 2144 13357 2208
rect 13421 2144 13437 2208
rect 13501 2144 13517 2208
rect 13581 2144 13597 2208
rect 13661 2144 13669 2208
rect 13349 1120 13669 2144
rect 13349 1056 13357 1120
rect 13421 1056 13437 1120
rect 13501 1056 13517 1120
rect 13581 1056 13597 1120
rect 13661 1056 13669 1120
rect 13349 496 13669 1056
rect 15200 14720 15520 15280
rect 15200 14656 15208 14720
rect 15272 14656 15288 14720
rect 15352 14656 15368 14720
rect 15432 14656 15448 14720
rect 15512 14656 15520 14720
rect 15200 13632 15520 14656
rect 15200 13568 15208 13632
rect 15272 13568 15288 13632
rect 15352 13568 15368 13632
rect 15432 13568 15448 13632
rect 15512 13568 15520 13632
rect 15200 12544 15520 13568
rect 15200 12480 15208 12544
rect 15272 12480 15288 12544
rect 15352 12480 15368 12544
rect 15432 12480 15448 12544
rect 15512 12480 15520 12544
rect 15200 11456 15520 12480
rect 15200 11392 15208 11456
rect 15272 11392 15288 11456
rect 15352 11392 15368 11456
rect 15432 11392 15448 11456
rect 15512 11392 15520 11456
rect 15200 10368 15520 11392
rect 15200 10304 15208 10368
rect 15272 10304 15288 10368
rect 15352 10304 15368 10368
rect 15432 10304 15448 10368
rect 15512 10304 15520 10368
rect 15200 9280 15520 10304
rect 15200 9216 15208 9280
rect 15272 9216 15288 9280
rect 15352 9216 15368 9280
rect 15432 9216 15448 9280
rect 15512 9216 15520 9280
rect 15200 8192 15520 9216
rect 15200 8128 15208 8192
rect 15272 8128 15288 8192
rect 15352 8128 15368 8192
rect 15432 8128 15448 8192
rect 15512 8128 15520 8192
rect 15200 7104 15520 8128
rect 15200 7040 15208 7104
rect 15272 7040 15288 7104
rect 15352 7040 15368 7104
rect 15432 7040 15448 7104
rect 15512 7040 15520 7104
rect 15200 6016 15520 7040
rect 15200 5952 15208 6016
rect 15272 5952 15288 6016
rect 15352 5952 15368 6016
rect 15432 5952 15448 6016
rect 15512 5952 15520 6016
rect 15200 4928 15520 5952
rect 15200 4864 15208 4928
rect 15272 4864 15288 4928
rect 15352 4864 15368 4928
rect 15432 4864 15448 4928
rect 15512 4864 15520 4928
rect 15200 3840 15520 4864
rect 15200 3776 15208 3840
rect 15272 3776 15288 3840
rect 15352 3776 15368 3840
rect 15432 3776 15448 3840
rect 15512 3776 15520 3840
rect 15200 2752 15520 3776
rect 15200 2688 15208 2752
rect 15272 2688 15288 2752
rect 15352 2688 15368 2752
rect 15432 2688 15448 2752
rect 15512 2688 15520 2752
rect 15200 1664 15520 2688
rect 15200 1600 15208 1664
rect 15272 1600 15288 1664
rect 15352 1600 15368 1664
rect 15432 1600 15448 1664
rect 15512 1600 15520 1664
rect 15200 576 15520 1600
rect 15200 512 15208 576
rect 15272 512 15288 576
rect 15352 512 15368 576
rect 15432 512 15448 576
rect 15512 512 15520 576
rect 15200 496 15520 512
use sky130_fd_sc_hd__a221o_1  _163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13340 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _166_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13432 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12328 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12604 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13156 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _172_
timestamp 1688980957
transform -1 0 12328 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _173_
timestamp 1688980957
transform 1 0 12328 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _174_
timestamp 1688980957
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _175_
timestamp 1688980957
transform -1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12788 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11316 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12788 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _179_
timestamp 1688980957
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _180_
timestamp 1688980957
transform -1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12236 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _182_
timestamp 1688980957
transform 1 0 11868 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _183_
timestamp 1688980957
transform 1 0 12236 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _184_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12972 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _186_
timestamp 1688980957
transform 1 0 10580 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10856 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _188_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10948 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _191_
timestamp 1688980957
transform -1 0 10488 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _192_
timestamp 1688980957
transform -1 0 10856 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _193_
timestamp 1688980957
transform -1 0 13432 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13524 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11592 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _196_
timestamp 1688980957
transform 1 0 11684 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10948 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _198_
timestamp 1688980957
transform -1 0 10396 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp 1688980957
transform 1 0 11684 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _200_
timestamp 1688980957
transform 1 0 10120 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _201_
timestamp 1688980957
transform -1 0 8648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _202_
timestamp 1688980957
transform -1 0 8280 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _203_
timestamp 1688980957
transform -1 0 9568 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _204_
timestamp 1688980957
transform 1 0 7636 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9016 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _206_
timestamp 1688980957
transform 1 0 8924 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8280 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _208_
timestamp 1688980957
transform 1 0 6900 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _209_
timestamp 1688980957
transform -1 0 6072 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _210_
timestamp 1688980957
transform 1 0 6532 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8188 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6900 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _213_
timestamp 1688980957
transform -1 0 7544 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _214_
timestamp 1688980957
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _215_
timestamp 1688980957
transform 1 0 7636 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _216_
timestamp 1688980957
transform -1 0 8648 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _217_
timestamp 1688980957
transform 1 0 7268 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1688980957
transform -1 0 6348 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _219_
timestamp 1688980957
transform 1 0 6164 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _220_
timestamp 1688980957
transform -1 0 6072 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _221_
timestamp 1688980957
transform 1 0 7728 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _222_
timestamp 1688980957
transform -1 0 7728 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _223_
timestamp 1688980957
transform 1 0 8372 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _224_
timestamp 1688980957
transform 1 0 8188 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9200 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1688980957
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _227_
timestamp 1688980957
transform -1 0 7452 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _228_
timestamp 1688980957
transform -1 0 6992 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _229_
timestamp 1688980957
transform 1 0 5796 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _230_
timestamp 1688980957
transform 1 0 4600 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _231_
timestamp 1688980957
transform 1 0 5336 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _232_
timestamp 1688980957
transform 1 0 6440 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _234_
timestamp 1688980957
transform 1 0 4968 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _235_
timestamp 1688980957
transform -1 0 6256 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _236_
timestamp 1688980957
transform 1 0 6716 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _237_
timestamp 1688980957
transform -1 0 7636 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _238_
timestamp 1688980957
transform 1 0 5980 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _239_
timestamp 1688980957
transform -1 0 5520 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _240_
timestamp 1688980957
transform 1 0 7820 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _241_
timestamp 1688980957
transform 1 0 7544 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _242_
timestamp 1688980957
transform 1 0 9108 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _243_
timestamp 1688980957
transform -1 0 9108 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _244_
timestamp 1688980957
transform 1 0 9016 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _245_
timestamp 1688980957
transform -1 0 9752 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _246_
timestamp 1688980957
transform 1 0 7084 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _247_
timestamp 1688980957
transform -1 0 8004 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _248_
timestamp 1688980957
transform 1 0 6716 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _249_
timestamp 1688980957
transform -1 0 5428 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _250_
timestamp 1688980957
transform -1 0 10120 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _251_
timestamp 1688980957
transform 1 0 8372 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _252_
timestamp 1688980957
transform -1 0 9016 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _253_
timestamp 1688980957
transform -1 0 9752 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1688980957
transform -1 0 10672 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _255_
timestamp 1688980957
transform -1 0 10396 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1688980957
transform 1 0 14352 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _258_
timestamp 1688980957
transform -1 0 5520 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _259_
timestamp 1688980957
transform -1 0 11684 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _260_
timestamp 1688980957
transform -1 0 11316 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10672 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _262_
timestamp 1688980957
transform -1 0 11040 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _263_
timestamp 1688980957
transform 1 0 10120 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _264_
timestamp 1688980957
transform -1 0 9016 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _265_
timestamp 1688980957
transform 1 0 8556 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _266_
timestamp 1688980957
transform 1 0 7636 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _267_
timestamp 1688980957
transform 1 0 8372 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _268_
timestamp 1688980957
transform -1 0 7912 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _269_
timestamp 1688980957
transform 1 0 6348 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1688980957
transform 1 0 7176 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7176 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _272_
timestamp 1688980957
transform -1 0 6532 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _273_
timestamp 1688980957
transform -1 0 5244 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _274_
timestamp 1688980957
transform 1 0 4324 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _275_
timestamp 1688980957
transform -1 0 4876 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _276_
timestamp 1688980957
transform 1 0 3864 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1688980957
transform 1 0 7544 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8464 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9476 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _280_
timestamp 1688980957
transform 1 0 8464 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _281_
timestamp 1688980957
transform -1 0 9292 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1688980957
transform 1 0 6716 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8464 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _284_
timestamp 1688980957
transform 1 0 4508 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _285_
timestamp 1688980957
transform 1 0 3772 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _286_
timestamp 1688980957
transform 1 0 4324 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _287_
timestamp 1688980957
transform 1 0 4876 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1688980957
transform -1 0 7820 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _289_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7544 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _290_
timestamp 1688980957
transform 1 0 6256 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _291_
timestamp 1688980957
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _292_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1688980957
transform -1 0 7544 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _294_
timestamp 1688980957
transform 1 0 6440 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1688980957
transform -1 0 6624 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _296_
timestamp 1688980957
transform 1 0 3772 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _297_
timestamp 1688980957
transform -1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6440 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _299_
timestamp 1688980957
transform 1 0 7084 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _300_
timestamp 1688980957
transform 1 0 8372 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _301_
timestamp 1688980957
transform 1 0 11132 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _302_
timestamp 1688980957
transform 1 0 12512 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _303_
timestamp 1688980957
transform -1 0 12512 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1688980957
transform 1 0 14536 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _305_
timestamp 1688980957
transform 1 0 12972 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _306_
timestamp 1688980957
transform 1 0 13524 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _307_
timestamp 1688980957
transform 1 0 7360 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _308_
timestamp 1688980957
transform 1 0 9108 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _309_
timestamp 1688980957
transform -1 0 12788 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _310_
timestamp 1688980957
transform 1 0 12052 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11408 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _312_
timestamp 1688980957
transform 1 0 12144 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _313_
timestamp 1688980957
transform -1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _314_
timestamp 1688980957
transform -1 0 12788 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _315_
timestamp 1688980957
transform 1 0 11224 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _316_
timestamp 1688980957
transform 1 0 10764 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _317_
timestamp 1688980957
transform -1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _318_
timestamp 1688980957
transform -1 0 12420 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _319_
timestamp 1688980957
transform -1 0 12052 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _320_
timestamp 1688980957
transform -1 0 11592 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _321_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _322_
timestamp 1688980957
transform 1 0 12696 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _323_
timestamp 1688980957
transform -1 0 13432 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _324_
timestamp 1688980957
transform 1 0 12328 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9016 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _326_
timestamp 1688980957
transform -1 0 12420 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _327_
timestamp 1688980957
transform -1 0 9568 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _328_
timestamp 1688980957
transform -1 0 8648 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _329_
timestamp 1688980957
transform -1 0 7268 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _330_
timestamp 1688980957
transform 1 0 5244 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _331_
timestamp 1688980957
transform -1 0 5152 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _332_
timestamp 1688980957
transform -1 0 4692 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _333_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _334_
timestamp 1688980957
transform 1 0 12788 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _335_
timestamp 1688980957
transform 1 0 13340 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _336_
timestamp 1688980957
transform 1 0 13340 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _337_
timestamp 1688980957
transform 1 0 13340 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _338_
timestamp 1688980957
transform 1 0 13340 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _339_
timestamp 1688980957
transform 1 0 13340 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _340_
timestamp 1688980957
transform 1 0 13340 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _341_
timestamp 1688980957
transform 1 0 10948 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _342_
timestamp 1688980957
transform 1 0 9936 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _343_
timestamp 1688980957
transform 1 0 11960 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _344_
timestamp 1688980957
transform 1 0 8648 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _345_
timestamp 1688980957
transform -1 0 9844 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _346_
timestamp 1688980957
transform 1 0 5428 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _347_
timestamp 1688980957
transform 1 0 4232 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _348_
timestamp 1688980957
transform 1 0 4232 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _349_
timestamp 1688980957
transform -1 0 10120 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _350_
timestamp 1688980957
transform 1 0 4140 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _351_
timestamp 1688980957
transform -1 0 4968 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _352_
timestamp 1688980957
transform -1 0 5244 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _353_
timestamp 1688980957
transform -1 0 10856 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _354_
timestamp 1688980957
transform 1 0 4876 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _355_
timestamp 1688980957
transform -1 0 10764 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _356_
timestamp 1688980957
transform 1 0 9660 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _357__12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12788 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _357_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10304 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1688980957
transform -1 0 7636 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1688980957
transform 1 0 10948 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1688980957
transform -1 0 7084 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1688980957
transform 1 0 10396 0 1 10336
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1688980957
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14628 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_157
timestamp 1688980957
transform 1 0 14996 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_149 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14260 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_157
timestamp 1688980957
transform 1 0 14996 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_153
timestamp 1688980957
transform 1 0 14628 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_157
timestamp 1688980957
transform 1 0 14996 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_60
timestamp 1688980957
transform 1 0 6072 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_72
timestamp 1688980957
transform 1 0 7176 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_84
timestamp 1688980957
transform 1 0 8280 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_96
timestamp 1688980957
transform 1 0 9384 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_104
timestamp 1688980957
transform 1 0 10120 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_108
timestamp 1688980957
transform 1 0 10488 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14260 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_157
timestamp 1688980957
transform 1 0 14996 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_101
timestamp 1688980957
transform 1 0 9844 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_118
timestamp 1688980957
transform 1 0 11408 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_130
timestamp 1688980957
transform 1 0 12512 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_153
timestamp 1688980957
transform 1 0 14628 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_157
timestamp 1688980957
transform 1 0 14996 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_69
timestamp 1688980957
transform 1 0 6900 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_80
timestamp 1688980957
transform 1 0 7912 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_121
timestamp 1688980957
transform 1 0 11684 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_133
timestamp 1688980957
transform 1 0 12788 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_145
timestamp 1688980957
transform 1 0 13892 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_157
timestamp 1688980957
transform 1 0 14996 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3220 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_37
timestamp 1688980957
transform 1 0 3956 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_56
timestamp 1688980957
transform 1 0 5704 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_68
timestamp 1688980957
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_76
timestamp 1688980957
transform 1 0 7544 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8372 0 1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_98
timestamp 1688980957
transform 1 0 9568 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_110
timestamp 1688980957
transform 1 0 10672 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_118
timestamp 1688980957
transform 1 0 11408 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_124
timestamp 1688980957
transform 1 0 11960 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_136
timestamp 1688980957
transform 1 0 13064 0 1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_153
timestamp 1688980957
transform 1 0 14628 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_157
timestamp 1688980957
transform 1 0 14996 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 1688980957
transform 1 0 5796 0 -1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_88
timestamp 1688980957
transform 1 0 8648 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_100
timestamp 1688980957
transform 1 0 9752 0 -1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_140
timestamp 1688980957
transform 1 0 13432 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_152
timestamp 1688980957
transform 1 0 14536 0 -1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5428 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_71
timestamp 1688980957
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_80
timestamp 1688980957
transform 1 0 7912 0 1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_144
timestamp 1688980957
transform 1 0 13800 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_156
timestamp 1688980957
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4140 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_77
timestamp 1688980957
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_83
timestamp 1688980957
transform 1 0 8188 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_95
timestamp 1688980957
transform 1 0 9292 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_107
timestamp 1688980957
transform 1 0 10396 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_152
timestamp 1688980957
transform 1 0 14536 0 -1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3220 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_37
timestamp 1688980957
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_55
timestamp 1688980957
transform 1 0 5612 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_61
timestamp 1688980957
transform 1 0 6164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_65
timestamp 1688980957
transform 1 0 6532 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_71
timestamp 1688980957
transform 1 0 7084 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 1688980957
transform 1 0 7912 0 1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_94
timestamp 1688980957
transform 1 0 9200 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_106
timestamp 1688980957
transform 1 0 10304 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_113
timestamp 1688980957
transform 1 0 10948 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_125
timestamp 1688980957
transform 1 0 12052 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_145
timestamp 1688980957
transform 1 0 13892 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_157
timestamp 1688980957
transform 1 0 14996 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4140 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_43
timestamp 1688980957
transform 1 0 4508 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_47
timestamp 1688980957
transform 1 0 4876 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_104
timestamp 1688980957
transform 1 0 10120 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_133
timestamp 1688980957
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_65
timestamp 1688980957
transform 1 0 6532 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_73
timestamp 1688980957
transform 1 0 7268 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 1688980957
transform 1 0 8004 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_99
timestamp 1688980957
transform 1 0 9660 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_111
timestamp 1688980957
transform 1 0 10764 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_125
timestamp 1688980957
transform 1 0 12052 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 12788 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_153
timestamp 1688980957
transform 1 0 14628 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_157
timestamp 1688980957
transform 1 0 14996 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3036 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_31
timestamp 1688980957
transform 1 0 3404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_74
timestamp 1688980957
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_86
timestamp 1688980957
transform 1 0 8464 0 -1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_100
timestamp 1688980957
transform 1 0 9752 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_113
timestamp 1688980957
transform 1 0 10948 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_117
timestamp 1688980957
transform 1 0 11316 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_128
timestamp 1688980957
transform 1 0 12328 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_136
timestamp 1688980957
transform 1 0 13064 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_51
timestamp 1688980957
transform 1 0 5244 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_57
timestamp 1688980957
transform 1 0 5796 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_62
timestamp 1688980957
transform 1 0 6256 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_70
timestamp 1688980957
transform 1 0 6992 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_112
timestamp 1688980957
transform 1 0 10856 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_118
timestamp 1688980957
transform 1 0 11408 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_123
timestamp 1688980957
transform 1 0 11868 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_129
timestamp 1688980957
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_149
timestamp 1688980957
transform 1 0 14260 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3036 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1688980957
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_57
timestamp 1688980957
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_70
timestamp 1688980957
transform 1 0 6992 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_75
timestamp 1688980957
transform 1 0 7452 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_79
timestamp 1688980957
transform 1 0 7820 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_85
timestamp 1688980957
transform 1 0 8372 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_106
timestamp 1688980957
transform 1 0 10304 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12052 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_133
timestamp 1688980957
transform 1 0 12788 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4324 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_63
timestamp 1688980957
transform 1 0 6348 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_75
timestamp 1688980957
transform 1 0 7452 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1688980957
transform 1 0 8004 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_90
timestamp 1688980957
transform 1 0 8832 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_94
timestamp 1688980957
transform 1 0 9200 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_114
timestamp 1688980957
transform 1 0 11040 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_119
timestamp 1688980957
transform 1 0 11500 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_127
timestamp 1688980957
transform 1 0 12236 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_149
timestamp 1688980957
transform 1 0 14260 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_157
timestamp 1688980957
transform 1 0 14996 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4140 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_47
timestamp 1688980957
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1688980957
transform 1 0 5428 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_66
timestamp 1688980957
transform 1 0 6624 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_72
timestamp 1688980957
transform 1 0 7176 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_79
timestamp 1688980957
transform 1 0 7820 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_85
timestamp 1688980957
transform 1 0 8372 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_104
timestamp 1688980957
transform 1 0 10120 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_113
timestamp 1688980957
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_122
timestamp 1688980957
transform 1 0 11776 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_126
timestamp 1688980957
transform 1 0 12144 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_49
timestamp 1688980957
transform 1 0 5060 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_71
timestamp 1688980957
transform 1 0 7084 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_97
timestamp 1688980957
transform 1 0 9476 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_127
timestamp 1688980957
transform 1 0 12236 0 1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_153
timestamp 1688980957
transform 1 0 14628 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_157
timestamp 1688980957
transform 1 0 14996 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3036 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1688980957
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_80
timestamp 1688980957
transform 1 0 7912 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_92
timestamp 1688980957
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_98
timestamp 1688980957
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp 1688980957
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_113
timestamp 1688980957
transform 1 0 10948 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_136
timestamp 1688980957
transform 1 0 13064 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3220 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_42
timestamp 1688980957
transform 1 0 4416 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_48
timestamp 1688980957
transform 1 0 4968 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_57
timestamp 1688980957
transform 1 0 5796 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_61
timestamp 1688980957
transform 1 0 6164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_95
timestamp 1688980957
transform 1 0 9292 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_123
timestamp 1688980957
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_128
timestamp 1688980957
transform 1 0 12328 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1688980957
transform 1 0 13156 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_149
timestamp 1688980957
transform 1 0 14260 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_157
timestamp 1688980957
transform 1 0 14996 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4140 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_47
timestamp 1688980957
transform 1 0 4876 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_69
timestamp 1688980957
transform 1 0 6900 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_77
timestamp 1688980957
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_92
timestamp 1688980957
transform 1 0 9016 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_96
timestamp 1688980957
transform 1 0 9384 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_103
timestamp 1688980957
transform 1 0 10028 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 10948 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_132
timestamp 1688980957
transform 1 0 12696 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_138
timestamp 1688980957
transform 1 0 13248 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_45
timestamp 1688980957
transform 1 0 4692 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_75
timestamp 1688980957
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_93
timestamp 1688980957
transform 1 0 9108 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_101
timestamp 1688980957
transform 1 0 9844 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_138
timestamp 1688980957
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_149
timestamp 1688980957
transform 1 0 14260 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_157
timestamp 1688980957
transform 1 0 14996 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3036 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_35
timestamp 1688980957
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_44
timestamp 1688980957
transform 1 0 4600 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_65
timestamp 1688980957
transform 1 0 6532 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_71
timestamp 1688980957
transform 1 0 7084 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_88
timestamp 1688980957
transform 1 0 8648 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_108
timestamp 1688980957
transform 1 0 10488 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_113
timestamp 1688980957
transform 1 0 10948 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_127
timestamp 1688980957
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_133
timestamp 1688980957
transform 1 0 12788 0 -1 13600
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_49
timestamp 1688980957
transform 1 0 5060 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_61
timestamp 1688980957
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_71
timestamp 1688980957
transform 1 0 7084 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_95
timestamp 1688980957
transform 1 0 9292 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_114
timestamp 1688980957
transform 1 0 11040 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_121
timestamp 1688980957
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_129
timestamp 1688980957
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_135
timestamp 1688980957
transform 1 0 12972 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_141
timestamp 1688980957
transform 1 0 13524 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_155
timestamp 1688980957
transform 1 0 14812 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3036 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_33
timestamp 1688980957
transform 1 0 3588 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp 1688980957
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_80
timestamp 1688980957
transform 1 0 7912 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_98
timestamp 1688980957
transform 1 0 9568 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_153
timestamp 1688980957
transform 1 0 14628 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_157
timestamp 1688980957
transform 1 0 14996 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_3
timestamp 1688980957
transform 1 0 828 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_8
timestamp 1688980957
transform 1 0 1288 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_16
timestamp 1688980957
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_22
timestamp 1688980957
transform 1 0 2576 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3220 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_35
timestamp 1688980957
transform 1 0 3772 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_43
timestamp 1688980957
transform 1 0 4508 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_54
timestamp 1688980957
transform 1 0 5520 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_57
timestamp 1688980957
transform 1 0 5796 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_63
timestamp 1688980957
transform 1 0 6348 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_71
timestamp 1688980957
transform 1 0 7084 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1688980957
transform 1 0 7636 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_95
timestamp 1688980957
transform 1 0 9292 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_101
timestamp 1688980957
transform 1 0 9844 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_105
timestamp 1688980957
transform 1 0 10212 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_111
timestamp 1688980957
transform 1 0 10764 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_113
timestamp 1688980957
transform 1 0 10948 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_119
timestamp 1688980957
transform 1 0 11500 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_127
timestamp 1688980957
transform 1 0 12236 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_136
timestamp 1688980957
transform 1 0 13064 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_141
timestamp 1688980957
transform 1 0 13524 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_147
timestamp 1688980957
transform 1 0 14076 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_155
timestamp 1688980957
transform 1 0 14812 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 9016 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 4508 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 12328 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 7084 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 12052 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 11868 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 15088 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 14536 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12788 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 11224 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 9936 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 9016 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 7360 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 6072 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 5244 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform 1 0 3496 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2208 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1688980957
transform 1 0 920 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 14076 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 15364 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 15364 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 15364 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 15364 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 15364 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 15364 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 15364 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 15364 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 15364 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 15364 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 15364 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 15364 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 15364 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 15364 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 15364 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 15364 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 15364 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 15364 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 15364 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 15364 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 15364 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 15364 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 15364 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 15364 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 15364 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 15364 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 15364 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 5704 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 10856 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 13432 0 1 14688
box -38 -48 130 592
<< labels >>
flabel metal4 s 4094 496 4414 15280 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7796 496 8116 15280 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11498 496 11818 15280 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15200 496 15520 15280 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2243 496 2563 15280 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5945 496 6265 15280 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9647 496 9967 15280 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13349 496 13669 15280 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 15014 15600 15070 16000 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal2 s 12438 15600 12494 16000 0 FreeSans 224 90 0 0 data[0]
port 3 nsew signal input
flabel metal2 s 11150 15600 11206 16000 0 FreeSans 224 90 0 0 data[1]
port 4 nsew signal input
flabel metal2 s 9862 15600 9918 16000 0 FreeSans 224 90 0 0 data[2]
port 5 nsew signal input
flabel metal2 s 8574 15600 8630 16000 0 FreeSans 224 90 0 0 data[3]
port 6 nsew signal input
flabel metal2 s 7286 15600 7342 16000 0 FreeSans 224 90 0 0 data[4]
port 7 nsew signal input
flabel metal2 s 5998 15600 6054 16000 0 FreeSans 224 90 0 0 data[5]
port 8 nsew signal input
flabel metal2 s 4710 15600 4766 16000 0 FreeSans 224 90 0 0 data[6]
port 9 nsew signal input
flabel metal2 s 3422 15600 3478 16000 0 FreeSans 224 90 0 0 data[7]
port 10 nsew signal input
flabel metal2 s 2134 15600 2190 16000 0 FreeSans 224 90 0 0 ext_data
port 11 nsew signal input
flabel metal2 s 846 15600 902 16000 0 FreeSans 224 90 0 0 load_divider
port 12 nsew signal input
flabel metal2 s 13726 15600 13782 16000 0 FreeSans 224 90 0 0 n_rst
port 13 nsew signal input
flabel metal3 s 15600 1096 16000 1216 0 FreeSans 480 0 0 0 r2r_out[0]
port 14 nsew signal tristate
flabel metal3 s 15600 3000 16000 3120 0 FreeSans 480 0 0 0 r2r_out[1]
port 15 nsew signal tristate
flabel metal3 s 15600 4904 16000 5024 0 FreeSans 480 0 0 0 r2r_out[2]
port 16 nsew signal tristate
flabel metal3 s 15600 6808 16000 6928 0 FreeSans 480 0 0 0 r2r_out[3]
port 17 nsew signal tristate
flabel metal3 s 15600 8712 16000 8832 0 FreeSans 480 0 0 0 r2r_out[4]
port 18 nsew signal tristate
flabel metal3 s 15600 10616 16000 10736 0 FreeSans 480 0 0 0 r2r_out[5]
port 19 nsew signal tristate
flabel metal3 s 15600 12520 16000 12640 0 FreeSans 480 0 0 0 r2r_out[6]
port 20 nsew signal tristate
flabel metal3 s 15600 14424 16000 14544 0 FreeSans 480 0 0 0 r2r_out[7]
port 21 nsew signal tristate
rlabel via1 8036 14688 8036 14688 0 VGND
rlabel metal1 7958 15232 7958 15232 0 VPWR
rlabel metal1 14168 14382 14168 14382 0 _000_
rlabel metal1 9660 12954 9660 12954 0 _001_
rlabel metal1 11458 14450 11458 14450 0 _002_
rlabel metal2 9246 14246 9246 14246 0 _003_
rlabel metal1 8878 12954 8878 12954 0 _004_
rlabel metal1 6992 14042 6992 14042 0 _005_
rlabel metal1 5699 12750 5699 12750 0 _006_
rlabel metal2 5014 14246 5014 14246 0 _007_
rlabel metal1 4472 12750 4472 12750 0 _008_
rlabel metal1 13708 6766 13708 6766 0 _009_
rlabel metal1 13064 5678 13064 5678 0 _010_
rlabel metal2 13662 8092 13662 8092 0 _011_
rlabel metal2 13662 9180 13662 9180 0 _012_
rlabel metal1 13570 10030 13570 10030 0 _013_
rlabel metal2 13662 11356 13662 11356 0 _014_
rlabel metal2 13662 12444 13662 12444 0 _015_
rlabel metal1 13294 13294 13294 13294 0 _016_
rlabel metal1 10994 6936 10994 6936 0 _017_
rlabel metal2 10350 2754 10350 2754 0 _018_
rlabel metal1 11776 4250 11776 4250 0 _019_
rlabel metal1 8724 5066 8724 5066 0 _020_
rlabel metal1 9250 2958 9250 2958 0 _021_
rlabel metal2 5934 2754 5934 2754 0 _022_
rlabel metal1 4917 4046 4917 4046 0 _023_
rlabel metal1 5796 5338 5796 5338 0 _024_
rlabel metal1 9338 6426 9338 6426 0 _025_
rlabel via1 4457 6154 4457 6154 0 _026_
rlabel metal1 4891 7990 4891 7990 0 _027_
rlabel metal1 5244 8942 5244 8942 0 _028_
rlabel metal2 9706 8194 9706 8194 0 _029_
rlabel via1 5193 9486 5193 9486 0 _030_
rlabel metal1 10308 9486 10308 9486 0 _031_
rlabel metal2 9706 11458 9706 11458 0 _032_
rlabel metal2 9246 11866 9246 11866 0 _033_
rlabel metal1 8188 11322 8188 11322 0 _034_
rlabel via1 7020 11662 7020 11662 0 _035_
rlabel metal1 8142 11186 8142 11186 0 _036_
rlabel metal1 5106 10778 5106 10778 0 _037_
rlabel metal1 5474 11696 5474 11696 0 _038_
rlabel metal1 5106 11322 5106 11322 0 _039_
rlabel metal1 5474 11084 5474 11084 0 _040_
rlabel metal1 7866 11628 7866 11628 0 _041_
rlabel metal1 7544 11050 7544 11050 0 _042_
rlabel metal1 6394 11526 6394 11526 0 _043_
rlabel metal1 7452 11186 7452 11186 0 _044_
rlabel metal1 7268 8398 7268 8398 0 _045_
rlabel metal1 7222 10234 7222 10234 0 _046_
rlabel metal1 6302 11050 6302 11050 0 _047_
rlabel metal1 5290 11628 5290 11628 0 _048_
rlabel metal1 4462 11322 4462 11322 0 _049_
rlabel metal1 5842 11186 5842 11186 0 _050_
rlabel metal1 6762 8398 6762 8398 0 _051_
rlabel metal1 7636 5746 7636 5746 0 _052_
rlabel metal1 10074 10064 10074 10064 0 _053_
rlabel metal1 8372 8398 8372 8398 0 _054_
rlabel metal1 12558 7242 12558 7242 0 _055_
rlabel metal2 13110 7140 13110 7140 0 _056_
rlabel metal2 9062 7276 9062 7276 0 _057_
rlabel metal1 13386 6222 13386 6222 0 _058_
rlabel metal2 8694 8398 8694 8398 0 _059_
rlabel metal1 10350 6766 10350 6766 0 _060_
rlabel metal2 12558 6426 12558 6426 0 _061_
rlabel metal1 11914 7990 11914 7990 0 _062_
rlabel via1 12185 6222 12185 6222 0 _063_
rlabel metal1 12466 6290 12466 6290 0 _064_
rlabel metal1 5336 9010 5336 9010 0 _065_
rlabel metal1 6711 4046 6711 4046 0 _066_
rlabel metal2 10994 9180 10994 9180 0 _067_
rlabel metal2 11822 8704 11822 8704 0 _068_
rlabel metal2 12006 8806 12006 8806 0 _069_
rlabel metal1 11500 9010 11500 9010 0 _070_
rlabel metal1 12742 8398 12742 8398 0 _071_
rlabel metal1 13386 9452 13386 9452 0 _072_
rlabel metal1 13294 9690 13294 9690 0 _073_
rlabel metal1 12696 9078 12696 9078 0 _074_
rlabel metal1 14030 9554 14030 9554 0 _075_
rlabel metal1 12926 10030 12926 10030 0 _076_
rlabel metal1 13248 10778 13248 10778 0 _077_
rlabel metal2 10672 5372 10672 5372 0 _078_
rlabel metal1 12374 10982 12374 10982 0 _079_
rlabel metal2 12650 10982 12650 10982 0 _080_
rlabel metal1 12006 12784 12006 12784 0 _081_
rlabel via1 12466 11186 12466 11186 0 _082_
rlabel metal1 13524 11322 13524 11322 0 _083_
rlabel metal1 12236 12274 12236 12274 0 _084_
rlabel metal1 12880 12750 12880 12750 0 _085_
rlabel metal1 12098 12716 12098 12716 0 _086_
rlabel metal1 14030 12784 14030 12784 0 _087_
rlabel metal1 12144 13362 12144 13362 0 _088_
rlabel metal1 12052 13498 12052 13498 0 _089_
rlabel metal1 12374 13770 12374 13770 0 _090_
rlabel metal1 12604 12410 12604 12410 0 _091_
rlabel metal1 12696 13498 12696 13498 0 _092_
rlabel metal2 10626 6630 10626 6630 0 _093_
rlabel metal1 8372 3366 8372 3366 0 _094_
rlabel metal1 11454 3570 11454 3570 0 _095_
rlabel metal1 10718 2482 10718 2482 0 _096_
rlabel metal1 10672 4794 10672 4794 0 _097_
rlabel metal1 12006 5236 12006 5236 0 _098_
rlabel metal1 12282 5100 12282 5100 0 _099_
rlabel metal1 11730 4080 11730 4080 0 _100_
rlabel metal2 10442 4845 10442 4845 0 _101_
rlabel metal1 10534 4522 10534 4522 0 _102_
rlabel metal2 10810 4828 10810 4828 0 _103_
rlabel metal1 9384 5134 9384 5134 0 _104_
rlabel metal1 8648 3706 8648 3706 0 _105_
rlabel metal2 9430 3740 9430 3740 0 _106_
rlabel metal1 8418 3638 8418 3638 0 _107_
rlabel metal1 9430 3706 9430 3706 0 _108_
rlabel metal1 7590 3026 7590 3026 0 _109_
rlabel metal1 6486 2482 6486 2482 0 _110_
rlabel metal2 6302 4488 6302 4488 0 _111_
rlabel metal1 7222 4692 7222 4692 0 _112_
rlabel metal1 7222 4250 7222 4250 0 _113_
rlabel metal1 5566 4556 5566 4556 0 _114_
rlabel metal1 6946 4522 6946 4522 0 _115_
rlabel metal1 7958 4794 7958 4794 0 _116_
rlabel metal1 7590 5066 7590 5066 0 _117_
rlabel metal1 6854 4692 6854 4692 0 _118_
rlabel metal1 6118 4794 6118 4794 0 _119_
rlabel metal1 8234 6970 8234 6970 0 _120_
rlabel metal1 7912 6902 7912 6902 0 _121_
rlabel metal1 8418 6902 8418 6902 0 _122_
rlabel metal1 8786 6222 8786 6222 0 _123_
rlabel metal1 6532 6834 6532 6834 0 _124_
rlabel metal1 6256 6698 6256 6698 0 _125_
rlabel metal1 6210 6868 6210 6868 0 _126_
rlabel metal1 4646 6800 4646 6800 0 _127_
rlabel metal1 5336 7990 5336 7990 0 _128_
rlabel metal1 6302 7888 6302 7888 0 _129_
rlabel metal1 5290 7888 5290 7888 0 _130_
rlabel metal2 6302 8738 6302 8738 0 _131_
rlabel metal1 7774 7344 7774 7344 0 _132_
rlabel metal1 7866 8296 7866 8296 0 _133_
rlabel metal1 5566 8976 5566 8976 0 _134_
rlabel metal1 8786 8296 8786 8296 0 _135_
rlabel metal2 9154 7956 9154 7956 0 _136_
rlabel metal1 8878 8364 8878 8364 0 _137_
rlabel metal1 9154 7922 9154 7922 0 _138_
rlabel metal1 9476 7922 9476 7922 0 _139_
rlabel metal1 7084 8874 7084 8874 0 _140_
rlabel metal1 9798 10132 9798 10132 0 _141_
rlabel metal1 6302 9690 6302 9690 0 _142_
rlabel metal2 10074 10472 10074 10472 0 _143_
rlabel metal1 8648 9622 8648 9622 0 _144_
rlabel metal1 9246 10064 9246 10064 0 _145_
rlabel metal1 9890 11220 9890 11220 0 _146_
rlabel metal1 10258 10778 10258 10778 0 _147_
rlabel metal1 4646 13838 4646 13838 0 _148_
rlabel metal1 5336 4658 5336 4658 0 _149_
rlabel metal1 10672 12614 10672 12614 0 _150_
rlabel metal1 10304 14042 10304 14042 0 _151_
rlabel metal1 8510 13906 8510 13906 0 _152_
rlabel metal1 8326 12614 8326 12614 0 _153_
rlabel metal1 6854 13906 6854 13906 0 _154_
rlabel metal2 7314 12206 7314 12206 0 _155_
rlabel metal1 6624 12954 6624 12954 0 _156_
rlabel metal1 4508 13906 4508 13906 0 _157_
rlabel metal2 4324 12852 4324 12852 0 _158_
rlabel metal2 8142 11951 8142 11951 0 _159_
rlabel metal2 8970 11458 8970 11458 0 _160_
rlabel viali 9153 11662 9153 11662 0 _161_
rlabel metal1 10258 9112 10258 9112 0 clk
rlabel metal1 9292 5814 9292 5814 0 clknet_0_clk
rlabel metal1 4278 5610 4278 5610 0 clknet_2_0__leaf_clk
rlabel metal1 10994 2958 10994 2958 0 clknet_2_1__leaf_clk
rlabel metal1 5106 14484 5106 14484 0 clknet_2_2__leaf_clk
rlabel metal1 9614 11730 9614 11730 0 clknet_2_3__leaf_clk
rlabel metal1 11224 4114 11224 4114 0 counter\[0\]
rlabel metal2 4554 8228 4554 8228 0 counter\[10\]
rlabel metal1 6210 8432 6210 8432 0 counter\[11\]
rlabel metal1 9384 8398 9384 8398 0 counter\[12\]
rlabel metal2 6302 10608 6302 10608 0 counter\[13\]
rlabel metal1 4462 10642 4462 10642 0 counter\[14\]
rlabel metal1 3910 11186 3910 11186 0 counter\[15\]
rlabel metal1 11132 4046 11132 4046 0 counter\[1\]
rlabel metal2 12374 4964 12374 4964 0 counter\[2\]
rlabel metal1 10120 4658 10120 4658 0 counter\[3\]
rlabel metal1 8096 4726 8096 4726 0 counter\[4\]
rlabel metal1 8188 4658 8188 4658 0 counter\[5\]
rlabel metal1 8372 4590 8372 4590 0 counter\[6\]
rlabel metal2 6946 5372 6946 5372 0 counter\[7\]
rlabel via1 8891 7310 8891 7310 0 counter\[8\]
rlabel metal1 8602 11186 8602 11186 0 counter\[9\]
rlabel metal1 12604 14926 12604 14926 0 data[0]
rlabel metal1 11224 14926 11224 14926 0 data[1]
rlabel metal1 10028 14926 10028 14926 0 data[2]
rlabel metal1 9062 14960 9062 14960 0 data[3]
rlabel metal1 7360 14926 7360 14926 0 data[4]
rlabel metal1 5980 14926 5980 14926 0 data[5]
rlabel metal1 5290 14892 5290 14892 0 data[6]
rlabel metal1 3496 14926 3496 14926 0 data[7]
rlabel metal2 10442 12648 10442 12648 0 divider\[0\]
rlabel metal2 8786 11560 8786 11560 0 divider\[1\]
rlabel metal1 8556 14586 8556 14586 0 divider\[2\]
rlabel metal1 7682 12784 7682 12784 0 divider\[3\]
rlabel metal1 7866 14518 7866 14518 0 divider\[4\]
rlabel metal1 6808 11798 6808 11798 0 divider\[5\]
rlabel metal1 5198 14960 5198 14960 0 divider\[6\]
rlabel metal1 3588 11730 3588 11730 0 divider\[7\]
rlabel metal1 2254 14926 2254 14926 0 ext_data
rlabel metal1 966 14926 966 14926 0 load_divider
rlabel metal1 13800 14926 13800 14926 0 n_rst
rlabel metal1 10166 12682 10166 12682 0 net1
rlabel metal1 4830 14926 4830 14926 0 net10
rlabel metal1 14214 14450 14214 14450 0 net11
rlabel metal1 12788 14518 12788 14518 0 net12
rlabel metal1 6532 4046 6532 4046 0 net13
rlabel metal1 8280 3570 8280 3570 0 net14
rlabel metal2 5382 8092 5382 8092 0 net15
rlabel metal1 11592 4658 11592 4658 0 net16
rlabel metal1 13570 5168 13570 5168 0 net17
rlabel metal1 6348 5134 6348 5134 0 net18
rlabel metal1 10442 6834 10442 6834 0 net19
rlabel metal1 11592 7854 11592 7854 0 net2
rlabel metal2 11178 11356 11178 11356 0 net20
rlabel metal1 14306 8398 14306 8398 0 net21
rlabel metal1 12788 13294 12788 13294 0 net22
rlabel metal1 10488 14790 10488 14790 0 net3
rlabel metal1 8970 12750 8970 12750 0 net4
rlabel metal1 7866 13838 7866 13838 0 net5
rlabel viali 6026 13290 6026 13290 0 net6
rlabel metal1 4830 13804 4830 13804 0 net7
rlabel metal1 4278 13260 4278 13260 0 net8
rlabel metal1 6578 10166 6578 10166 0 net9
rlabel metal3 15372 1156 15372 1156 0 r2r_out[0]
rlabel metal3 15096 3060 15096 3060 0 r2r_out[1]
rlabel metal1 12650 8330 12650 8330 0 r2r_out[2]
rlabel metal1 14996 8806 14996 8806 0 r2r_out[3]
rlabel metal1 15042 9894 15042 9894 0 r2r_out[4]
rlabel metal3 15418 10676 15418 10676 0 r2r_out[5]
rlabel metal1 15088 12342 15088 12342 0 r2r_out[6]
rlabel metal1 15042 13498 15042 13498 0 r2r_out[7]
rlabel metal1 4922 14008 4922 14008 0 rst
<< properties >>
string FIXED_BBOX 0 0 16000 16000
<< end >>
