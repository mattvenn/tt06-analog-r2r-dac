* NGSPICE file created from r2r_parax.ext - technology: sky130A

.subckt r2r_parax b0 b1 b2 b3 b4 b5 b6 b7 out GND
X0 a_766_6998# a_1366_2566# a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=20
X1 b0.t0 a_n1834_10998# a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=40
X2 b6.t0 a_1966_6998# a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=40
X3 b3.t0 a_166_2566# a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=40
X4 b5.t0 a_1366_2566# a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=40
X5 a_n1834_10998# a_n1034_2566# a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=20
X6 a_n1834_10998# GND.t0 a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=40
X7 b1.t0 a_n1034_2566# a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=40
X8 a_1966_6998# out.t0 a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=20
X9 a_766_6998# a_166_2566# a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=20
X10 a_1966_6998# a_1366_2566# a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=20
X11 b2.t0 a_n434_6998# a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=40
X12 b4.t0 a_766_6998# a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=40
X13 a_n434_6998# a_n1034_2566# a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=20
X14 b7.t0 out.t1 a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=40
X15 a_n434_6998# a_166_2566# a_n1964_2436# sky130_fd_pr__res_high_po_0p35 l=20
R0 b0 b0.t0 43.7238
R1 b6 b6.t0 43.7238
R2 b3 b3.t0 43.7238
R3 b5 b5.t0 43.7238
R4 GND GND.t0 43.6798
R5 b1 b1.t0 43.7238
R6 out.n0 out.t0 50.8673
R7 out.n0 out.t1 43.5548
R8 out out.n0 2.05675
R9 b2 b2.t0 43.7238
R10 b4 b4.t0 43.7238
R11 b7 b7.t0 43.7238
C0 a_166_2566# a_1366_2566# 0.182372f
C1 b0 b1 0.098267f
C2 a_n1834_10998# a_n434_6998# 1.8e-21
C3 b2 b1 0.098267f
C4 b5 b4 0.098267f
C5 b7 b6 0.098267f
C6 a_1966_6998# out 0.106769f
C7 a_n1834_10998# a_n1034_2566# 0.20932f
C8 a_n434_6998# a_n1034_2566# 0.131455f
C9 b5 b6 0.098267f
C10 a_1966_6998# a_1366_2566# 0.131485f
C11 a_n434_6998# a_166_2566# 0.209322f
C12 b3 b4 0.098267f
C13 a_766_6998# a_1366_2566# 0.209322f
C14 GND a_n1034_2566# 0.023658f
C15 out a_1366_2566# 0.151801f
C16 a_766_6998# a_166_2566# 0.131455f
C17 b3 b2 0.098267f
C18 a_n1034_2566# a_166_2566# 0.182372f
C19 out a_n1964_2436# 4.20278f
C20 b7 a_n1964_2436# 0.971435f
C21 b6 a_n1964_2436# 0.866417f
C22 b5 a_n1964_2436# 0.866417f
C23 b4 a_n1964_2436# 0.866417f
C24 b3 a_n1964_2436# 0.866417f
C25 b2 a_n1964_2436# 0.866417f
C26 b1 a_n1964_2436# 0.866417f
C27 b0 a_n1964_2436# 0.971438f
C28 GND a_n1964_2436# 0.991776f
C29 a_1966_6998# a_n1964_2436# 2.02255f
C30 a_1366_2566# a_n1964_2436# 3.90969f
C31 a_766_6998# a_n1964_2436# 1.95966f
C32 a_166_2566# a_n1964_2436# 3.87524f
C33 a_n434_6998# a_n1964_2436# 1.95966f
C34 a_n1034_2566# a_n1964_2436# 4.05843f
C35 a_n1834_10998# a_n1964_2436# 3.79668f
.ends

