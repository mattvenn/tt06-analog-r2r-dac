** sch_path: /home/matt/work/asic-workshop/shuttle-2404/tt06-analog-r2r-dac/xschem/r2r.sch
.subckt r2r b1 b0 b2 b3 b5 out b4 b6 b7
*.ipin b1
*.ipin b0
*.ipin b2
*.ipin b3
*.ipin b5
*.opin out
*.ipin b4
*.ipin b6
*.ipin b7
R1 b0 net1 1k m=1
R2 b1 net2 1k m=1
R3 b2 net3 1k m=1
R4 net1 GND 1k m=1
R5 b3 net4 1k m=1
R6 net2 net1 500 m=1
R7 net3 net2 500 m=1
R8 net4 net3 500 m=1
R9 b4 net5 1k m=1
R10 b5 net6 1k m=1
R11 b6 net7 1k m=1
R12 b7 out 1k m=1
R13 net6 net5 500 m=1
R14 net7 net6 500 m=1
R15 out net7 500 m=1
R16 net5 net4 500 m=1
.ends
.GLOBAL GND
.end
