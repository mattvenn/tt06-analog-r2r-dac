VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_mattvenn_r2r_dac
  CLASS BLOCK ;
  FOREIGN tt_um_mattvenn_r2r_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 8.440 5.520 9.940 221.280 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 18.090 204.925 92.530 206.530 ;
      LAYER pwell ;
        RECT 18.285 203.725 19.655 204.535 ;
        RECT 19.665 203.725 25.175 204.535 ;
        RECT 27.485 203.725 28.855 204.505 ;
        RECT 28.865 203.725 30.695 204.535 ;
        RECT 31.175 203.810 31.605 204.595 ;
        RECT 31.625 203.725 32.995 204.535 ;
        RECT 33.005 203.725 34.835 204.405 ;
        RECT 34.845 203.725 38.515 204.535 ;
        RECT 39.445 203.725 41.275 204.405 ;
        RECT 41.285 203.725 44.035 204.535 ;
        RECT 44.055 203.810 44.485 204.595 ;
        RECT 44.505 204.435 45.450 204.635 ;
        RECT 46.785 204.435 47.715 204.635 ;
        RECT 44.505 203.955 47.715 204.435 ;
        RECT 44.505 203.755 47.575 203.955 ;
        RECT 44.505 203.725 45.450 203.755 ;
        RECT 18.425 203.515 18.595 203.725 ;
        RECT 19.805 203.515 19.975 203.725 ;
        RECT 23.495 203.560 23.655 203.670 ;
        RECT 24.405 203.515 24.575 203.705 ;
        RECT 25.335 203.570 25.495 203.680 ;
        RECT 26.245 203.535 26.415 203.705 ;
        RECT 27.625 203.535 27.795 203.725 ;
        RECT 29.005 203.535 29.175 203.725 ;
        RECT 30.840 203.565 30.960 203.675 ;
        RECT 31.765 203.535 31.935 203.725 ;
        RECT 33.145 203.535 33.315 203.725 ;
        RECT 34.065 203.515 34.235 203.705 ;
        RECT 34.985 203.535 35.155 203.725 ;
        RECT 36.825 203.515 36.995 203.705 ;
        RECT 38.675 203.570 38.835 203.680 ;
        RECT 39.585 203.535 39.755 203.725 ;
        RECT 41.425 203.535 41.595 203.725 ;
        RECT 44.640 203.565 44.760 203.675 ;
        RECT 45.105 203.535 45.275 203.705 ;
        RECT 47.405 203.535 47.575 203.755 ;
        RECT 47.725 203.725 49.095 204.505 ;
        RECT 49.105 203.725 51.855 204.535 ;
        RECT 52.325 203.725 53.695 204.505 ;
        RECT 53.705 203.725 56.455 204.535 ;
        RECT 56.935 203.810 57.365 204.595 ;
        RECT 57.385 204.435 58.315 204.635 ;
        RECT 59.650 204.435 60.595 204.635 ;
        RECT 57.385 203.955 60.595 204.435 ;
        RECT 57.525 203.755 60.595 203.955 ;
        RECT 47.875 203.535 48.045 203.725 ;
        RECT 45.105 203.515 45.305 203.535 ;
        RECT 48.785 203.515 48.955 203.705 ;
        RECT 49.245 203.535 49.415 203.725 ;
        RECT 52.000 203.565 52.120 203.675 ;
        RECT 52.475 203.535 52.645 203.725 ;
        RECT 53.845 203.535 54.015 203.725 ;
        RECT 56.600 203.565 56.720 203.675 ;
        RECT 57.525 203.515 57.695 203.755 ;
        RECT 59.650 203.725 60.595 203.755 ;
        RECT 60.605 203.725 61.975 204.505 ;
        RECT 61.985 203.725 63.355 204.535 ;
        RECT 63.365 204.435 64.310 204.635 ;
        RECT 65.645 204.435 66.575 204.635 ;
        RECT 63.365 203.955 66.575 204.435 ;
        RECT 63.365 203.755 66.435 203.955 ;
        RECT 63.365 203.725 64.310 203.755 ;
        RECT 57.985 203.515 58.155 203.705 ;
        RECT 59.820 203.565 59.940 203.675 ;
        RECT 61.655 203.535 61.825 203.725 ;
        RECT 62.125 203.535 62.295 203.725 ;
        RECT 66.265 203.535 66.435 203.755 ;
        RECT 66.585 203.725 67.955 204.505 ;
        RECT 67.965 203.725 69.795 204.535 ;
        RECT 69.815 203.810 70.245 204.595 ;
        RECT 70.265 203.725 72.095 204.535 ;
        RECT 72.105 204.435 73.050 204.635 ;
        RECT 74.385 204.435 75.315 204.635 ;
        RECT 72.105 203.955 75.315 204.435 ;
        RECT 72.105 203.755 75.175 203.955 ;
        RECT 72.105 203.725 73.050 203.755 ;
        RECT 66.735 203.535 66.905 203.725 ;
        RECT 67.185 203.515 67.355 203.705 ;
        RECT 67.645 203.515 67.815 203.705 ;
        RECT 68.105 203.535 68.275 203.725 ;
        RECT 69.480 203.565 69.600 203.675 ;
        RECT 70.405 203.535 70.575 203.725 ;
        RECT 75.005 203.535 75.175 203.755 ;
        RECT 75.325 203.725 76.695 204.505 ;
        RECT 76.705 203.725 78.075 204.535 ;
        RECT 78.085 203.725 79.455 204.505 ;
        RECT 79.465 203.725 81.295 204.535 ;
        RECT 81.325 203.725 82.675 204.635 ;
        RECT 82.695 203.810 83.125 204.595 ;
        RECT 83.145 203.725 84.515 204.535 ;
        RECT 84.525 203.725 85.895 204.505 ;
        RECT 85.905 203.725 89.575 204.535 ;
        RECT 89.585 203.725 90.955 204.505 ;
        RECT 90.965 203.725 92.335 204.535 ;
        RECT 75.475 203.535 75.645 203.725 ;
        RECT 76.845 203.535 77.015 203.725 ;
        RECT 77.305 203.515 77.475 203.705 ;
        RECT 77.775 203.560 77.935 203.670 ;
        RECT 78.235 203.535 78.405 203.725 ;
        RECT 79.605 203.535 79.775 203.725 ;
        RECT 81.440 203.535 81.610 203.725 ;
        RECT 81.900 203.515 82.070 203.705 ;
        RECT 82.365 203.515 82.535 203.705 ;
        RECT 83.285 203.535 83.455 203.725 ;
        RECT 84.665 203.535 84.835 203.725 ;
        RECT 86.045 203.535 86.215 203.725 ;
        RECT 90.635 203.535 90.805 203.725 ;
        RECT 92.025 203.515 92.195 203.725 ;
        RECT 18.285 202.705 19.655 203.515 ;
        RECT 19.665 202.705 23.335 203.515 ;
        RECT 24.265 202.835 33.875 203.515 ;
        RECT 33.925 202.835 36.665 203.515 ;
        RECT 36.685 202.835 43.995 203.515 ;
        RECT 28.775 202.615 29.705 202.835 ;
        RECT 32.535 202.605 33.875 202.835 ;
        RECT 40.200 202.615 41.110 202.835 ;
        RECT 42.645 202.605 43.995 202.835 ;
        RECT 44.055 202.645 44.485 203.430 ;
        RECT 45.105 202.835 48.635 203.515 ;
        RECT 48.645 202.835 50.475 203.515 ;
        RECT 45.810 202.605 48.635 202.835 ;
        RECT 49.130 202.605 50.475 202.835 ;
        RECT 50.525 202.835 57.835 203.515 ;
        RECT 50.525 202.605 51.875 202.835 ;
        RECT 53.410 202.615 54.320 202.835 ;
        RECT 57.845 202.705 59.675 203.515 ;
        RECT 60.185 202.835 67.495 203.515 ;
        RECT 60.185 202.605 61.535 202.835 ;
        RECT 63.070 202.615 63.980 202.835 ;
        RECT 67.505 202.705 69.335 203.515 ;
        RECT 69.815 202.645 70.245 203.430 ;
        RECT 70.305 202.835 77.615 203.515 ;
        RECT 70.305 202.605 71.655 202.835 ;
        RECT 73.190 202.615 74.100 202.835 ;
        RECT 78.545 202.605 82.215 203.515 ;
        RECT 82.225 202.835 90.925 203.515 ;
        RECT 85.770 202.615 86.680 202.835 ;
        RECT 88.220 202.605 90.925 202.835 ;
        RECT 90.965 202.705 92.335 203.515 ;
      LAYER nwell ;
        RECT 18.090 199.485 92.530 202.315 ;
      LAYER pwell ;
        RECT 18.285 198.285 19.655 199.095 ;
        RECT 19.665 198.285 25.175 199.095 ;
        RECT 25.185 198.285 27.935 199.095 ;
        RECT 27.955 198.285 29.305 199.195 ;
        RECT 29.325 198.285 31.155 199.095 ;
        RECT 31.175 198.370 31.605 199.155 ;
        RECT 31.625 198.285 32.995 199.095 ;
        RECT 36.520 198.965 37.430 199.185 ;
        RECT 38.965 198.965 40.315 199.195 ;
        RECT 33.005 198.285 40.315 198.965 ;
        RECT 40.365 198.285 43.115 199.095 ;
        RECT 43.125 198.965 45.950 199.195 ;
        RECT 46.805 198.995 47.750 199.195 ;
        RECT 49.085 198.995 50.015 199.195 ;
        RECT 43.125 198.285 46.655 198.965 ;
        RECT 46.805 198.515 50.015 198.995 ;
        RECT 46.805 198.315 49.875 198.515 ;
        RECT 46.805 198.285 47.750 198.315 ;
        RECT 18.425 198.075 18.595 198.285 ;
        RECT 19.805 198.075 19.975 198.285 ;
        RECT 25.325 198.075 25.495 198.285 ;
        RECT 29.005 198.095 29.175 198.285 ;
        RECT 29.465 198.095 29.635 198.285 ;
        RECT 30.845 198.075 31.015 198.265 ;
        RECT 31.765 198.095 31.935 198.285 ;
        RECT 33.145 198.095 33.315 198.285 ;
        RECT 36.365 198.075 36.535 198.265 ;
        RECT 40.505 198.095 40.675 198.285 ;
        RECT 46.455 198.265 46.655 198.285 ;
        RECT 41.885 198.075 42.055 198.265 ;
        RECT 43.720 198.125 43.840 198.235 ;
        RECT 44.645 198.075 44.815 198.265 ;
        RECT 46.485 198.095 46.655 198.265 ;
        RECT 47.400 198.125 47.520 198.235 ;
        RECT 47.865 198.075 48.035 198.265 ;
        RECT 49.245 198.075 49.415 198.265 ;
        RECT 49.705 198.095 49.875 198.315 ;
        RECT 50.025 198.285 55.535 199.095 ;
        RECT 55.545 198.285 56.915 199.095 ;
        RECT 56.935 198.370 57.365 199.155 ;
        RECT 57.385 198.965 60.210 199.195 ;
        RECT 57.385 198.285 60.915 198.965 ;
        RECT 61.065 198.285 62.895 199.095 ;
        RECT 64.210 198.965 67.035 199.195 ;
        RECT 63.505 198.285 67.035 198.965 ;
        RECT 67.045 198.285 70.715 199.095 ;
        RECT 70.725 198.285 72.095 199.095 ;
        RECT 72.950 198.965 75.775 199.195 ;
        RECT 72.245 198.285 75.775 198.965 ;
        RECT 75.785 198.285 79.455 199.095 ;
        RECT 80.405 198.285 81.755 199.195 ;
        RECT 82.695 198.370 83.125 199.155 ;
        RECT 83.160 198.285 84.975 199.195 ;
        RECT 86.000 198.965 86.920 199.195 ;
        RECT 86.000 198.285 89.465 198.965 ;
        RECT 89.585 198.285 90.955 199.095 ;
        RECT 90.965 198.285 92.335 199.095 ;
        RECT 50.165 198.095 50.335 198.285 ;
        RECT 52.920 198.125 53.040 198.235 ;
        RECT 55.685 198.095 55.855 198.285 ;
        RECT 60.715 198.265 60.915 198.285 ;
        RECT 56.605 198.095 56.775 198.265 ;
        RECT 56.575 198.075 56.775 198.095 ;
        RECT 18.285 197.265 19.655 198.075 ;
        RECT 19.665 197.265 25.175 198.075 ;
        RECT 25.185 197.265 30.695 198.075 ;
        RECT 30.705 197.265 36.215 198.075 ;
        RECT 36.225 197.265 41.735 198.075 ;
        RECT 41.745 197.265 43.575 198.075 ;
        RECT 44.055 197.205 44.485 197.990 ;
        RECT 44.505 197.265 47.255 198.075 ;
        RECT 47.735 197.165 49.085 198.075 ;
        RECT 49.105 197.265 52.775 198.075 ;
        RECT 53.245 197.395 56.775 198.075 ;
        RECT 56.925 198.045 57.870 198.075 ;
        RECT 59.825 198.045 59.995 198.265 ;
        RECT 60.285 198.075 60.455 198.265 ;
        RECT 60.745 198.095 60.915 198.265 ;
        RECT 61.205 198.095 61.375 198.285 ;
        RECT 63.505 198.265 63.705 198.285 ;
        RECT 63.040 198.125 63.160 198.235 ;
        RECT 63.505 198.095 63.675 198.265 ;
        RECT 67.185 198.095 67.355 198.285 ;
        RECT 67.155 198.075 67.355 198.095 ;
        RECT 67.645 198.075 67.815 198.265 ;
        RECT 69.480 198.125 69.600 198.235 ;
        RECT 70.405 198.075 70.575 198.265 ;
        RECT 70.865 198.095 71.035 198.285 ;
        RECT 72.245 198.265 72.445 198.285 ;
        RECT 71.785 198.095 71.955 198.265 ;
        RECT 72.245 198.095 72.415 198.265 ;
        RECT 71.785 198.075 71.985 198.095 ;
        RECT 75.465 198.075 75.635 198.265 ;
        RECT 75.925 198.095 76.095 198.285 ;
        RECT 79.155 198.120 79.315 198.230 ;
        RECT 79.615 198.130 79.775 198.240 ;
        RECT 80.070 198.075 80.240 198.265 ;
        RECT 81.440 198.095 81.610 198.285 ;
        RECT 81.915 198.130 82.075 198.240 ;
        RECT 83.285 198.095 83.455 198.285 ;
        RECT 85.120 198.240 85.290 198.265 ;
        RECT 85.120 198.130 85.295 198.240 ;
        RECT 85.120 198.075 85.290 198.130 ;
        RECT 85.585 198.095 85.755 198.265 ;
        RECT 85.605 198.075 85.755 198.095 ;
        RECT 87.885 198.075 88.055 198.265 ;
        RECT 89.265 198.095 89.435 198.285 ;
        RECT 89.725 198.095 89.895 198.285 ;
        RECT 90.640 198.125 90.760 198.235 ;
        RECT 92.025 198.075 92.195 198.285 ;
        RECT 56.925 197.845 59.995 198.045 ;
        RECT 53.245 197.165 56.070 197.395 ;
        RECT 56.925 197.365 60.135 197.845 ;
        RECT 56.925 197.165 57.870 197.365 ;
        RECT 59.205 197.165 60.135 197.365 ;
        RECT 60.145 197.265 63.815 198.075 ;
        RECT 63.825 197.395 67.355 198.075 ;
        RECT 63.825 197.165 66.650 197.395 ;
        RECT 67.505 197.265 69.335 198.075 ;
        RECT 69.815 197.205 70.245 197.990 ;
        RECT 70.265 197.265 71.635 198.075 ;
        RECT 71.785 197.395 75.315 198.075 ;
        RECT 72.490 197.165 75.315 197.395 ;
        RECT 75.325 197.265 78.995 198.075 ;
        RECT 79.925 197.165 81.755 198.075 ;
        RECT 81.960 197.165 85.435 198.075 ;
        RECT 85.605 197.255 87.535 198.075 ;
        RECT 87.745 197.265 90.495 198.075 ;
        RECT 90.965 197.265 92.335 198.075 ;
        RECT 86.585 197.165 87.535 197.255 ;
      LAYER nwell ;
        RECT 18.090 194.045 92.530 196.875 ;
      LAYER pwell ;
        RECT 18.285 192.845 19.655 193.655 ;
        RECT 19.665 192.845 25.175 193.655 ;
        RECT 25.185 192.845 30.695 193.655 ;
        RECT 31.175 192.930 31.605 193.715 ;
        RECT 36.060 193.525 36.970 193.745 ;
        RECT 38.505 193.525 39.855 193.755 ;
        RECT 32.545 192.845 39.855 193.525 ;
        RECT 39.905 192.845 41.735 193.655 ;
        RECT 43.550 193.555 44.495 193.755 ;
        RECT 41.745 192.875 44.495 193.555 ;
        RECT 46.325 193.525 47.255 193.755 ;
        RECT 18.425 192.635 18.595 192.845 ;
        RECT 19.805 192.635 19.975 192.845 ;
        RECT 25.325 192.655 25.495 192.845 ;
        RECT 26.245 192.635 26.415 192.825 ;
        RECT 30.840 192.685 30.960 192.795 ;
        RECT 31.775 192.690 31.935 192.800 ;
        RECT 32.685 192.655 32.855 192.845 ;
        RECT 33.600 192.685 33.720 192.795 ;
        RECT 34.980 192.635 35.150 192.825 ;
        RECT 35.445 192.635 35.615 192.825 ;
        RECT 36.825 192.635 36.995 192.825 ;
        RECT 38.205 192.635 38.375 192.825 ;
        RECT 40.045 192.635 40.215 192.845 ;
        RECT 41.890 192.655 42.060 192.875 ;
        RECT 43.550 192.845 44.495 192.875 ;
        RECT 44.505 192.845 47.255 193.525 ;
        RECT 48.225 193.525 49.575 193.755 ;
        RECT 51.110 193.525 52.020 193.745 ;
        RECT 48.225 192.845 55.535 193.525 ;
        RECT 55.545 192.845 56.915 193.655 ;
        RECT 56.935 192.930 57.365 193.715 ;
        RECT 57.385 192.845 58.755 193.655 ;
        RECT 58.775 192.845 60.125 193.755 ;
        RECT 60.185 193.525 61.535 193.755 ;
        RECT 63.070 193.525 63.980 193.745 ;
        RECT 60.185 192.845 67.495 193.525 ;
        RECT 67.505 192.845 69.335 193.655 ;
        RECT 69.385 193.525 70.735 193.755 ;
        RECT 72.270 193.525 73.180 193.745 ;
        RECT 69.385 192.845 76.695 193.525 ;
        RECT 76.705 192.845 78.075 193.655 ;
        RECT 79.135 193.525 80.065 193.755 ;
        RECT 78.230 192.845 80.065 193.525 ;
        RECT 80.585 193.665 81.535 193.755 ;
        RECT 80.585 192.845 82.515 193.665 ;
        RECT 82.695 192.930 83.125 193.715 ;
        RECT 83.145 192.845 86.815 193.755 ;
        RECT 86.845 192.845 88.195 193.755 ;
        RECT 88.205 192.845 90.955 193.655 ;
        RECT 90.965 192.845 92.335 193.655 ;
        RECT 44.645 192.795 44.815 192.845 ;
        RECT 43.720 192.685 43.840 192.795 ;
        RECT 44.640 192.685 44.815 192.795 ;
        RECT 44.645 192.655 44.815 192.685 ;
        RECT 45.110 192.635 45.280 192.825 ;
        RECT 47.415 192.690 47.575 192.800 ;
        RECT 48.785 192.635 48.955 192.825 ;
        RECT 54.305 192.635 54.475 192.825 ;
        RECT 54.765 192.635 54.935 192.825 ;
        RECT 55.225 192.655 55.395 192.845 ;
        RECT 55.685 192.655 55.855 192.845 ;
        RECT 57.525 192.655 57.695 192.845 ;
        RECT 59.825 192.655 59.995 192.845 ;
        RECT 60.285 192.635 60.455 192.825 ;
        RECT 18.285 191.825 19.655 192.635 ;
        RECT 19.665 191.825 25.175 192.635 ;
        RECT 26.105 191.955 33.415 192.635 ;
        RECT 29.620 191.735 30.530 191.955 ;
        RECT 32.065 191.725 33.415 191.955 ;
        RECT 33.945 191.725 35.295 192.635 ;
        RECT 35.305 191.825 36.675 192.635 ;
        RECT 36.695 191.725 38.045 192.635 ;
        RECT 38.065 191.825 39.895 192.635 ;
        RECT 40.015 191.955 43.480 192.635 ;
        RECT 42.560 191.725 43.480 191.955 ;
        RECT 44.055 191.765 44.485 192.550 ;
        RECT 44.965 191.725 48.620 192.635 ;
        RECT 48.645 191.825 51.395 192.635 ;
        RECT 51.405 191.725 54.615 192.635 ;
        RECT 54.625 191.825 60.135 192.635 ;
        RECT 60.145 191.825 62.895 192.635 ;
        RECT 63.040 192.605 63.210 192.825 ;
        RECT 65.345 192.635 65.515 192.825 ;
        RECT 67.185 192.655 67.355 192.845 ;
        RECT 67.645 192.655 67.815 192.845 ;
        RECT 69.035 192.680 69.195 192.790 ;
        RECT 70.415 192.680 70.575 192.790 ;
        RECT 64.240 192.605 65.195 192.635 ;
        RECT 62.915 191.925 65.195 192.605 ;
        RECT 64.240 191.725 65.195 191.925 ;
        RECT 65.205 191.825 68.875 192.635 ;
        RECT 71.185 192.605 72.130 192.635 ;
        RECT 74.085 192.605 74.255 192.825 ;
        RECT 74.545 192.635 74.715 192.825 ;
        RECT 76.385 192.655 76.555 192.845 ;
        RECT 76.845 192.655 77.015 192.845 ;
        RECT 78.230 192.825 78.395 192.845 ;
        RECT 82.365 192.825 82.515 192.845 ;
        RECT 78.225 192.655 78.395 192.825 ;
        RECT 80.065 192.635 80.235 192.825 ;
        RECT 81.900 192.685 82.020 192.795 ;
        RECT 82.365 192.635 82.535 192.825 ;
        RECT 83.285 192.655 83.455 192.845 ;
        RECT 86.960 192.655 87.130 192.845 ;
        RECT 88.345 192.655 88.515 192.845 ;
        RECT 92.025 192.635 92.195 192.845 ;
        RECT 69.815 191.765 70.245 192.550 ;
        RECT 71.185 192.405 74.255 192.605 ;
        RECT 71.185 191.925 74.395 192.405 ;
        RECT 71.185 191.725 72.130 191.925 ;
        RECT 73.465 191.725 74.395 191.925 ;
        RECT 74.405 191.825 79.915 192.635 ;
        RECT 79.925 191.825 81.755 192.635 ;
        RECT 82.225 191.955 90.925 192.635 ;
        RECT 85.770 191.735 86.680 191.955 ;
        RECT 88.220 191.725 90.925 191.955 ;
        RECT 90.965 191.825 92.335 192.635 ;
      LAYER nwell ;
        RECT 18.090 188.605 92.530 191.435 ;
      LAYER pwell ;
        RECT 18.285 187.405 19.655 188.215 ;
        RECT 19.665 187.405 25.175 188.215 ;
        RECT 25.185 187.405 27.935 188.215 ;
        RECT 27.945 187.405 29.295 188.315 ;
        RECT 29.325 187.405 31.155 188.215 ;
        RECT 31.175 187.490 31.605 188.275 ;
        RECT 31.625 187.405 32.995 188.215 ;
        RECT 33.175 187.405 36.675 188.315 ;
        RECT 39.680 188.085 40.815 188.315 ;
        RECT 43.105 188.085 44.035 188.315 ;
        RECT 37.605 187.405 40.815 188.085 ;
        RECT 41.285 187.405 44.035 188.085 ;
        RECT 44.055 187.405 45.405 188.315 ;
        RECT 45.425 187.405 47.255 188.215 ;
        RECT 47.265 187.405 48.635 188.185 ;
        RECT 48.645 187.405 52.315 188.215 ;
        RECT 53.245 187.405 56.900 188.315 ;
        RECT 56.935 187.490 57.365 188.275 ;
        RECT 57.395 187.405 61.515 188.315 ;
        RECT 61.525 188.085 62.445 188.315 ;
        RECT 65.205 188.085 66.135 188.315 ;
        RECT 70.705 188.085 71.635 188.315 ;
        RECT 61.525 187.405 65.110 188.085 ;
        RECT 65.205 187.405 67.955 188.085 ;
        RECT 68.885 187.405 71.635 188.085 ;
        RECT 71.655 187.405 73.005 188.315 ;
        RECT 73.485 188.115 74.430 188.315 ;
        RECT 73.485 187.435 76.235 188.115 ;
        RECT 73.485 187.405 74.430 187.435 ;
        RECT 18.425 187.195 18.595 187.405 ;
        RECT 19.805 187.215 19.975 187.405 ;
        RECT 25.325 187.215 25.495 187.405 ;
        RECT 27.625 187.195 27.795 187.385 ;
        RECT 28.090 187.215 28.260 187.405 ;
        RECT 29.465 187.215 29.635 187.405 ;
        RECT 31.765 187.385 31.935 187.405 ;
        RECT 33.175 187.385 33.310 187.405 ;
        RECT 31.305 187.195 31.475 187.385 ;
        RECT 31.755 187.215 31.935 187.385 ;
        RECT 33.140 187.215 33.310 187.385 ;
        RECT 31.755 187.195 31.925 187.215 ;
        RECT 34.990 187.195 35.160 187.385 ;
        RECT 36.360 187.215 36.530 187.385 ;
        RECT 36.835 187.250 36.995 187.360 ;
        RECT 37.745 187.215 37.915 187.405 ;
        RECT 36.395 187.195 36.530 187.215 ;
        RECT 40.045 187.195 40.215 187.385 ;
        RECT 40.960 187.245 41.080 187.355 ;
        RECT 41.425 187.215 41.595 187.405 ;
        RECT 42.805 187.195 42.975 187.385 ;
        RECT 43.275 187.240 43.435 187.350 ;
        RECT 44.185 187.215 44.355 187.405 ;
        RECT 44.655 187.240 44.815 187.350 ;
        RECT 45.565 187.195 45.735 187.405 ;
        RECT 48.325 187.215 48.495 187.405 ;
        RECT 48.785 187.215 48.955 187.405 ;
        RECT 52.475 187.250 52.635 187.360 ;
        RECT 52.925 187.195 53.095 187.385 ;
        RECT 53.390 187.215 53.560 187.405 ;
        RECT 58.445 187.195 58.615 187.385 ;
        RECT 59.365 187.215 59.535 187.405 ;
        RECT 61.205 187.215 61.375 187.405 ;
        RECT 61.670 187.215 61.840 187.405 ;
        RECT 63.045 187.195 63.215 187.385 ;
        RECT 63.505 187.195 63.675 187.385 ;
        RECT 66.720 187.245 66.840 187.355 ;
        RECT 18.285 186.385 19.655 187.195 ;
        RECT 20.625 186.515 27.935 187.195 ;
        RECT 28.040 186.515 31.505 187.195 ;
        RECT 20.625 186.285 21.975 186.515 ;
        RECT 23.510 186.295 24.420 186.515 ;
        RECT 28.040 186.285 28.960 186.515 ;
        RECT 31.625 186.285 34.835 187.195 ;
        RECT 34.845 186.285 36.195 187.195 ;
        RECT 36.395 186.285 39.895 187.195 ;
        RECT 39.920 186.285 41.735 187.195 ;
        RECT 41.755 186.285 43.105 187.195 ;
        RECT 44.055 186.325 44.485 187.110 ;
        RECT 45.425 186.515 52.735 187.195 ;
        RECT 48.940 186.295 49.850 186.515 ;
        RECT 51.385 186.285 52.735 186.515 ;
        RECT 52.785 186.385 58.295 187.195 ;
        RECT 58.305 186.385 60.135 187.195 ;
        RECT 60.145 186.285 63.355 187.195 ;
        RECT 63.445 186.285 66.445 187.195 ;
        RECT 67.190 187.165 67.360 187.385 ;
        RECT 67.645 187.215 67.815 187.405 ;
        RECT 68.115 187.250 68.275 187.360 ;
        RECT 69.025 187.215 69.195 187.405 ;
        RECT 72.705 187.215 72.875 187.405 ;
        RECT 73.165 187.355 73.335 187.385 ;
        RECT 73.160 187.245 73.335 187.355 ;
        RECT 68.850 187.165 69.795 187.195 ;
        RECT 67.045 186.485 69.795 187.165 ;
        RECT 70.265 187.165 71.210 187.195 ;
        RECT 73.165 187.165 73.335 187.245 ;
        RECT 75.920 187.215 76.090 187.435 ;
        RECT 76.245 187.405 81.755 188.215 ;
        RECT 82.695 187.490 83.125 188.275 ;
        RECT 83.145 187.405 88.655 188.215 ;
        RECT 88.665 187.405 90.495 188.215 ;
        RECT 90.965 187.405 92.335 188.215 ;
        RECT 76.385 187.195 76.555 187.405 ;
        RECT 76.840 187.245 76.960 187.355 ;
        RECT 78.220 187.195 78.390 187.385 ;
        RECT 78.690 187.195 78.860 187.385 ;
        RECT 81.915 187.250 82.075 187.360 ;
        RECT 82.365 187.195 82.535 187.385 ;
        RECT 83.285 187.215 83.455 187.405 ;
        RECT 88.805 187.215 88.975 187.405 ;
        RECT 90.640 187.245 90.760 187.355 ;
        RECT 92.025 187.195 92.195 187.405 ;
        RECT 68.850 186.285 69.795 186.485 ;
        RECT 69.815 186.325 70.245 187.110 ;
        RECT 70.265 186.965 73.335 187.165 ;
        RECT 70.265 186.485 73.475 186.965 ;
        RECT 70.265 186.285 71.210 186.485 ;
        RECT 72.545 186.285 73.475 186.485 ;
        RECT 73.485 186.285 76.655 187.195 ;
        RECT 77.185 186.285 78.535 187.195 ;
        RECT 78.545 186.285 82.200 187.195 ;
        RECT 82.225 186.515 90.925 187.195 ;
        RECT 85.770 186.295 86.680 186.515 ;
        RECT 88.220 186.285 90.925 186.515 ;
        RECT 90.965 186.385 92.335 187.195 ;
      LAYER nwell ;
        RECT 18.090 183.165 92.530 185.995 ;
      LAYER pwell ;
        RECT 18.285 181.965 19.655 182.775 ;
        RECT 19.665 181.965 25.175 182.775 ;
        RECT 25.185 181.965 27.015 182.775 ;
        RECT 27.040 181.965 28.855 182.875 ;
        RECT 28.885 181.965 30.235 182.875 ;
        RECT 31.175 182.050 31.605 182.835 ;
        RECT 41.025 182.785 41.975 182.875 ;
        RECT 31.710 181.965 40.815 182.645 ;
        RECT 41.025 181.965 42.955 182.785 ;
        RECT 44.175 182.645 45.105 182.875 ;
        RECT 46.565 182.785 47.515 182.875 ;
        RECT 18.425 181.755 18.595 181.965 ;
        RECT 19.805 181.755 19.975 181.965 ;
        RECT 25.325 181.755 25.495 181.965 ;
        RECT 27.165 181.775 27.335 181.965 ;
        RECT 29.000 181.775 29.170 181.965 ;
        RECT 30.395 181.810 30.555 181.920 ;
        RECT 30.845 181.755 31.015 181.945 ;
        RECT 36.375 181.800 36.535 181.910 ;
        RECT 39.125 181.755 39.295 181.945 ;
        RECT 39.585 181.755 39.755 181.945 ;
        RECT 40.505 181.775 40.675 181.965 ;
        RECT 42.805 181.945 42.955 181.965 ;
        RECT 43.270 181.965 45.105 182.645 ;
        RECT 45.585 181.965 47.515 182.785 ;
        RECT 47.725 181.965 51.395 182.875 ;
        RECT 51.405 181.965 55.075 182.775 ;
        RECT 55.555 181.965 56.905 182.875 ;
        RECT 56.935 182.050 57.365 182.835 ;
        RECT 57.385 181.965 66.490 182.645 ;
        RECT 66.585 181.965 67.955 182.775 ;
        RECT 67.965 181.965 71.440 182.875 ;
        RECT 71.645 181.965 74.385 182.645 ;
        RECT 74.405 181.965 79.915 182.775 ;
        RECT 79.935 181.965 82.665 182.875 ;
        RECT 82.695 182.050 83.125 182.835 ;
        RECT 83.145 181.965 86.620 182.875 ;
        RECT 86.825 182.645 87.745 182.875 ;
        RECT 86.825 181.965 89.115 182.645 ;
        RECT 89.125 181.965 90.955 182.775 ;
        RECT 90.965 181.965 92.335 182.775 ;
        RECT 43.270 181.945 43.435 181.965 ;
        RECT 45.585 181.945 45.735 181.965 ;
        RECT 41.420 181.805 41.540 181.915 ;
        RECT 42.805 181.775 42.980 181.945 ;
        RECT 43.265 181.775 43.435 181.945 ;
        RECT 42.810 181.755 42.980 181.775 ;
        RECT 44.645 181.755 44.815 181.945 ;
        RECT 45.565 181.775 45.735 181.945 ;
        RECT 47.870 181.775 48.040 181.965 ;
        RECT 50.165 181.755 50.335 181.945 ;
        RECT 51.545 181.775 51.715 181.965 ;
        RECT 55.220 181.805 55.340 181.915 ;
        RECT 55.685 181.755 55.855 181.945 ;
        RECT 56.605 181.775 56.775 181.965 ;
        RECT 57.525 181.775 57.695 181.965 ;
        RECT 60.285 181.775 60.455 181.945 ;
        RECT 60.285 181.755 60.435 181.775 ;
        RECT 61.670 181.755 61.840 181.945 ;
        RECT 62.125 181.755 62.295 181.945 ;
        RECT 64.885 181.755 65.055 181.945 ;
        RECT 66.725 181.775 66.895 181.965 ;
        RECT 68.110 181.775 68.280 181.965 ;
        RECT 68.565 181.755 68.735 181.945 ;
        RECT 70.415 181.800 70.575 181.910 ;
        RECT 71.785 181.775 71.955 181.965 ;
        RECT 74.080 181.755 74.250 181.945 ;
        RECT 74.545 181.755 74.715 181.965 ;
        RECT 80.065 181.755 80.235 181.965 ;
        RECT 83.290 181.775 83.460 181.965 ;
        RECT 85.585 181.755 85.755 181.945 ;
        RECT 88.805 181.775 88.975 181.965 ;
        RECT 89.265 181.775 89.435 181.965 ;
        RECT 92.025 181.755 92.195 181.965 ;
        RECT 18.285 180.945 19.655 181.755 ;
        RECT 19.665 180.945 25.175 181.755 ;
        RECT 25.185 180.945 30.695 181.755 ;
        RECT 30.705 180.945 36.215 181.755 ;
        RECT 37.145 181.075 39.435 181.755 ;
        RECT 37.145 180.845 38.065 181.075 ;
        RECT 39.445 180.945 41.275 181.755 ;
        RECT 41.745 180.845 43.095 181.755 ;
        RECT 44.055 180.885 44.485 181.670 ;
        RECT 44.505 180.945 50.015 181.755 ;
        RECT 50.025 180.945 55.535 181.755 ;
        RECT 55.545 180.945 58.295 181.755 ;
        RECT 58.505 180.935 60.435 181.755 ;
        RECT 58.505 180.845 59.455 180.935 ;
        RECT 60.605 180.845 61.955 181.755 ;
        RECT 61.985 181.075 64.725 181.755 ;
        RECT 64.745 180.945 68.415 181.755 ;
        RECT 68.425 180.945 69.795 181.755 ;
        RECT 69.815 180.885 70.245 181.670 ;
        RECT 71.475 180.845 74.395 181.755 ;
        RECT 74.405 180.945 79.915 181.755 ;
        RECT 79.925 180.945 85.435 181.755 ;
        RECT 85.445 180.945 90.955 181.755 ;
        RECT 90.965 180.945 92.335 181.755 ;
      LAYER nwell ;
        RECT 18.090 177.725 92.530 180.555 ;
      LAYER pwell ;
        RECT 18.285 176.525 19.655 177.335 ;
        RECT 19.665 176.525 23.335 177.335 ;
        RECT 27.320 177.205 28.230 177.425 ;
        RECT 29.765 177.205 31.115 177.435 ;
        RECT 23.805 176.525 31.115 177.205 ;
        RECT 31.175 176.610 31.605 177.395 ;
        RECT 31.795 176.525 35.295 177.435 ;
        RECT 37.960 177.205 38.880 177.435 ;
        RECT 40.355 177.205 41.275 177.435 ;
        RECT 42.885 177.345 43.835 177.435 ;
        RECT 35.415 176.525 38.880 177.205 ;
        RECT 38.985 176.525 41.275 177.205 ;
        RECT 41.905 176.525 43.835 177.345 ;
        RECT 44.530 177.205 45.875 177.435 ;
        RECT 44.045 176.525 45.875 177.205 ;
        RECT 46.805 176.525 48.175 177.305 ;
        RECT 49.105 176.525 52.775 177.435 ;
        RECT 53.095 177.205 54.025 177.435 ;
        RECT 53.095 176.525 54.930 177.205 ;
        RECT 55.085 176.525 56.435 177.435 ;
        RECT 56.935 176.610 57.365 177.395 ;
        RECT 58.755 177.205 59.675 177.435 ;
        RECT 61.055 177.205 61.975 177.435 ;
        RECT 57.385 176.525 59.675 177.205 ;
        RECT 59.685 176.525 61.975 177.205 ;
        RECT 61.985 176.525 64.725 177.205 ;
        RECT 64.745 176.525 68.415 177.335 ;
        RECT 69.355 176.525 70.705 177.435 ;
        RECT 74.240 177.205 75.150 177.425 ;
        RECT 76.685 177.205 78.035 177.435 ;
        RECT 70.725 176.525 78.035 177.205 ;
        RECT 78.180 177.205 79.100 177.435 ;
        RECT 78.180 176.525 81.645 177.205 ;
        RECT 82.695 176.610 83.125 177.395 ;
        RECT 83.145 177.205 84.075 177.435 ;
        RECT 83.145 176.525 87.045 177.205 ;
        RECT 87.305 176.525 88.655 177.435 ;
        RECT 88.665 176.525 90.495 177.335 ;
        RECT 90.965 176.525 92.335 177.335 ;
        RECT 18.425 176.315 18.595 176.525 ;
        RECT 19.805 176.315 19.975 176.525 ;
        RECT 23.480 176.365 23.600 176.475 ;
        RECT 23.945 176.335 24.115 176.525 ;
        RECT 31.795 176.505 31.930 176.525 ;
        RECT 28.545 176.315 28.715 176.505 ;
        RECT 29.005 176.315 29.175 176.505 ;
        RECT 31.760 176.335 31.940 176.505 ;
        RECT 31.770 176.315 31.940 176.335 ;
        RECT 33.145 176.315 33.315 176.505 ;
        RECT 35.445 176.335 35.615 176.525 ;
        RECT 35.900 176.315 36.070 176.505 ;
        RECT 36.365 176.315 36.535 176.505 ;
        RECT 39.125 176.475 39.295 176.525 ;
        RECT 41.905 176.505 42.055 176.525 ;
        RECT 39.120 176.365 39.295 176.475 ;
        RECT 39.125 176.335 39.295 176.365 ;
        RECT 39.585 176.315 39.755 176.505 ;
        RECT 40.965 176.315 41.135 176.505 ;
        RECT 41.420 176.365 41.540 176.475 ;
        RECT 41.885 176.335 42.055 176.505 ;
        RECT 43.720 176.365 43.840 176.475 ;
        RECT 44.185 176.335 44.355 176.525 ;
        RECT 44.645 176.315 44.815 176.505 ;
        RECT 46.035 176.370 46.195 176.480 ;
        RECT 47.865 176.335 48.035 176.525 ;
        RECT 48.335 176.370 48.495 176.480 ;
        RECT 49.250 176.335 49.420 176.525 ;
        RECT 54.765 176.505 54.930 176.525 ;
        RECT 52.005 176.315 52.175 176.505 ;
        RECT 54.765 176.335 54.935 176.505 ;
        RECT 56.150 176.335 56.320 176.525 ;
        RECT 56.600 176.365 56.720 176.475 ;
        RECT 57.525 176.335 57.695 176.525 ;
        RECT 59.825 176.335 59.995 176.525 ;
        RECT 62.125 176.335 62.295 176.525 ;
        RECT 63.505 176.315 63.675 176.505 ;
        RECT 64.885 176.335 65.055 176.525 ;
        RECT 67.180 176.315 67.350 176.505 ;
        RECT 67.645 176.315 67.815 176.505 ;
        RECT 68.575 176.370 68.735 176.480 ;
        RECT 69.480 176.365 69.600 176.475 ;
        RECT 70.405 176.335 70.575 176.525 ;
        RECT 70.865 176.335 71.035 176.525 ;
        RECT 73.625 176.315 73.795 176.505 ;
        RECT 74.080 176.315 74.250 176.505 ;
        RECT 77.760 176.365 77.880 176.475 ;
        RECT 78.225 176.335 78.395 176.505 ;
        RECT 81.445 176.335 81.615 176.525 ;
        RECT 81.915 176.370 82.075 176.480 ;
        RECT 78.235 176.315 78.395 176.335 ;
        RECT 82.365 176.315 82.535 176.505 ;
        RECT 83.560 176.335 83.730 176.525 ;
        RECT 87.420 176.335 87.590 176.525 ;
        RECT 88.805 176.335 88.975 176.525 ;
        RECT 90.640 176.365 90.760 176.475 ;
        RECT 92.025 176.315 92.195 176.525 ;
        RECT 18.285 175.505 19.655 176.315 ;
        RECT 19.665 175.505 25.175 176.315 ;
        RECT 25.280 175.635 28.745 176.315 ;
        RECT 25.280 175.405 26.200 175.635 ;
        RECT 28.865 175.505 31.615 176.315 ;
        RECT 31.625 175.405 32.975 176.315 ;
        RECT 33.005 175.505 34.835 176.315 ;
        RECT 34.865 175.405 36.215 176.315 ;
        RECT 36.225 175.505 38.975 176.315 ;
        RECT 39.455 175.405 40.805 176.315 ;
        RECT 40.825 175.505 43.575 176.315 ;
        RECT 44.055 175.445 44.485 176.230 ;
        RECT 44.505 175.635 51.815 176.315 ;
        RECT 51.865 175.635 60.970 176.315 ;
        RECT 48.020 175.415 48.930 175.635 ;
        RECT 50.465 175.405 51.815 175.635 ;
        RECT 61.075 175.405 63.805 176.315 ;
        RECT 64.020 175.405 67.495 176.315 ;
        RECT 67.520 175.405 69.335 176.315 ;
        RECT 69.815 175.445 70.245 176.230 ;
        RECT 70.360 175.635 73.825 176.315 ;
        RECT 70.360 175.405 71.280 175.635 ;
        RECT 73.955 175.405 77.615 176.315 ;
        RECT 78.235 175.405 81.890 176.315 ;
        RECT 82.225 175.635 90.925 176.315 ;
        RECT 85.770 175.415 86.680 175.635 ;
        RECT 88.220 175.405 90.925 175.635 ;
        RECT 90.965 175.505 92.335 176.315 ;
      LAYER nwell ;
        RECT 18.090 172.285 92.530 175.115 ;
      LAYER pwell ;
        RECT 18.285 171.085 19.655 171.895 ;
        RECT 19.665 171.085 22.415 171.895 ;
        RECT 26.400 171.765 27.310 171.985 ;
        RECT 28.845 171.765 30.195 171.995 ;
        RECT 22.885 171.085 30.195 171.765 ;
        RECT 31.175 171.170 31.605 171.955 ;
        RECT 31.640 171.085 33.455 171.995 ;
        RECT 33.465 171.085 35.295 171.895 ;
        RECT 35.305 171.795 36.250 171.995 ;
        RECT 37.585 171.795 38.515 171.995 ;
        RECT 35.305 171.315 38.515 171.795 ;
        RECT 40.600 171.765 41.735 171.995 ;
        RECT 43.150 171.765 44.495 171.995 ;
        RECT 47.005 171.905 47.955 171.995 ;
        RECT 35.305 171.115 38.375 171.315 ;
        RECT 35.305 171.085 36.250 171.115 ;
        RECT 18.425 170.875 18.595 171.085 ;
        RECT 19.805 170.875 19.975 171.085 ;
        RECT 22.560 170.925 22.680 171.035 ;
        RECT 23.025 170.895 23.195 171.085 ;
        RECT 25.325 170.875 25.495 171.065 ;
        RECT 27.160 170.875 27.330 171.065 ;
        RECT 30.395 170.930 30.555 171.040 ;
        RECT 31.765 170.895 31.935 171.085 ;
        RECT 33.605 170.895 33.775 171.085 ;
        RECT 37.285 170.875 37.455 171.065 ;
        RECT 38.205 170.895 38.375 171.115 ;
        RECT 38.525 171.085 41.735 171.765 ;
        RECT 42.665 171.085 44.495 171.765 ;
        RECT 44.505 171.085 46.335 171.895 ;
        RECT 47.005 171.085 48.935 171.905 ;
        RECT 49.105 171.085 54.615 171.895 ;
        RECT 54.625 171.085 56.455 171.895 ;
        RECT 56.935 171.170 57.365 171.955 ;
        RECT 57.555 171.085 61.055 171.995 ;
        RECT 61.065 171.085 62.880 171.995 ;
        RECT 62.915 171.085 64.265 171.995 ;
        RECT 68.260 171.765 69.170 171.985 ;
        RECT 70.705 171.765 72.055 171.995 ;
        RECT 64.745 171.085 72.055 171.765 ;
        RECT 72.105 171.085 77.615 171.895 ;
        RECT 77.625 171.085 81.295 171.895 ;
        RECT 81.305 171.085 82.655 171.995 ;
        RECT 82.695 171.170 83.125 171.955 ;
        RECT 83.145 171.085 84.495 171.995 ;
        RECT 84.525 171.085 90.035 171.895 ;
        RECT 90.965 171.085 92.335 171.895 ;
        RECT 38.665 170.895 38.835 171.085 ;
        RECT 40.500 170.875 40.670 171.065 ;
        RECT 40.965 170.875 41.135 171.065 ;
        RECT 41.895 170.930 42.055 171.040 ;
        RECT 42.805 170.895 42.975 171.085 ;
        RECT 43.720 170.925 43.840 171.035 ;
        RECT 44.645 170.875 44.815 171.085 ;
        RECT 48.785 171.065 48.935 171.085 ;
        RECT 46.480 170.925 46.600 171.035 ;
        RECT 48.785 170.895 48.955 171.065 ;
        RECT 49.245 170.895 49.415 171.085 ;
        RECT 50.165 170.875 50.335 171.065 ;
        RECT 52.000 170.925 52.120 171.035 ;
        RECT 52.465 170.875 52.635 171.065 ;
        RECT 54.765 170.895 54.935 171.085 ;
        RECT 57.555 171.065 57.690 171.085 ;
        RECT 56.600 170.925 56.720 171.035 ;
        RECT 57.520 170.895 57.690 171.065 ;
        RECT 59.820 170.875 59.990 171.065 ;
        RECT 61.205 170.875 61.375 171.065 ;
        RECT 62.585 170.895 62.755 171.085 ;
        RECT 63.965 170.895 64.135 171.085 ;
        RECT 64.420 170.925 64.540 171.035 ;
        RECT 64.885 170.895 65.055 171.085 ;
        RECT 66.725 170.875 66.895 171.065 ;
        RECT 69.480 170.925 69.600 171.035 ;
        RECT 70.405 170.875 70.575 171.065 ;
        RECT 72.245 170.895 72.415 171.085 ;
        RECT 74.080 170.925 74.200 171.035 ;
        RECT 77.300 170.875 77.470 171.065 ;
        RECT 77.765 170.895 77.935 171.085 ;
        RECT 18.285 170.065 19.655 170.875 ;
        RECT 19.665 170.065 25.175 170.875 ;
        RECT 25.185 170.065 27.015 170.875 ;
        RECT 27.045 169.965 28.395 170.875 ;
        RECT 28.490 170.195 37.595 170.875 ;
        RECT 37.895 169.965 40.815 170.875 ;
        RECT 40.825 170.065 43.575 170.875 ;
        RECT 44.055 170.005 44.485 170.790 ;
        RECT 44.505 170.065 50.015 170.875 ;
        RECT 50.025 170.065 51.855 170.875 ;
        RECT 52.325 170.195 59.635 170.875 ;
        RECT 55.840 169.975 56.750 170.195 ;
        RECT 58.285 169.965 59.635 170.195 ;
        RECT 59.705 169.965 61.055 170.875 ;
        RECT 61.065 170.065 66.575 170.875 ;
        RECT 66.585 170.065 69.335 170.875 ;
        RECT 69.815 170.005 70.245 170.790 ;
        RECT 70.265 170.065 73.935 170.875 ;
        RECT 74.695 169.965 77.615 170.875 ;
        RECT 77.625 170.845 78.580 170.875 ;
        RECT 79.610 170.845 79.780 171.065 ;
        RECT 80.070 170.875 80.240 171.065 ;
        RECT 81.450 170.895 81.620 171.085 ;
        RECT 83.290 170.895 83.460 171.085 ;
        RECT 83.745 170.875 83.915 171.065 ;
        RECT 84.665 170.895 84.835 171.085 ;
        RECT 89.265 170.875 89.435 171.065 ;
        RECT 90.195 170.930 90.355 171.040 ;
        RECT 92.025 170.875 92.195 171.085 ;
        RECT 77.625 170.165 79.905 170.845 ;
        RECT 77.625 169.965 78.580 170.165 ;
        RECT 79.925 169.965 83.580 170.875 ;
        RECT 83.605 170.065 89.115 170.875 ;
        RECT 89.125 170.065 90.955 170.875 ;
        RECT 90.965 170.065 92.335 170.875 ;
      LAYER nwell ;
        RECT 18.090 166.845 92.530 169.675 ;
      LAYER pwell ;
        RECT 18.285 165.645 19.655 166.455 ;
        RECT 19.665 165.645 25.175 166.455 ;
        RECT 25.185 165.645 30.695 166.455 ;
        RECT 31.175 165.730 31.605 166.515 ;
        RECT 31.625 165.645 34.375 166.455 ;
        RECT 36.460 166.325 37.595 166.555 ;
        RECT 38.745 166.465 39.695 166.555 ;
        RECT 34.385 165.645 37.595 166.325 ;
        RECT 37.765 165.645 39.695 166.465 ;
        RECT 43.880 166.325 44.790 166.545 ;
        RECT 46.325 166.325 47.675 166.555 ;
        RECT 40.365 165.645 47.675 166.325 ;
        RECT 47.725 165.645 49.555 166.455 ;
        RECT 52.220 166.325 53.140 166.555 ;
        RECT 49.675 165.645 53.140 166.325 ;
        RECT 53.725 165.645 55.075 166.555 ;
        RECT 55.095 165.645 56.445 166.555 ;
        RECT 56.935 165.730 57.365 166.515 ;
        RECT 57.385 165.645 61.055 166.455 ;
        RECT 61.065 165.645 62.435 166.455 ;
        RECT 62.445 165.645 64.260 166.555 ;
        RECT 64.285 165.645 66.115 166.555 ;
        RECT 66.140 165.645 67.955 166.555 ;
        RECT 67.965 165.645 69.335 166.455 ;
        RECT 69.345 165.645 72.555 166.555 ;
        RECT 72.565 165.645 73.915 166.555 ;
        RECT 74.875 165.645 77.615 166.325 ;
        RECT 77.625 165.645 78.975 166.555 ;
        RECT 80.975 166.325 81.905 166.555 ;
        RECT 80.070 165.645 81.905 166.325 ;
        RECT 82.695 165.730 83.125 166.515 ;
        RECT 83.145 165.645 86.620 166.555 ;
        RECT 86.825 165.645 90.495 166.455 ;
        RECT 90.965 165.645 92.335 166.455 ;
        RECT 18.425 165.435 18.595 165.645 ;
        RECT 19.805 165.435 19.975 165.645 ;
        RECT 25.325 165.435 25.495 165.645 ;
        RECT 29.000 165.485 29.120 165.595 ;
        RECT 29.470 165.435 29.640 165.625 ;
        RECT 30.840 165.485 30.960 165.595 ;
        RECT 31.765 165.455 31.935 165.645 ;
        RECT 34.525 165.455 34.695 165.645 ;
        RECT 37.765 165.625 37.915 165.645 ;
        RECT 35.905 165.435 36.075 165.625 ;
        RECT 37.290 165.435 37.460 165.625 ;
        RECT 37.745 165.435 37.915 165.625 ;
        RECT 40.040 165.485 40.160 165.595 ;
        RECT 40.505 165.455 40.675 165.645 ;
        RECT 47.865 165.625 48.035 165.645 ;
        RECT 41.420 165.485 41.540 165.595 ;
        RECT 42.800 165.435 42.970 165.625 ;
        RECT 43.275 165.480 43.435 165.590 ;
        RECT 44.645 165.435 44.815 165.625 ;
        RECT 46.490 165.435 46.660 165.625 ;
        RECT 47.860 165.455 48.035 165.625 ;
        RECT 49.705 165.455 49.875 165.645 ;
        RECT 47.895 165.435 48.030 165.455 ;
        RECT 51.545 165.435 51.715 165.625 ;
        RECT 53.380 165.485 53.500 165.595 ;
        RECT 54.760 165.455 54.930 165.645 ;
        RECT 55.225 165.455 55.395 165.645 ;
        RECT 56.600 165.485 56.720 165.595 ;
        RECT 57.065 165.435 57.235 165.625 ;
        RECT 57.525 165.455 57.695 165.645 ;
        RECT 61.205 165.455 61.375 165.645 ;
        RECT 62.585 165.435 62.755 165.625 ;
        RECT 63.965 165.455 64.135 165.645 ;
        RECT 64.430 165.455 64.600 165.645 ;
        RECT 66.265 165.455 66.435 165.645 ;
        RECT 68.105 165.435 68.275 165.645 ;
        RECT 70.405 165.435 70.575 165.625 ;
        RECT 72.245 165.455 72.415 165.645 ;
        RECT 72.710 165.455 72.880 165.645 ;
        RECT 74.085 165.435 74.255 165.625 ;
        RECT 76.845 165.435 77.015 165.625 ;
        RECT 77.305 165.455 77.475 165.645 ;
        RECT 77.770 165.455 77.940 165.645 ;
        RECT 80.070 165.625 80.235 165.645 ;
        RECT 79.155 165.490 79.315 165.600 ;
        RECT 80.065 165.435 80.235 165.625 ;
        RECT 80.525 165.435 80.695 165.625 ;
        RECT 82.365 165.595 82.535 165.625 ;
        RECT 82.360 165.485 82.535 165.595 ;
        RECT 82.365 165.435 82.535 165.485 ;
        RECT 83.290 165.455 83.460 165.645 ;
        RECT 86.965 165.455 87.135 165.645 ;
        RECT 90.640 165.485 90.760 165.595 ;
        RECT 92.025 165.435 92.195 165.645 ;
        RECT 18.285 164.625 19.655 165.435 ;
        RECT 19.665 164.625 25.175 165.435 ;
        RECT 25.185 164.625 28.855 165.435 ;
        RECT 29.325 164.755 32.995 165.435 ;
        RECT 29.325 164.525 30.250 164.755 ;
        RECT 33.005 164.525 36.175 165.435 ;
        RECT 36.225 164.525 37.575 165.435 ;
        RECT 37.605 164.625 41.275 165.435 ;
        RECT 41.765 164.525 43.115 165.435 ;
        RECT 44.055 164.565 44.485 165.350 ;
        RECT 44.505 164.625 46.335 165.435 ;
        RECT 46.345 164.525 47.695 165.435 ;
        RECT 47.895 164.525 51.395 165.435 ;
        RECT 51.405 164.625 56.915 165.435 ;
        RECT 56.925 164.625 62.435 165.435 ;
        RECT 62.445 164.625 67.955 165.435 ;
        RECT 67.965 164.625 69.795 165.435 ;
        RECT 69.815 164.565 70.245 165.350 ;
        RECT 70.265 164.625 73.935 165.435 ;
        RECT 73.945 164.625 75.315 165.435 ;
        RECT 75.325 164.525 77.140 165.435 ;
        RECT 78.085 164.755 80.375 165.435 ;
        RECT 78.085 164.525 79.005 164.755 ;
        RECT 80.385 164.625 82.215 165.435 ;
        RECT 82.225 164.755 90.925 165.435 ;
        RECT 85.770 164.535 86.680 164.755 ;
        RECT 88.220 164.525 90.925 164.755 ;
        RECT 90.965 164.625 92.335 165.435 ;
      LAYER nwell ;
        RECT 18.090 161.405 92.530 164.235 ;
      LAYER pwell ;
        RECT 18.285 160.205 19.655 161.015 ;
        RECT 19.665 160.205 22.415 161.015 ;
        RECT 25.940 160.885 26.850 161.105 ;
        RECT 28.385 160.885 29.735 161.115 ;
        RECT 22.425 160.205 29.735 160.885 ;
        RECT 29.785 160.205 31.135 161.115 ;
        RECT 31.175 160.290 31.605 161.075 ;
        RECT 31.625 160.205 34.375 161.015 ;
        RECT 34.845 160.915 35.790 161.115 ;
        RECT 37.125 160.915 38.055 161.115 ;
        RECT 34.845 160.435 38.055 160.915 ;
        RECT 34.845 160.235 37.915 160.435 ;
        RECT 34.845 160.205 35.790 160.235 ;
        RECT 18.425 159.995 18.595 160.205 ;
        RECT 19.805 159.995 19.975 160.205 ;
        RECT 22.565 160.015 22.735 160.205 ;
        RECT 25.325 159.995 25.495 160.185 ;
        RECT 29.930 160.015 30.100 160.205 ;
        RECT 30.845 159.995 31.015 160.185 ;
        RECT 31.765 160.015 31.935 160.205 ;
        RECT 33.600 160.045 33.720 160.155 ;
        RECT 34.065 159.995 34.235 160.185 ;
        RECT 34.520 160.045 34.640 160.155 ;
        RECT 36.830 159.995 37.000 160.185 ;
        RECT 37.295 160.040 37.455 160.150 ;
        RECT 37.745 160.015 37.915 160.235 ;
        RECT 38.065 160.205 39.415 161.115 ;
        RECT 39.445 160.205 43.115 161.015 ;
        RECT 44.215 160.205 47.715 161.115 ;
        RECT 49.805 160.885 51.395 161.115 ;
        RECT 47.725 160.205 51.395 160.885 ;
        RECT 51.415 160.205 52.765 161.115 ;
        RECT 53.345 160.205 56.455 161.115 ;
        RECT 56.935 160.290 57.365 161.075 ;
        RECT 60.130 160.885 61.055 161.115 ;
        RECT 57.385 160.205 61.055 160.885 ;
        RECT 61.985 160.205 64.735 161.115 ;
        RECT 64.760 160.205 66.575 161.115 ;
        RECT 66.585 160.205 69.335 161.015 ;
        RECT 69.805 160.205 71.635 161.115 ;
        RECT 71.665 160.205 73.015 161.115 ;
        RECT 73.025 160.205 76.695 161.015 ;
        RECT 76.705 160.205 78.075 161.015 ;
        RECT 78.165 160.205 81.615 161.115 ;
        RECT 82.695 160.290 83.125 161.075 ;
        RECT 83.240 160.885 84.160 161.115 ;
        RECT 86.825 160.885 87.960 161.115 ;
        RECT 83.240 160.205 86.705 160.885 ;
        RECT 86.825 160.205 90.035 160.885 ;
        RECT 90.965 160.205 92.335 161.015 ;
        RECT 38.210 160.015 38.380 160.205 ;
        RECT 39.585 160.015 39.755 160.205 ;
        RECT 44.215 160.185 44.350 160.205 ;
        RECT 41.425 159.995 41.595 160.185 ;
        RECT 42.800 159.995 42.970 160.185 ;
        RECT 43.275 160.040 43.435 160.160 ;
        RECT 44.180 160.015 44.350 160.185 ;
        RECT 44.655 160.040 44.815 160.150 ;
        RECT 45.565 159.995 45.735 160.185 ;
        RECT 47.870 160.015 48.040 160.205 ;
        RECT 49.245 159.995 49.415 160.185 ;
        RECT 49.705 159.995 49.875 160.185 ;
        RECT 52.465 160.015 52.635 160.205 ;
        RECT 52.920 160.045 53.040 160.155 ;
        RECT 53.385 160.015 53.555 160.205 ;
        RECT 54.300 159.995 54.470 160.185 ;
        RECT 54.765 159.995 54.935 160.185 ;
        RECT 56.600 160.045 56.720 160.155 ;
        RECT 60.740 160.015 60.910 160.205 ;
        RECT 61.215 160.050 61.375 160.160 ;
        RECT 62.125 160.015 62.295 160.205 ;
        RECT 63.965 159.995 64.135 160.185 ;
        RECT 64.885 160.015 65.055 160.205 ;
        RECT 66.725 160.015 66.895 160.205 ;
        RECT 69.025 159.995 69.195 160.185 ;
        RECT 69.480 160.045 69.600 160.155 ;
        RECT 69.950 160.015 70.120 160.205 ;
        RECT 70.405 159.995 70.575 160.185 ;
        RECT 71.780 160.015 71.950 160.205 ;
        RECT 73.165 159.995 73.335 160.205 ;
        RECT 73.625 159.995 73.795 160.185 ;
        RECT 75.465 159.995 75.635 160.185 ;
        RECT 76.845 160.015 77.015 160.205 ;
        RECT 78.225 159.995 78.395 160.205 ;
        RECT 79.605 159.995 79.775 160.185 ;
        RECT 81.915 160.050 82.075 160.160 ;
        RECT 86.505 160.015 86.675 160.205 ;
        RECT 88.345 159.995 88.515 160.185 ;
        RECT 89.725 160.015 89.895 160.205 ;
        RECT 90.195 160.050 90.355 160.160 ;
        RECT 92.025 159.995 92.195 160.205 ;
        RECT 18.285 159.185 19.655 159.995 ;
        RECT 19.665 159.185 25.175 159.995 ;
        RECT 25.185 159.185 30.695 159.995 ;
        RECT 30.705 159.185 33.455 159.995 ;
        RECT 33.940 159.085 35.755 159.995 ;
        RECT 35.765 159.085 37.115 159.995 ;
        RECT 38.160 159.315 41.625 159.995 ;
        RECT 38.160 159.085 39.080 159.315 ;
        RECT 41.765 159.085 43.115 159.995 ;
        RECT 44.055 159.125 44.485 159.910 ;
        RECT 45.440 159.085 47.255 159.995 ;
        RECT 47.265 159.315 49.555 159.995 ;
        RECT 49.675 159.315 53.140 159.995 ;
        RECT 47.265 159.085 48.185 159.315 ;
        RECT 52.220 159.085 53.140 159.315 ;
        RECT 53.265 159.085 54.615 159.995 ;
        RECT 54.625 159.315 63.730 159.995 ;
        RECT 63.825 159.185 65.655 159.995 ;
        RECT 65.760 159.315 69.225 159.995 ;
        RECT 65.760 159.085 66.680 159.315 ;
        RECT 69.815 159.125 70.245 159.910 ;
        RECT 70.265 159.185 71.635 159.995 ;
        RECT 71.645 159.085 73.460 159.995 ;
        RECT 73.485 159.185 75.315 159.995 ;
        RECT 75.325 159.315 78.065 159.995 ;
        RECT 78.085 159.185 79.455 159.995 ;
        RECT 79.465 159.315 88.165 159.995 ;
        RECT 83.010 159.095 83.920 159.315 ;
        RECT 85.460 159.085 88.165 159.315 ;
        RECT 88.205 159.185 90.955 159.995 ;
        RECT 90.965 159.185 92.335 159.995 ;
      LAYER nwell ;
        RECT 18.090 155.965 92.530 158.795 ;
      LAYER pwell ;
        RECT 18.285 154.765 19.655 155.575 ;
        RECT 19.665 154.765 25.175 155.575 ;
        RECT 25.185 154.765 30.695 155.575 ;
        RECT 31.175 154.850 31.605 155.635 ;
        RECT 35.600 155.445 36.510 155.665 ;
        RECT 38.045 155.445 39.395 155.675 ;
        RECT 43.880 155.445 44.790 155.665 ;
        RECT 46.325 155.445 47.675 155.675 ;
        RECT 32.085 154.765 39.395 155.445 ;
        RECT 40.365 154.765 47.675 155.445 ;
        RECT 47.725 154.765 49.555 155.575 ;
        RECT 49.605 155.445 50.955 155.675 ;
        RECT 52.490 155.445 53.400 155.665 ;
        RECT 49.605 154.765 56.915 155.445 ;
        RECT 56.935 154.850 57.365 155.635 ;
        RECT 57.385 154.765 60.135 155.575 ;
        RECT 63.660 155.445 64.570 155.665 ;
        RECT 66.105 155.445 67.455 155.675 ;
        RECT 60.145 154.765 67.455 155.445 ;
        RECT 67.505 154.765 71.175 155.575 ;
        RECT 75.650 155.445 76.560 155.665 ;
        RECT 78.100 155.445 80.805 155.675 ;
        RECT 72.105 154.765 80.805 155.445 ;
        RECT 80.845 154.765 82.675 155.575 ;
        RECT 82.695 154.850 83.125 155.635 ;
        RECT 83.145 154.765 88.655 155.575 ;
        RECT 88.665 154.765 90.495 155.575 ;
        RECT 90.965 154.765 92.335 155.575 ;
        RECT 18.425 154.555 18.595 154.765 ;
        RECT 19.805 154.555 19.975 154.765 ;
        RECT 25.325 154.555 25.495 154.765 ;
        RECT 30.845 154.715 31.015 154.745 ;
        RECT 30.840 154.605 31.015 154.715 ;
        RECT 31.760 154.605 31.880 154.715 ;
        RECT 30.845 154.555 31.015 154.605 ;
        RECT 32.225 154.575 32.395 154.765 ;
        RECT 36.365 154.555 36.535 154.745 ;
        RECT 39.595 154.610 39.755 154.720 ;
        RECT 40.505 154.575 40.675 154.765 ;
        RECT 41.885 154.555 42.055 154.745 ;
        RECT 43.720 154.605 43.840 154.715 ;
        RECT 44.645 154.555 44.815 154.745 ;
        RECT 47.865 154.575 48.035 154.765 ;
        RECT 50.165 154.555 50.335 154.745 ;
        RECT 55.685 154.555 55.855 154.745 ;
        RECT 56.605 154.575 56.775 154.765 ;
        RECT 57.525 154.575 57.695 154.765 ;
        RECT 60.285 154.575 60.455 154.765 ;
        RECT 61.205 154.555 61.375 154.745 ;
        RECT 66.725 154.555 66.895 154.745 ;
        RECT 67.645 154.575 67.815 154.765 ;
        RECT 69.480 154.605 69.600 154.715 ;
        RECT 70.405 154.555 70.575 154.745 ;
        RECT 71.335 154.610 71.495 154.720 ;
        RECT 72.245 154.575 72.415 154.765 ;
        RECT 75.925 154.555 76.095 154.745 ;
        RECT 80.985 154.575 81.155 154.765 ;
        RECT 81.445 154.555 81.615 154.745 ;
        RECT 83.285 154.575 83.455 154.765 ;
        RECT 86.965 154.555 87.135 154.745 ;
        RECT 88.805 154.575 88.975 154.765 ;
        RECT 90.640 154.605 90.760 154.715 ;
        RECT 92.025 154.555 92.195 154.765 ;
        RECT 18.285 153.745 19.655 154.555 ;
        RECT 19.665 153.745 25.175 154.555 ;
        RECT 25.185 153.745 30.695 154.555 ;
        RECT 30.705 153.745 36.215 154.555 ;
        RECT 36.225 153.745 41.735 154.555 ;
        RECT 41.745 153.745 43.575 154.555 ;
        RECT 44.055 153.685 44.485 154.470 ;
        RECT 44.505 153.745 50.015 154.555 ;
        RECT 50.025 153.745 55.535 154.555 ;
        RECT 55.545 153.745 61.055 154.555 ;
        RECT 61.065 153.745 66.575 154.555 ;
        RECT 66.585 153.745 69.335 154.555 ;
        RECT 69.815 153.685 70.245 154.470 ;
        RECT 70.265 153.745 75.775 154.555 ;
        RECT 75.785 153.745 81.295 154.555 ;
        RECT 81.305 153.745 86.815 154.555 ;
        RECT 86.825 153.745 90.495 154.555 ;
        RECT 90.965 153.745 92.335 154.555 ;
      LAYER nwell ;
        RECT 18.090 150.525 92.530 153.355 ;
      LAYER pwell ;
        RECT 18.285 149.325 19.655 150.135 ;
        RECT 19.665 149.325 25.175 150.135 ;
        RECT 25.185 149.325 30.695 150.135 ;
        RECT 31.175 149.410 31.605 150.195 ;
        RECT 31.625 149.325 37.135 150.135 ;
        RECT 37.145 149.325 42.655 150.135 ;
        RECT 42.665 149.325 48.175 150.135 ;
        RECT 48.185 149.325 53.695 150.135 ;
        RECT 53.705 149.325 56.455 150.135 ;
        RECT 56.935 149.410 57.365 150.195 ;
        RECT 57.385 149.325 62.895 150.135 ;
        RECT 67.370 150.005 68.280 150.225 ;
        RECT 69.820 150.005 72.525 150.235 ;
        RECT 63.825 149.325 72.525 150.005 ;
        RECT 72.565 149.325 78.075 150.135 ;
        RECT 78.085 149.325 81.755 150.135 ;
        RECT 82.695 149.410 83.125 150.195 ;
        RECT 83.145 149.325 88.655 150.135 ;
        RECT 88.665 149.325 90.495 150.135 ;
        RECT 90.965 149.325 92.335 150.135 ;
        RECT 18.425 149.115 18.595 149.325 ;
        RECT 19.805 149.115 19.975 149.325 ;
        RECT 25.325 149.115 25.495 149.325 ;
        RECT 30.845 149.275 31.015 149.305 ;
        RECT 30.840 149.165 31.015 149.275 ;
        RECT 30.845 149.115 31.015 149.165 ;
        RECT 31.765 149.135 31.935 149.325 ;
        RECT 36.365 149.115 36.535 149.305 ;
        RECT 37.285 149.135 37.455 149.325 ;
        RECT 41.885 149.115 42.055 149.305 ;
        RECT 42.805 149.135 42.975 149.325 ;
        RECT 43.720 149.165 43.840 149.275 ;
        RECT 44.645 149.115 44.815 149.305 ;
        RECT 48.325 149.135 48.495 149.325 ;
        RECT 50.165 149.115 50.335 149.305 ;
        RECT 53.845 149.135 54.015 149.325 ;
        RECT 55.685 149.115 55.855 149.305 ;
        RECT 56.600 149.165 56.720 149.275 ;
        RECT 57.525 149.135 57.695 149.325 ;
        RECT 61.205 149.115 61.375 149.305 ;
        RECT 63.055 149.170 63.215 149.280 ;
        RECT 63.965 149.135 64.135 149.325 ;
        RECT 66.725 149.115 66.895 149.305 ;
        RECT 69.480 149.165 69.600 149.275 ;
        RECT 70.405 149.115 70.575 149.305 ;
        RECT 72.705 149.135 72.875 149.325 ;
        RECT 75.925 149.115 76.095 149.305 ;
        RECT 78.225 149.135 78.395 149.325 ;
        RECT 81.445 149.115 81.615 149.305 ;
        RECT 81.915 149.170 82.075 149.280 ;
        RECT 83.285 149.135 83.455 149.325 ;
        RECT 86.965 149.115 87.135 149.305 ;
        RECT 88.805 149.135 88.975 149.325 ;
        RECT 90.640 149.165 90.760 149.275 ;
        RECT 92.025 149.115 92.195 149.325 ;
        RECT 18.285 148.305 19.655 149.115 ;
        RECT 19.665 148.305 25.175 149.115 ;
        RECT 25.185 148.305 30.695 149.115 ;
        RECT 30.705 148.305 36.215 149.115 ;
        RECT 36.225 148.305 41.735 149.115 ;
        RECT 41.745 148.305 43.575 149.115 ;
        RECT 44.055 148.245 44.485 149.030 ;
        RECT 44.505 148.305 50.015 149.115 ;
        RECT 50.025 148.305 55.535 149.115 ;
        RECT 55.545 148.305 61.055 149.115 ;
        RECT 61.065 148.305 66.575 149.115 ;
        RECT 66.585 148.305 69.335 149.115 ;
        RECT 69.815 148.245 70.245 149.030 ;
        RECT 70.265 148.305 75.775 149.115 ;
        RECT 75.785 148.305 81.295 149.115 ;
        RECT 81.305 148.305 86.815 149.115 ;
        RECT 86.825 148.305 90.495 149.115 ;
        RECT 90.965 148.305 92.335 149.115 ;
      LAYER nwell ;
        RECT 18.090 145.085 92.530 147.915 ;
      LAYER pwell ;
        RECT 18.285 143.885 19.655 144.695 ;
        RECT 19.665 143.885 25.175 144.695 ;
        RECT 25.185 143.885 30.695 144.695 ;
        RECT 31.175 143.970 31.605 144.755 ;
        RECT 31.625 143.885 37.135 144.695 ;
        RECT 37.145 143.885 42.655 144.695 ;
        RECT 42.665 143.885 48.175 144.695 ;
        RECT 48.185 143.885 53.695 144.695 ;
        RECT 53.705 143.885 56.455 144.695 ;
        RECT 56.935 143.970 57.365 144.755 ;
        RECT 57.385 143.885 62.895 144.695 ;
        RECT 62.905 143.885 68.415 144.695 ;
        RECT 68.425 143.885 73.935 144.695 ;
        RECT 73.945 143.885 79.455 144.695 ;
        RECT 79.465 143.885 82.215 144.695 ;
        RECT 82.695 143.970 83.125 144.755 ;
        RECT 83.145 143.885 88.655 144.695 ;
        RECT 88.665 143.885 90.495 144.695 ;
        RECT 90.965 143.885 92.335 144.695 ;
        RECT 18.425 143.675 18.595 143.885 ;
        RECT 19.805 143.675 19.975 143.885 ;
        RECT 25.325 143.675 25.495 143.885 ;
        RECT 30.845 143.835 31.015 143.865 ;
        RECT 30.840 143.725 31.015 143.835 ;
        RECT 30.845 143.675 31.015 143.725 ;
        RECT 31.765 143.695 31.935 143.885 ;
        RECT 36.365 143.675 36.535 143.865 ;
        RECT 37.285 143.695 37.455 143.885 ;
        RECT 41.885 143.675 42.055 143.865 ;
        RECT 42.805 143.695 42.975 143.885 ;
        RECT 43.720 143.725 43.840 143.835 ;
        RECT 44.645 143.675 44.815 143.865 ;
        RECT 48.325 143.695 48.495 143.885 ;
        RECT 50.165 143.675 50.335 143.865 ;
        RECT 53.845 143.695 54.015 143.885 ;
        RECT 55.685 143.675 55.855 143.865 ;
        RECT 56.600 143.725 56.720 143.835 ;
        RECT 57.525 143.695 57.695 143.885 ;
        RECT 61.205 143.675 61.375 143.865 ;
        RECT 63.045 143.695 63.215 143.885 ;
        RECT 66.725 143.675 66.895 143.865 ;
        RECT 68.565 143.695 68.735 143.885 ;
        RECT 69.480 143.725 69.600 143.835 ;
        RECT 70.405 143.675 70.575 143.865 ;
        RECT 74.085 143.695 74.255 143.885 ;
        RECT 75.925 143.675 76.095 143.865 ;
        RECT 79.605 143.695 79.775 143.885 ;
        RECT 81.445 143.675 81.615 143.865 ;
        RECT 82.360 143.725 82.480 143.835 ;
        RECT 83.285 143.695 83.455 143.885 ;
        RECT 86.965 143.675 87.135 143.865 ;
        RECT 88.805 143.695 88.975 143.885 ;
        RECT 90.640 143.725 90.760 143.835 ;
        RECT 92.025 143.675 92.195 143.885 ;
        RECT 18.285 142.865 19.655 143.675 ;
        RECT 19.665 142.865 25.175 143.675 ;
        RECT 25.185 142.865 30.695 143.675 ;
        RECT 30.705 142.865 36.215 143.675 ;
        RECT 36.225 142.865 41.735 143.675 ;
        RECT 41.745 142.865 43.575 143.675 ;
        RECT 44.055 142.805 44.485 143.590 ;
        RECT 44.505 142.865 50.015 143.675 ;
        RECT 50.025 142.865 55.535 143.675 ;
        RECT 55.545 142.865 61.055 143.675 ;
        RECT 61.065 142.865 66.575 143.675 ;
        RECT 66.585 142.865 69.335 143.675 ;
        RECT 69.815 142.805 70.245 143.590 ;
        RECT 70.265 142.865 75.775 143.675 ;
        RECT 75.785 142.865 81.295 143.675 ;
        RECT 81.305 142.865 86.815 143.675 ;
        RECT 86.825 142.865 90.495 143.675 ;
        RECT 90.965 142.865 92.335 143.675 ;
      LAYER nwell ;
        RECT 18.090 139.645 92.530 142.475 ;
      LAYER pwell ;
        RECT 18.285 138.445 19.655 139.255 ;
        RECT 19.665 138.445 25.175 139.255 ;
        RECT 25.185 138.445 30.695 139.255 ;
        RECT 31.175 138.530 31.605 139.315 ;
        RECT 31.625 138.445 37.135 139.255 ;
        RECT 37.145 138.445 42.655 139.255 ;
        RECT 42.665 138.445 48.175 139.255 ;
        RECT 48.185 138.445 53.695 139.255 ;
        RECT 53.705 138.445 56.455 139.255 ;
        RECT 56.935 138.530 57.365 139.315 ;
        RECT 57.385 138.445 62.895 139.255 ;
        RECT 62.905 138.445 68.415 139.255 ;
        RECT 68.425 138.445 73.935 139.255 ;
        RECT 73.945 138.445 79.455 139.255 ;
        RECT 79.465 138.445 82.215 139.255 ;
        RECT 82.695 138.530 83.125 139.315 ;
        RECT 83.145 138.445 88.655 139.255 ;
        RECT 88.665 138.445 90.495 139.255 ;
        RECT 90.965 138.445 92.335 139.255 ;
        RECT 18.425 138.235 18.595 138.445 ;
        RECT 19.805 138.235 19.975 138.445 ;
        RECT 25.325 138.235 25.495 138.445 ;
        RECT 30.845 138.395 31.015 138.425 ;
        RECT 30.840 138.285 31.015 138.395 ;
        RECT 30.845 138.235 31.015 138.285 ;
        RECT 31.765 138.255 31.935 138.445 ;
        RECT 36.365 138.235 36.535 138.425 ;
        RECT 37.285 138.255 37.455 138.445 ;
        RECT 41.885 138.235 42.055 138.425 ;
        RECT 42.805 138.255 42.975 138.445 ;
        RECT 43.720 138.285 43.840 138.395 ;
        RECT 44.645 138.235 44.815 138.425 ;
        RECT 48.325 138.255 48.495 138.445 ;
        RECT 50.165 138.235 50.335 138.425 ;
        RECT 53.845 138.255 54.015 138.445 ;
        RECT 55.685 138.235 55.855 138.425 ;
        RECT 56.600 138.285 56.720 138.395 ;
        RECT 57.525 138.255 57.695 138.445 ;
        RECT 61.205 138.235 61.375 138.425 ;
        RECT 63.045 138.255 63.215 138.445 ;
        RECT 66.725 138.235 66.895 138.425 ;
        RECT 68.565 138.255 68.735 138.445 ;
        RECT 69.480 138.285 69.600 138.395 ;
        RECT 70.405 138.235 70.575 138.425 ;
        RECT 74.085 138.255 74.255 138.445 ;
        RECT 75.925 138.235 76.095 138.425 ;
        RECT 79.605 138.255 79.775 138.445 ;
        RECT 81.445 138.235 81.615 138.425 ;
        RECT 82.360 138.285 82.480 138.395 ;
        RECT 83.285 138.255 83.455 138.445 ;
        RECT 86.965 138.235 87.135 138.425 ;
        RECT 88.805 138.255 88.975 138.445 ;
        RECT 90.640 138.285 90.760 138.395 ;
        RECT 92.025 138.235 92.195 138.445 ;
        RECT 18.285 137.425 19.655 138.235 ;
        RECT 19.665 137.425 25.175 138.235 ;
        RECT 25.185 137.425 30.695 138.235 ;
        RECT 30.705 137.425 36.215 138.235 ;
        RECT 36.225 137.425 41.735 138.235 ;
        RECT 41.745 137.425 43.575 138.235 ;
        RECT 44.055 137.365 44.485 138.150 ;
        RECT 44.505 137.425 50.015 138.235 ;
        RECT 50.025 137.425 55.535 138.235 ;
        RECT 55.545 137.425 61.055 138.235 ;
        RECT 61.065 137.425 66.575 138.235 ;
        RECT 66.585 137.425 69.335 138.235 ;
        RECT 69.815 137.365 70.245 138.150 ;
        RECT 70.265 137.425 75.775 138.235 ;
        RECT 75.785 137.425 81.295 138.235 ;
        RECT 81.305 137.425 86.815 138.235 ;
        RECT 86.825 137.425 90.495 138.235 ;
        RECT 90.965 137.425 92.335 138.235 ;
      LAYER nwell ;
        RECT 18.090 134.205 92.530 137.035 ;
      LAYER pwell ;
        RECT 18.285 133.005 19.655 133.815 ;
        RECT 19.665 133.005 25.175 133.815 ;
        RECT 25.185 133.005 30.695 133.815 ;
        RECT 31.175 133.090 31.605 133.875 ;
        RECT 31.625 133.005 37.135 133.815 ;
        RECT 37.145 133.005 42.655 133.815 ;
        RECT 42.665 133.005 44.035 133.815 ;
        RECT 44.055 133.090 44.485 133.875 ;
        RECT 44.505 133.005 50.015 133.815 ;
        RECT 50.025 133.005 55.535 133.815 ;
        RECT 55.545 133.005 56.915 133.815 ;
        RECT 56.935 133.090 57.365 133.875 ;
        RECT 57.385 133.005 62.895 133.815 ;
        RECT 62.905 133.005 68.415 133.815 ;
        RECT 68.425 133.005 69.795 133.815 ;
        RECT 69.815 133.090 70.245 133.875 ;
        RECT 70.265 133.005 75.775 133.815 ;
        RECT 75.785 133.005 81.295 133.815 ;
        RECT 81.305 133.005 82.675 133.815 ;
        RECT 82.695 133.090 83.125 133.875 ;
        RECT 83.145 133.005 88.655 133.815 ;
        RECT 88.665 133.005 90.495 133.815 ;
        RECT 90.965 133.005 92.335 133.815 ;
        RECT 18.425 132.815 18.595 133.005 ;
        RECT 19.805 132.815 19.975 133.005 ;
        RECT 25.325 132.815 25.495 133.005 ;
        RECT 30.840 132.845 30.960 132.955 ;
        RECT 31.765 132.815 31.935 133.005 ;
        RECT 37.285 132.815 37.455 133.005 ;
        RECT 42.805 132.815 42.975 133.005 ;
        RECT 44.645 132.815 44.815 133.005 ;
        RECT 50.165 132.815 50.335 133.005 ;
        RECT 55.685 132.815 55.855 133.005 ;
        RECT 57.525 132.815 57.695 133.005 ;
        RECT 63.045 132.815 63.215 133.005 ;
        RECT 68.565 132.815 68.735 133.005 ;
        RECT 70.405 132.815 70.575 133.005 ;
        RECT 75.925 132.815 76.095 133.005 ;
        RECT 81.445 132.815 81.615 133.005 ;
        RECT 83.285 132.815 83.455 133.005 ;
        RECT 88.805 132.815 88.975 133.005 ;
        RECT 90.640 132.845 90.760 132.955 ;
        RECT 92.025 132.815 92.195 133.005 ;
      LAYER li1 ;
        RECT 18.280 206.255 92.340 206.425 ;
        RECT 18.365 205.165 19.575 206.255 ;
        RECT 19.745 205.820 25.090 206.255 ;
        RECT 18.365 204.455 18.885 204.995 ;
        RECT 19.055 204.625 19.575 205.165 ;
        RECT 18.365 203.705 19.575 204.455 ;
        RECT 21.330 204.250 21.670 205.080 ;
        RECT 23.150 204.570 23.500 205.820 ;
        RECT 26.375 205.530 26.705 206.255 ;
        RECT 19.745 203.705 25.090 204.250 ;
        RECT 26.185 203.875 26.705 205.360 ;
        RECT 26.875 204.535 27.395 206.085 ;
        RECT 27.655 205.325 27.825 206.085 ;
        RECT 28.005 205.495 28.335 206.255 ;
        RECT 27.655 205.155 28.320 205.325 ;
        RECT 28.505 205.180 28.775 206.085 ;
        RECT 28.150 205.010 28.320 205.155 ;
        RECT 27.585 204.605 27.915 204.975 ;
        RECT 28.150 204.680 28.435 205.010 ;
        RECT 28.150 204.425 28.320 204.680 ;
        RECT 26.875 203.705 27.215 204.365 ;
        RECT 27.655 204.255 28.320 204.425 ;
        RECT 28.605 204.380 28.775 205.180 ;
        RECT 28.945 205.165 30.615 206.255 ;
        RECT 27.655 203.875 27.825 204.255 ;
        RECT 28.005 203.705 28.335 204.085 ;
        RECT 28.515 203.875 28.775 204.380 ;
        RECT 28.945 204.475 29.695 204.995 ;
        RECT 29.865 204.645 30.615 205.165 ;
        RECT 31.245 205.090 31.535 206.255 ;
        RECT 31.705 205.165 32.915 206.255 ;
        RECT 28.945 203.705 30.615 204.475 ;
        RECT 31.705 204.455 32.225 204.995 ;
        RECT 32.395 204.625 32.915 205.165 ;
        RECT 33.085 205.285 33.355 206.055 ;
        RECT 33.525 205.475 33.855 206.255 ;
        RECT 34.060 205.650 34.245 206.055 ;
        RECT 34.415 205.830 34.750 206.255 ;
        RECT 34.060 205.475 34.725 205.650 ;
        RECT 33.085 205.115 34.215 205.285 ;
        RECT 31.245 203.705 31.535 204.430 ;
        RECT 31.705 203.705 32.915 204.455 ;
        RECT 33.085 204.205 33.255 205.115 ;
        RECT 33.425 204.365 33.785 204.945 ;
        RECT 33.965 204.615 34.215 205.115 ;
        RECT 34.385 204.445 34.725 205.475 ;
        RECT 34.925 205.165 38.435 206.255 ;
        RECT 34.040 204.275 34.725 204.445 ;
        RECT 34.925 204.475 36.575 204.995 ;
        RECT 36.745 204.645 38.435 205.165 ;
        RECT 39.525 205.285 39.795 206.055 ;
        RECT 39.965 205.475 40.295 206.255 ;
        RECT 40.500 205.650 40.685 206.055 ;
        RECT 40.855 205.830 41.190 206.255 ;
        RECT 40.500 205.475 41.165 205.650 ;
        RECT 39.525 205.115 40.655 205.285 ;
        RECT 33.085 203.875 33.345 204.205 ;
        RECT 33.555 203.705 33.830 204.185 ;
        RECT 34.040 203.875 34.245 204.275 ;
        RECT 34.415 203.705 34.750 204.105 ;
        RECT 34.925 203.705 38.435 204.475 ;
        RECT 39.525 204.205 39.695 205.115 ;
        RECT 39.865 204.365 40.225 204.945 ;
        RECT 40.405 204.615 40.655 205.115 ;
        RECT 40.825 204.445 41.165 205.475 ;
        RECT 41.365 205.165 43.955 206.255 ;
        RECT 40.480 204.275 41.165 204.445 ;
        RECT 41.365 204.475 42.575 204.995 ;
        RECT 42.745 204.645 43.955 205.165 ;
        RECT 44.125 205.090 44.415 206.255 ;
        RECT 44.585 205.115 44.860 206.085 ;
        RECT 45.070 205.455 45.350 206.255 ;
        RECT 45.520 205.745 47.135 206.075 ;
        RECT 45.520 205.405 46.695 205.575 ;
        RECT 45.520 205.285 45.690 205.405 ;
        RECT 45.030 205.115 45.690 205.285 ;
        RECT 39.525 203.875 39.785 204.205 ;
        RECT 39.995 203.705 40.270 204.185 ;
        RECT 40.480 203.875 40.685 204.275 ;
        RECT 40.855 203.705 41.190 204.105 ;
        RECT 41.365 203.705 43.955 204.475 ;
        RECT 44.125 203.705 44.415 204.430 ;
        RECT 44.585 204.380 44.755 205.115 ;
        RECT 45.030 204.945 45.200 205.115 ;
        RECT 45.950 204.945 46.195 205.235 ;
        RECT 46.365 205.115 46.695 205.405 ;
        RECT 46.955 204.945 47.125 205.505 ;
        RECT 47.375 205.115 47.635 206.255 ;
        RECT 47.885 205.325 48.065 206.085 ;
        RECT 48.245 205.495 48.575 206.255 ;
        RECT 47.885 205.155 48.560 205.325 ;
        RECT 48.745 205.180 49.015 206.085 ;
        RECT 48.390 205.010 48.560 205.155 ;
        RECT 44.925 204.615 45.200 204.945 ;
        RECT 45.370 204.615 46.195 204.945 ;
        RECT 46.410 204.615 47.125 204.945 ;
        RECT 47.295 204.695 47.630 204.945 ;
        RECT 45.030 204.445 45.200 204.615 ;
        RECT 46.875 204.525 47.125 204.615 ;
        RECT 47.825 204.605 48.165 204.975 ;
        RECT 48.390 204.680 48.665 205.010 ;
        RECT 44.585 204.035 44.860 204.380 ;
        RECT 45.030 204.275 46.695 204.445 ;
        RECT 45.050 203.705 45.425 204.105 ;
        RECT 45.595 203.925 45.765 204.275 ;
        RECT 45.935 203.705 46.265 204.105 ;
        RECT 46.435 203.875 46.695 204.275 ;
        RECT 46.875 204.105 47.205 204.525 ;
        RECT 47.375 203.705 47.635 204.525 ;
        RECT 48.390 204.425 48.560 204.680 ;
        RECT 47.895 204.255 48.560 204.425 ;
        RECT 48.835 204.380 49.015 205.180 ;
        RECT 49.185 205.165 51.775 206.255 ;
        RECT 47.895 203.875 48.065 204.255 ;
        RECT 48.245 203.705 48.575 204.085 ;
        RECT 48.755 203.875 49.015 204.380 ;
        RECT 49.185 204.475 50.395 204.995 ;
        RECT 50.565 204.645 51.775 205.165 ;
        RECT 52.485 205.325 52.665 206.085 ;
        RECT 52.845 205.495 53.175 206.255 ;
        RECT 52.485 205.155 53.160 205.325 ;
        RECT 53.345 205.180 53.615 206.085 ;
        RECT 52.990 205.010 53.160 205.155 ;
        RECT 52.425 204.605 52.765 204.975 ;
        RECT 52.990 204.680 53.265 205.010 ;
        RECT 49.185 203.705 51.775 204.475 ;
        RECT 52.990 204.425 53.160 204.680 ;
        RECT 52.495 204.255 53.160 204.425 ;
        RECT 53.435 204.380 53.615 205.180 ;
        RECT 53.785 205.165 56.375 206.255 ;
        RECT 52.495 203.875 52.665 204.255 ;
        RECT 52.845 203.705 53.175 204.085 ;
        RECT 53.355 203.875 53.615 204.380 ;
        RECT 53.785 204.475 54.995 204.995 ;
        RECT 55.165 204.645 56.375 205.165 ;
        RECT 57.005 205.090 57.295 206.255 ;
        RECT 57.465 205.115 57.725 206.255 ;
        RECT 57.965 205.745 59.580 206.075 ;
        RECT 57.975 204.945 58.145 205.505 ;
        RECT 58.405 205.405 59.580 205.575 ;
        RECT 59.750 205.455 60.030 206.255 ;
        RECT 58.405 205.115 58.735 205.405 ;
        RECT 59.410 205.285 59.580 205.405 ;
        RECT 58.905 204.945 59.150 205.235 ;
        RECT 59.410 205.115 60.070 205.285 ;
        RECT 60.240 205.115 60.515 206.085 ;
        RECT 59.900 204.945 60.070 205.115 ;
        RECT 57.470 204.695 57.805 204.945 ;
        RECT 57.975 204.615 58.690 204.945 ;
        RECT 58.905 204.615 59.730 204.945 ;
        RECT 59.900 204.615 60.175 204.945 ;
        RECT 57.975 204.525 58.225 204.615 ;
        RECT 53.785 203.705 56.375 204.475 ;
        RECT 57.005 203.705 57.295 204.430 ;
        RECT 57.465 203.705 57.725 204.525 ;
        RECT 57.895 204.105 58.225 204.525 ;
        RECT 59.900 204.445 60.070 204.615 ;
        RECT 58.405 204.275 60.070 204.445 ;
        RECT 60.345 204.380 60.515 205.115 ;
        RECT 58.405 203.875 58.665 204.275 ;
        RECT 58.835 203.705 59.165 204.105 ;
        RECT 59.335 203.925 59.505 204.275 ;
        RECT 59.675 203.705 60.050 204.105 ;
        RECT 60.240 204.035 60.515 204.380 ;
        RECT 60.685 205.180 60.955 206.085 ;
        RECT 61.125 205.495 61.455 206.255 ;
        RECT 61.635 205.325 61.815 206.085 ;
        RECT 60.685 204.380 60.865 205.180 ;
        RECT 61.140 205.155 61.815 205.325 ;
        RECT 62.065 205.165 63.275 206.255 ;
        RECT 61.140 205.010 61.310 205.155 ;
        RECT 61.035 204.680 61.310 205.010 ;
        RECT 61.140 204.425 61.310 204.680 ;
        RECT 61.535 204.605 61.875 204.975 ;
        RECT 62.065 204.455 62.585 204.995 ;
        RECT 62.755 204.625 63.275 205.165 ;
        RECT 63.445 205.115 63.720 206.085 ;
        RECT 63.930 205.455 64.210 206.255 ;
        RECT 64.380 205.745 65.995 206.075 ;
        RECT 64.380 205.405 65.555 205.575 ;
        RECT 64.380 205.285 64.550 205.405 ;
        RECT 63.890 205.115 64.550 205.285 ;
        RECT 60.685 203.875 60.945 204.380 ;
        RECT 61.140 204.255 61.805 204.425 ;
        RECT 61.125 203.705 61.455 204.085 ;
        RECT 61.635 203.875 61.805 204.255 ;
        RECT 62.065 203.705 63.275 204.455 ;
        RECT 63.445 204.380 63.615 205.115 ;
        RECT 63.890 204.945 64.060 205.115 ;
        RECT 64.810 204.945 65.055 205.235 ;
        RECT 65.225 205.115 65.555 205.405 ;
        RECT 65.815 204.945 65.985 205.505 ;
        RECT 66.235 205.115 66.495 206.255 ;
        RECT 66.745 205.325 66.925 206.085 ;
        RECT 67.105 205.495 67.435 206.255 ;
        RECT 66.745 205.155 67.420 205.325 ;
        RECT 67.605 205.180 67.875 206.085 ;
        RECT 67.250 205.010 67.420 205.155 ;
        RECT 63.785 204.615 64.060 204.945 ;
        RECT 64.230 204.615 65.055 204.945 ;
        RECT 65.270 204.615 65.985 204.945 ;
        RECT 66.155 204.695 66.490 204.945 ;
        RECT 63.890 204.445 64.060 204.615 ;
        RECT 65.735 204.525 65.985 204.615 ;
        RECT 66.685 204.605 67.025 204.975 ;
        RECT 67.250 204.680 67.525 205.010 ;
        RECT 63.445 204.035 63.720 204.380 ;
        RECT 63.890 204.275 65.555 204.445 ;
        RECT 63.910 203.705 64.285 204.105 ;
        RECT 64.455 203.925 64.625 204.275 ;
        RECT 64.795 203.705 65.125 204.105 ;
        RECT 65.295 203.875 65.555 204.275 ;
        RECT 65.735 204.105 66.065 204.525 ;
        RECT 66.235 203.705 66.495 204.525 ;
        RECT 67.250 204.425 67.420 204.680 ;
        RECT 66.755 204.255 67.420 204.425 ;
        RECT 67.695 204.380 67.875 205.180 ;
        RECT 68.045 205.165 69.715 206.255 ;
        RECT 66.755 203.875 66.925 204.255 ;
        RECT 67.105 203.705 67.435 204.085 ;
        RECT 67.615 203.875 67.875 204.380 ;
        RECT 68.045 204.475 68.795 204.995 ;
        RECT 68.965 204.645 69.715 205.165 ;
        RECT 69.885 205.090 70.175 206.255 ;
        RECT 70.345 205.165 72.015 206.255 ;
        RECT 70.345 204.475 71.095 204.995 ;
        RECT 71.265 204.645 72.015 205.165 ;
        RECT 72.185 205.115 72.460 206.085 ;
        RECT 72.670 205.455 72.950 206.255 ;
        RECT 73.120 205.745 74.735 206.075 ;
        RECT 73.120 205.405 74.295 205.575 ;
        RECT 73.120 205.285 73.290 205.405 ;
        RECT 72.630 205.115 73.290 205.285 ;
        RECT 68.045 203.705 69.715 204.475 ;
        RECT 69.885 203.705 70.175 204.430 ;
        RECT 70.345 203.705 72.015 204.475 ;
        RECT 72.185 204.380 72.355 205.115 ;
        RECT 72.630 204.945 72.800 205.115 ;
        RECT 73.550 204.945 73.795 205.235 ;
        RECT 73.965 205.115 74.295 205.405 ;
        RECT 74.555 204.945 74.725 205.505 ;
        RECT 74.975 205.115 75.235 206.255 ;
        RECT 75.485 205.325 75.665 206.085 ;
        RECT 75.845 205.495 76.175 206.255 ;
        RECT 75.485 205.155 76.160 205.325 ;
        RECT 76.345 205.180 76.615 206.085 ;
        RECT 75.990 205.010 76.160 205.155 ;
        RECT 72.525 204.615 72.800 204.945 ;
        RECT 72.970 204.615 73.795 204.945 ;
        RECT 74.010 204.615 74.725 204.945 ;
        RECT 74.895 204.695 75.230 204.945 ;
        RECT 72.630 204.445 72.800 204.615 ;
        RECT 74.475 204.525 74.725 204.615 ;
        RECT 75.425 204.605 75.765 204.975 ;
        RECT 75.990 204.680 76.265 205.010 ;
        RECT 72.185 204.035 72.460 204.380 ;
        RECT 72.630 204.275 74.295 204.445 ;
        RECT 72.650 203.705 73.025 204.105 ;
        RECT 73.195 203.925 73.365 204.275 ;
        RECT 73.535 203.705 73.865 204.105 ;
        RECT 74.035 203.875 74.295 204.275 ;
        RECT 74.475 204.105 74.805 204.525 ;
        RECT 74.975 203.705 75.235 204.525 ;
        RECT 75.990 204.425 76.160 204.680 ;
        RECT 75.495 204.255 76.160 204.425 ;
        RECT 76.435 204.380 76.615 205.180 ;
        RECT 76.785 205.165 77.995 206.255 ;
        RECT 75.495 203.875 75.665 204.255 ;
        RECT 75.845 203.705 76.175 204.085 ;
        RECT 76.355 203.875 76.615 204.380 ;
        RECT 76.785 204.455 77.305 204.995 ;
        RECT 77.475 204.625 77.995 205.165 ;
        RECT 78.245 205.325 78.425 206.085 ;
        RECT 78.605 205.495 78.935 206.255 ;
        RECT 78.245 205.155 78.920 205.325 ;
        RECT 79.105 205.180 79.375 206.085 ;
        RECT 78.750 205.010 78.920 205.155 ;
        RECT 78.185 204.605 78.525 204.975 ;
        RECT 78.750 204.680 79.025 205.010 ;
        RECT 76.785 203.705 77.995 204.455 ;
        RECT 78.750 204.425 78.920 204.680 ;
        RECT 78.255 204.255 78.920 204.425 ;
        RECT 79.195 204.380 79.375 205.180 ;
        RECT 79.545 205.165 81.215 206.255 ;
        RECT 78.255 203.875 78.425 204.255 ;
        RECT 78.605 203.705 78.935 204.085 ;
        RECT 79.115 203.875 79.375 204.380 ;
        RECT 79.545 204.475 80.295 204.995 ;
        RECT 80.465 204.645 81.215 205.165 ;
        RECT 81.385 205.115 81.665 206.255 ;
        RECT 81.835 205.105 82.165 206.085 ;
        RECT 82.335 205.115 82.595 206.255 ;
        RECT 81.395 204.675 81.730 204.945 ;
        RECT 81.900 204.505 82.070 205.105 ;
        RECT 82.765 205.090 83.055 206.255 ;
        RECT 83.225 205.165 84.435 206.255 ;
        RECT 82.240 204.695 82.575 204.945 ;
        RECT 79.545 203.705 81.215 204.475 ;
        RECT 81.385 203.705 81.695 204.505 ;
        RECT 81.900 203.875 82.595 204.505 ;
        RECT 83.225 204.455 83.745 204.995 ;
        RECT 83.915 204.625 84.435 205.165 ;
        RECT 84.695 205.325 84.865 206.085 ;
        RECT 85.045 205.495 85.375 206.255 ;
        RECT 84.695 205.155 85.360 205.325 ;
        RECT 85.545 205.180 85.815 206.085 ;
        RECT 85.190 205.010 85.360 205.155 ;
        RECT 84.625 204.605 84.955 204.975 ;
        RECT 85.190 204.680 85.475 205.010 ;
        RECT 82.765 203.705 83.055 204.430 ;
        RECT 83.225 203.705 84.435 204.455 ;
        RECT 85.190 204.425 85.360 204.680 ;
        RECT 84.695 204.255 85.360 204.425 ;
        RECT 85.645 204.380 85.815 205.180 ;
        RECT 85.985 205.165 89.495 206.255 ;
        RECT 84.695 203.875 84.865 204.255 ;
        RECT 85.045 203.705 85.375 204.085 ;
        RECT 85.555 203.875 85.815 204.380 ;
        RECT 85.985 204.475 87.635 204.995 ;
        RECT 87.805 204.645 89.495 205.165 ;
        RECT 89.665 205.180 89.935 206.085 ;
        RECT 90.105 205.495 90.435 206.255 ;
        RECT 90.615 205.325 90.795 206.085 ;
        RECT 85.985 203.705 89.495 204.475 ;
        RECT 89.665 204.380 89.845 205.180 ;
        RECT 90.120 205.155 90.795 205.325 ;
        RECT 91.045 205.165 92.255 206.255 ;
        RECT 90.120 205.010 90.290 205.155 ;
        RECT 90.015 204.680 90.290 205.010 ;
        RECT 90.120 204.425 90.290 204.680 ;
        RECT 90.515 204.605 90.855 204.975 ;
        RECT 91.045 204.625 91.565 205.165 ;
        RECT 91.735 204.455 92.255 204.995 ;
        RECT 89.665 203.875 89.925 204.380 ;
        RECT 90.120 204.255 90.785 204.425 ;
        RECT 90.105 203.705 90.435 204.085 ;
        RECT 90.615 203.875 90.785 204.255 ;
        RECT 91.045 203.705 92.255 204.455 ;
        RECT 18.280 203.535 92.340 203.705 ;
        RECT 18.365 202.785 19.575 203.535 ;
        RECT 18.365 202.245 18.885 202.785 ;
        RECT 19.745 202.765 23.255 203.535 ;
        RECT 24.350 202.985 24.605 203.275 ;
        RECT 24.775 203.155 25.105 203.535 ;
        RECT 24.350 202.815 25.100 202.985 ;
        RECT 19.055 202.075 19.575 202.615 ;
        RECT 19.745 202.245 21.395 202.765 ;
        RECT 21.565 202.075 23.255 202.595 ;
        RECT 18.365 200.985 19.575 202.075 ;
        RECT 19.745 200.985 23.255 202.075 ;
        RECT 24.350 201.995 24.700 202.645 ;
        RECT 24.870 201.825 25.100 202.815 ;
        RECT 24.350 201.655 25.100 201.825 ;
        RECT 24.350 201.155 24.605 201.655 ;
        RECT 24.775 200.985 25.105 201.485 ;
        RECT 25.275 201.155 25.445 203.275 ;
        RECT 25.805 203.175 26.135 203.535 ;
        RECT 26.305 203.145 26.800 203.315 ;
        RECT 27.005 203.145 27.860 203.315 ;
        RECT 25.675 201.955 26.135 203.005 ;
        RECT 25.615 201.170 25.940 201.955 ;
        RECT 26.305 201.785 26.475 203.145 ;
        RECT 26.645 202.235 26.995 202.855 ;
        RECT 27.165 202.635 27.520 202.855 ;
        RECT 27.165 202.045 27.335 202.635 ;
        RECT 27.690 202.435 27.860 203.145 ;
        RECT 28.735 203.075 29.065 203.535 ;
        RECT 29.275 203.175 29.625 203.345 ;
        RECT 28.065 202.605 28.855 202.855 ;
        RECT 29.275 202.785 29.535 203.175 ;
        RECT 29.845 203.085 30.795 203.365 ;
        RECT 30.965 203.095 31.155 203.535 ;
        RECT 31.325 203.155 32.395 203.325 ;
        RECT 29.025 202.435 29.195 202.615 ;
        RECT 26.305 201.615 26.700 201.785 ;
        RECT 26.870 201.655 27.335 202.045 ;
        RECT 27.505 202.265 29.195 202.435 ;
        RECT 26.530 201.485 26.700 201.615 ;
        RECT 27.505 201.485 27.675 202.265 ;
        RECT 29.365 202.095 29.535 202.785 ;
        RECT 28.035 201.925 29.535 202.095 ;
        RECT 29.725 202.125 29.935 202.915 ;
        RECT 30.105 202.295 30.455 202.915 ;
        RECT 30.625 202.305 30.795 203.085 ;
        RECT 31.325 202.925 31.495 203.155 ;
        RECT 30.965 202.755 31.495 202.925 ;
        RECT 30.965 202.475 31.185 202.755 ;
        RECT 31.665 202.585 31.905 202.985 ;
        RECT 30.625 202.135 31.030 202.305 ;
        RECT 31.365 202.215 31.905 202.585 ;
        RECT 32.075 202.800 32.395 203.155 ;
        RECT 32.640 203.075 32.945 203.535 ;
        RECT 33.115 202.825 33.365 203.355 ;
        RECT 32.075 202.625 32.400 202.800 ;
        RECT 32.075 202.325 32.990 202.625 ;
        RECT 32.250 202.295 32.990 202.325 ;
        RECT 29.725 201.965 30.400 202.125 ;
        RECT 30.860 202.045 31.030 202.135 ;
        RECT 29.725 201.955 30.690 201.965 ;
        RECT 29.365 201.785 29.535 201.925 ;
        RECT 26.110 200.985 26.360 201.445 ;
        RECT 26.530 201.155 26.780 201.485 ;
        RECT 26.995 201.155 27.675 201.485 ;
        RECT 27.845 201.585 28.920 201.755 ;
        RECT 29.365 201.615 29.925 201.785 ;
        RECT 30.230 201.665 30.690 201.955 ;
        RECT 30.860 201.875 32.080 202.045 ;
        RECT 27.845 201.245 28.015 201.585 ;
        RECT 28.250 200.985 28.580 201.415 ;
        RECT 28.750 201.245 28.920 201.585 ;
        RECT 29.215 200.985 29.585 201.445 ;
        RECT 29.755 201.155 29.925 201.615 ;
        RECT 30.860 201.495 31.030 201.875 ;
        RECT 32.250 201.705 32.420 202.295 ;
        RECT 33.160 202.175 33.365 202.825 ;
        RECT 33.535 202.780 33.785 203.535 ;
        RECT 34.005 203.035 34.305 203.365 ;
        RECT 34.475 203.055 34.750 203.535 ;
        RECT 30.160 201.155 31.030 201.495 ;
        RECT 31.620 201.535 32.420 201.705 ;
        RECT 31.200 200.985 31.450 201.445 ;
        RECT 31.620 201.245 31.790 201.535 ;
        RECT 31.970 200.985 32.300 201.365 ;
        RECT 32.640 200.985 32.945 202.125 ;
        RECT 33.115 201.295 33.365 202.175 ;
        RECT 34.005 202.125 34.175 203.035 ;
        RECT 34.930 202.885 35.225 203.275 ;
        RECT 35.395 203.055 35.650 203.535 ;
        RECT 35.825 202.885 36.085 203.275 ;
        RECT 36.255 203.055 36.535 203.535 ;
        RECT 36.855 202.985 37.025 203.275 ;
        RECT 37.195 203.155 37.525 203.535 ;
        RECT 34.345 202.295 34.695 202.865 ;
        RECT 34.930 202.715 36.580 202.885 ;
        RECT 36.855 202.815 37.520 202.985 ;
        RECT 34.865 202.375 36.005 202.545 ;
        RECT 34.865 202.125 35.035 202.375 ;
        RECT 36.175 202.205 36.580 202.715 ;
        RECT 33.535 200.985 33.785 202.125 ;
        RECT 34.005 201.955 35.035 202.125 ;
        RECT 35.825 202.035 36.580 202.205 ;
        RECT 34.005 201.155 34.315 201.955 ;
        RECT 35.445 201.785 35.615 201.835 ;
        RECT 35.825 201.785 36.085 202.035 ;
        RECT 36.770 201.995 37.120 202.645 ;
        RECT 34.485 200.985 34.795 201.785 ;
        RECT 34.965 201.615 36.085 201.785 ;
        RECT 34.965 201.155 35.225 201.615 ;
        RECT 35.395 200.985 35.650 201.445 ;
        RECT 35.825 201.155 36.085 201.615 ;
        RECT 36.255 200.985 36.540 201.855 ;
        RECT 37.290 201.825 37.520 202.815 ;
        RECT 36.855 201.655 37.520 201.825 ;
        RECT 36.855 201.155 37.025 201.655 ;
        RECT 37.195 200.985 37.525 201.485 ;
        RECT 37.695 201.155 37.880 203.275 ;
        RECT 38.135 203.075 38.385 203.535 ;
        RECT 38.555 203.085 38.890 203.255 ;
        RECT 39.085 203.085 39.760 203.255 ;
        RECT 38.555 202.945 38.725 203.085 ;
        RECT 38.050 201.955 38.330 202.905 ;
        RECT 38.500 202.815 38.725 202.945 ;
        RECT 38.500 201.710 38.670 202.815 ;
        RECT 38.895 202.665 39.420 202.885 ;
        RECT 38.840 201.900 39.080 202.495 ;
        RECT 39.250 201.965 39.420 202.665 ;
        RECT 39.590 202.305 39.760 203.085 ;
        RECT 40.080 203.035 40.450 203.535 ;
        RECT 40.630 203.085 41.035 203.255 ;
        RECT 41.205 203.085 41.990 203.255 ;
        RECT 40.630 202.855 40.800 203.085 ;
        RECT 39.970 202.555 40.800 202.855 ;
        RECT 41.185 202.585 41.650 202.915 ;
        RECT 39.970 202.525 40.170 202.555 ;
        RECT 40.290 202.305 40.460 202.375 ;
        RECT 39.590 202.135 40.460 202.305 ;
        RECT 39.950 202.045 40.460 202.135 ;
        RECT 38.500 201.580 38.805 201.710 ;
        RECT 39.250 201.600 39.780 201.965 ;
        RECT 38.120 200.985 38.385 201.445 ;
        RECT 38.555 201.155 38.805 201.580 ;
        RECT 39.950 201.430 40.120 202.045 ;
        RECT 39.015 201.260 40.120 201.430 ;
        RECT 40.290 200.985 40.460 201.785 ;
        RECT 40.630 201.485 40.800 202.555 ;
        RECT 40.970 201.655 41.160 202.375 ;
        RECT 41.330 201.625 41.650 202.585 ;
        RECT 41.820 202.625 41.990 203.085 ;
        RECT 42.265 203.005 42.475 203.535 ;
        RECT 42.735 202.795 43.065 203.320 ;
        RECT 43.235 202.925 43.405 203.535 ;
        RECT 43.575 202.880 43.905 203.315 ;
        RECT 43.575 202.795 43.955 202.880 ;
        RECT 44.125 202.810 44.415 203.535 ;
        RECT 42.865 202.625 43.065 202.795 ;
        RECT 43.730 202.755 43.955 202.795 ;
        RECT 41.820 202.295 42.695 202.625 ;
        RECT 42.865 202.295 43.615 202.625 ;
        RECT 40.630 201.155 40.880 201.485 ;
        RECT 41.820 201.455 41.990 202.295 ;
        RECT 42.865 202.090 43.055 202.295 ;
        RECT 43.785 202.175 43.955 202.755 ;
        RECT 43.740 202.125 43.955 202.175 ;
        RECT 42.160 201.715 43.055 202.090 ;
        RECT 43.565 202.045 43.955 202.125 ;
        RECT 41.105 201.285 41.990 201.455 ;
        RECT 42.170 200.985 42.485 201.485 ;
        RECT 42.715 201.155 43.055 201.715 ;
        RECT 43.225 200.985 43.395 201.995 ;
        RECT 43.565 201.200 43.895 202.045 ;
        RECT 44.125 200.985 44.415 202.150 ;
        RECT 45.065 201.955 45.295 203.295 ;
        RECT 45.475 202.455 45.705 203.355 ;
        RECT 45.905 202.755 46.150 203.535 ;
        RECT 46.320 202.995 46.750 203.355 ;
        RECT 47.330 203.165 48.060 203.535 ;
        RECT 46.320 202.805 48.060 202.995 ;
        RECT 46.320 202.575 46.540 202.805 ;
        RECT 45.475 201.775 45.815 202.455 ;
        RECT 45.065 201.575 45.815 201.775 ;
        RECT 45.995 202.275 46.540 202.575 ;
        RECT 45.065 201.185 45.305 201.575 ;
        RECT 45.475 200.985 45.825 201.395 ;
        RECT 45.995 201.165 46.325 202.275 ;
        RECT 46.710 202.005 47.135 202.625 ;
        RECT 47.330 202.005 47.590 202.625 ;
        RECT 47.800 202.295 48.060 202.805 ;
        RECT 46.495 201.635 47.520 201.835 ;
        RECT 46.495 201.165 46.675 201.635 ;
        RECT 46.845 200.985 47.175 201.465 ;
        RECT 47.350 201.165 47.520 201.635 ;
        RECT 47.785 200.985 48.070 202.125 ;
        RECT 48.260 201.165 48.540 203.355 ;
        RECT 48.815 202.985 48.985 203.365 ;
        RECT 49.200 203.155 49.530 203.535 ;
        RECT 48.815 202.815 49.530 202.985 ;
        RECT 48.725 202.265 49.080 202.635 ;
        RECT 49.360 202.625 49.530 202.815 ;
        RECT 49.700 202.790 49.955 203.365 ;
        RECT 49.360 202.295 49.615 202.625 ;
        RECT 49.360 202.085 49.530 202.295 ;
        RECT 48.815 201.915 49.530 202.085 ;
        RECT 49.785 202.060 49.955 202.790 ;
        RECT 50.130 202.695 50.390 203.535 ;
        RECT 50.615 202.880 50.945 203.315 ;
        RECT 51.115 202.925 51.285 203.535 ;
        RECT 50.565 202.795 50.945 202.880 ;
        RECT 51.455 202.795 51.785 203.320 ;
        RECT 52.045 203.005 52.255 203.535 ;
        RECT 52.530 203.085 53.315 203.255 ;
        RECT 53.485 203.085 53.890 203.255 ;
        RECT 50.565 202.755 50.790 202.795 ;
        RECT 50.565 202.175 50.735 202.755 ;
        RECT 51.455 202.625 51.655 202.795 ;
        RECT 52.530 202.625 52.700 203.085 ;
        RECT 50.905 202.295 51.655 202.625 ;
        RECT 51.825 202.295 52.700 202.625 ;
        RECT 48.815 201.155 48.985 201.915 ;
        RECT 49.200 200.985 49.530 201.745 ;
        RECT 49.700 201.155 49.955 202.060 ;
        RECT 50.130 200.985 50.390 202.135 ;
        RECT 50.565 202.125 50.780 202.175 ;
        RECT 50.565 202.045 50.955 202.125 ;
        RECT 50.625 201.200 50.955 202.045 ;
        RECT 51.465 202.090 51.655 202.295 ;
        RECT 51.125 200.985 51.295 201.995 ;
        RECT 51.465 201.715 52.360 202.090 ;
        RECT 51.465 201.155 51.805 201.715 ;
        RECT 52.035 200.985 52.350 201.485 ;
        RECT 52.530 201.455 52.700 202.295 ;
        RECT 52.870 202.585 53.335 202.915 ;
        RECT 53.720 202.855 53.890 203.085 ;
        RECT 54.070 203.035 54.440 203.535 ;
        RECT 54.760 203.085 55.435 203.255 ;
        RECT 55.630 203.085 55.965 203.255 ;
        RECT 52.870 201.625 53.190 202.585 ;
        RECT 53.720 202.555 54.550 202.855 ;
        RECT 53.360 201.655 53.550 202.375 ;
        RECT 53.720 201.485 53.890 202.555 ;
        RECT 54.350 202.525 54.550 202.555 ;
        RECT 54.060 202.305 54.230 202.375 ;
        RECT 54.760 202.305 54.930 203.085 ;
        RECT 55.795 202.945 55.965 203.085 ;
        RECT 56.135 203.075 56.385 203.535 ;
        RECT 54.060 202.135 54.930 202.305 ;
        RECT 55.100 202.665 55.625 202.885 ;
        RECT 55.795 202.815 56.020 202.945 ;
        RECT 54.060 202.045 54.570 202.135 ;
        RECT 52.530 201.285 53.415 201.455 ;
        RECT 53.640 201.155 53.890 201.485 ;
        RECT 54.060 200.985 54.230 201.785 ;
        RECT 54.400 201.430 54.570 202.045 ;
        RECT 55.100 201.965 55.270 202.665 ;
        RECT 54.740 201.600 55.270 201.965 ;
        RECT 55.440 201.900 55.680 202.495 ;
        RECT 55.850 201.710 56.020 202.815 ;
        RECT 56.190 201.955 56.470 202.905 ;
        RECT 55.715 201.580 56.020 201.710 ;
        RECT 54.400 201.260 55.505 201.430 ;
        RECT 55.715 201.155 55.965 201.580 ;
        RECT 56.135 200.985 56.400 201.445 ;
        RECT 56.640 201.155 56.825 203.275 ;
        RECT 56.995 203.155 57.325 203.535 ;
        RECT 57.495 202.985 57.665 203.275 ;
        RECT 57.000 202.815 57.665 202.985 ;
        RECT 57.000 201.825 57.230 202.815 ;
        RECT 57.925 202.765 59.595 203.535 ;
        RECT 60.275 202.880 60.605 203.315 ;
        RECT 60.775 202.925 60.945 203.535 ;
        RECT 60.225 202.795 60.605 202.880 ;
        RECT 61.115 202.795 61.445 203.320 ;
        RECT 61.705 203.005 61.915 203.535 ;
        RECT 62.190 203.085 62.975 203.255 ;
        RECT 63.145 203.085 63.550 203.255 ;
        RECT 57.400 201.995 57.750 202.645 ;
        RECT 57.925 202.245 58.675 202.765 ;
        RECT 60.225 202.755 60.450 202.795 ;
        RECT 58.845 202.075 59.595 202.595 ;
        RECT 57.000 201.655 57.665 201.825 ;
        RECT 56.995 200.985 57.325 201.485 ;
        RECT 57.495 201.155 57.665 201.655 ;
        RECT 57.925 200.985 59.595 202.075 ;
        RECT 60.225 202.175 60.395 202.755 ;
        RECT 61.115 202.625 61.315 202.795 ;
        RECT 62.190 202.625 62.360 203.085 ;
        RECT 60.565 202.295 61.315 202.625 ;
        RECT 61.485 202.295 62.360 202.625 ;
        RECT 60.225 202.125 60.440 202.175 ;
        RECT 60.225 202.045 60.615 202.125 ;
        RECT 60.285 201.200 60.615 202.045 ;
        RECT 61.125 202.090 61.315 202.295 ;
        RECT 60.785 200.985 60.955 201.995 ;
        RECT 61.125 201.715 62.020 202.090 ;
        RECT 61.125 201.155 61.465 201.715 ;
        RECT 61.695 200.985 62.010 201.485 ;
        RECT 62.190 201.455 62.360 202.295 ;
        RECT 62.530 202.585 62.995 202.915 ;
        RECT 63.380 202.855 63.550 203.085 ;
        RECT 63.730 203.035 64.100 203.535 ;
        RECT 64.420 203.085 65.095 203.255 ;
        RECT 65.290 203.085 65.625 203.255 ;
        RECT 62.530 201.625 62.850 202.585 ;
        RECT 63.380 202.555 64.210 202.855 ;
        RECT 63.020 201.655 63.210 202.375 ;
        RECT 63.380 201.485 63.550 202.555 ;
        RECT 64.010 202.525 64.210 202.555 ;
        RECT 63.720 202.305 63.890 202.375 ;
        RECT 64.420 202.305 64.590 203.085 ;
        RECT 65.455 202.945 65.625 203.085 ;
        RECT 65.795 203.075 66.045 203.535 ;
        RECT 63.720 202.135 64.590 202.305 ;
        RECT 64.760 202.665 65.285 202.885 ;
        RECT 65.455 202.815 65.680 202.945 ;
        RECT 63.720 202.045 64.230 202.135 ;
        RECT 62.190 201.285 63.075 201.455 ;
        RECT 63.300 201.155 63.550 201.485 ;
        RECT 63.720 200.985 63.890 201.785 ;
        RECT 64.060 201.430 64.230 202.045 ;
        RECT 64.760 201.965 64.930 202.665 ;
        RECT 64.400 201.600 64.930 201.965 ;
        RECT 65.100 201.900 65.340 202.495 ;
        RECT 65.510 201.710 65.680 202.815 ;
        RECT 65.850 201.955 66.130 202.905 ;
        RECT 65.375 201.580 65.680 201.710 ;
        RECT 64.060 201.260 65.165 201.430 ;
        RECT 65.375 201.155 65.625 201.580 ;
        RECT 65.795 200.985 66.060 201.445 ;
        RECT 66.300 201.155 66.485 203.275 ;
        RECT 66.655 203.155 66.985 203.535 ;
        RECT 67.155 202.985 67.325 203.275 ;
        RECT 66.660 202.815 67.325 202.985 ;
        RECT 66.660 201.825 66.890 202.815 ;
        RECT 67.585 202.765 69.255 203.535 ;
        RECT 69.885 202.810 70.175 203.535 ;
        RECT 70.395 202.880 70.725 203.315 ;
        RECT 70.895 202.925 71.065 203.535 ;
        RECT 70.345 202.795 70.725 202.880 ;
        RECT 71.235 202.795 71.565 203.320 ;
        RECT 71.825 203.005 72.035 203.535 ;
        RECT 72.310 203.085 73.095 203.255 ;
        RECT 73.265 203.085 73.670 203.255 ;
        RECT 67.060 201.995 67.410 202.645 ;
        RECT 67.585 202.245 68.335 202.765 ;
        RECT 70.345 202.755 70.570 202.795 ;
        RECT 68.505 202.075 69.255 202.595 ;
        RECT 70.345 202.175 70.515 202.755 ;
        RECT 71.235 202.625 71.435 202.795 ;
        RECT 72.310 202.625 72.480 203.085 ;
        RECT 70.685 202.295 71.435 202.625 ;
        RECT 71.605 202.295 72.480 202.625 ;
        RECT 66.660 201.655 67.325 201.825 ;
        RECT 66.655 200.985 66.985 201.485 ;
        RECT 67.155 201.155 67.325 201.655 ;
        RECT 67.585 200.985 69.255 202.075 ;
        RECT 69.885 200.985 70.175 202.150 ;
        RECT 70.345 202.125 70.560 202.175 ;
        RECT 70.345 202.045 70.735 202.125 ;
        RECT 70.405 201.200 70.735 202.045 ;
        RECT 71.245 202.090 71.435 202.295 ;
        RECT 70.905 200.985 71.075 201.995 ;
        RECT 71.245 201.715 72.140 202.090 ;
        RECT 71.245 201.155 71.585 201.715 ;
        RECT 71.815 200.985 72.130 201.485 ;
        RECT 72.310 201.455 72.480 202.295 ;
        RECT 72.650 202.585 73.115 202.915 ;
        RECT 73.500 202.855 73.670 203.085 ;
        RECT 73.850 203.035 74.220 203.535 ;
        RECT 74.540 203.085 75.215 203.255 ;
        RECT 75.410 203.085 75.745 203.255 ;
        RECT 72.650 201.625 72.970 202.585 ;
        RECT 73.500 202.555 74.330 202.855 ;
        RECT 73.140 201.655 73.330 202.375 ;
        RECT 73.500 201.485 73.670 202.555 ;
        RECT 74.130 202.525 74.330 202.555 ;
        RECT 73.840 202.305 74.010 202.375 ;
        RECT 74.540 202.305 74.710 203.085 ;
        RECT 75.575 202.945 75.745 203.085 ;
        RECT 75.915 203.075 76.165 203.535 ;
        RECT 73.840 202.135 74.710 202.305 ;
        RECT 74.880 202.665 75.405 202.885 ;
        RECT 75.575 202.815 75.800 202.945 ;
        RECT 73.840 202.045 74.350 202.135 ;
        RECT 72.310 201.285 73.195 201.455 ;
        RECT 73.420 201.155 73.670 201.485 ;
        RECT 73.840 200.985 74.010 201.785 ;
        RECT 74.180 201.430 74.350 202.045 ;
        RECT 74.880 201.965 75.050 202.665 ;
        RECT 74.520 201.600 75.050 201.965 ;
        RECT 75.220 201.900 75.460 202.495 ;
        RECT 75.630 201.710 75.800 202.815 ;
        RECT 75.970 201.955 76.250 202.905 ;
        RECT 75.495 201.580 75.800 201.710 ;
        RECT 74.180 201.260 75.285 201.430 ;
        RECT 75.495 201.155 75.745 201.580 ;
        RECT 75.915 200.985 76.180 201.445 ;
        RECT 76.420 201.155 76.605 203.275 ;
        RECT 76.775 203.155 77.105 203.535 ;
        RECT 77.275 202.985 77.445 203.275 ;
        RECT 76.780 202.815 77.445 202.985 ;
        RECT 78.635 202.815 78.965 203.535 ;
        RECT 79.510 203.135 81.125 203.305 ;
        RECT 81.295 203.135 81.625 203.535 ;
        RECT 80.955 202.965 81.125 203.135 ;
        RECT 81.795 203.060 82.130 203.320 ;
        RECT 76.780 201.825 77.010 202.815 ;
        RECT 77.180 201.995 77.530 202.645 ;
        RECT 78.690 202.295 79.040 202.625 ;
        RECT 79.350 202.295 79.770 202.960 ;
        RECT 79.940 202.515 80.230 202.955 ;
        RECT 80.420 202.515 80.690 202.955 ;
        RECT 80.955 202.795 81.515 202.965 ;
        RECT 81.345 202.625 81.515 202.795 ;
        RECT 80.900 202.515 81.150 202.625 ;
        RECT 79.940 202.345 80.235 202.515 ;
        RECT 80.420 202.345 80.695 202.515 ;
        RECT 80.900 202.345 81.155 202.515 ;
        RECT 79.940 202.295 80.230 202.345 ;
        RECT 80.420 202.295 80.690 202.345 ;
        RECT 80.900 202.295 81.150 202.345 ;
        RECT 81.345 202.295 81.650 202.625 ;
        RECT 78.690 202.175 78.895 202.295 ;
        RECT 78.685 202.005 78.895 202.175 ;
        RECT 81.345 202.125 81.515 202.295 ;
        RECT 79.145 201.955 81.515 202.125 ;
        RECT 76.780 201.655 77.445 201.825 ;
        RECT 76.775 200.985 77.105 201.485 ;
        RECT 77.275 201.155 77.445 201.655 ;
        RECT 78.715 201.325 78.885 201.825 ;
        RECT 79.145 201.495 79.315 201.955 ;
        RECT 79.545 201.575 80.970 201.745 ;
        RECT 79.545 201.325 79.875 201.575 ;
        RECT 78.715 201.155 79.875 201.325 ;
        RECT 80.100 200.985 80.430 201.405 ;
        RECT 80.685 201.155 80.970 201.575 ;
        RECT 81.215 200.985 81.545 201.785 ;
        RECT 81.875 201.705 82.130 203.060 ;
        RECT 82.395 202.985 82.565 203.275 ;
        RECT 82.735 203.155 83.065 203.535 ;
        RECT 82.395 202.815 83.060 202.985 ;
        RECT 82.310 201.995 82.660 202.645 ;
        RECT 82.830 201.825 83.060 202.815 ;
        RECT 81.795 201.195 82.130 201.705 ;
        RECT 82.395 201.655 83.060 201.825 ;
        RECT 82.395 201.155 82.565 201.655 ;
        RECT 82.735 200.985 83.065 201.485 ;
        RECT 83.235 201.155 83.460 203.275 ;
        RECT 83.675 203.075 83.925 203.535 ;
        RECT 84.110 203.085 84.440 203.255 ;
        RECT 84.620 203.085 85.370 203.255 ;
        RECT 83.660 201.955 83.940 202.555 ;
        RECT 84.110 201.555 84.280 203.085 ;
        RECT 84.450 202.585 85.030 202.915 ;
        RECT 84.450 201.715 84.690 202.585 ;
        RECT 85.200 202.305 85.370 203.085 ;
        RECT 85.620 203.035 85.990 203.535 ;
        RECT 86.170 203.085 86.630 203.255 ;
        RECT 86.860 203.085 87.530 203.255 ;
        RECT 86.170 202.855 86.340 203.085 ;
        RECT 85.540 202.555 86.340 202.855 ;
        RECT 86.510 202.585 87.060 202.915 ;
        RECT 85.540 202.525 85.710 202.555 ;
        RECT 85.830 202.305 86.000 202.375 ;
        RECT 85.200 202.135 86.000 202.305 ;
        RECT 85.490 202.045 86.000 202.135 ;
        RECT 84.880 201.610 85.320 201.965 ;
        RECT 83.660 200.985 83.925 201.445 ;
        RECT 84.110 201.180 84.345 201.555 ;
        RECT 85.490 201.430 85.660 202.045 ;
        RECT 84.590 201.260 85.660 201.430 ;
        RECT 85.830 200.985 86.000 201.785 ;
        RECT 86.170 201.485 86.340 202.555 ;
        RECT 86.510 201.655 86.700 202.375 ;
        RECT 86.870 202.045 87.060 202.585 ;
        RECT 87.360 202.545 87.530 203.085 ;
        RECT 87.845 203.005 88.015 203.535 ;
        RECT 88.310 202.885 88.670 203.325 ;
        RECT 88.845 203.055 89.015 203.535 ;
        RECT 89.205 202.890 89.540 203.315 ;
        RECT 89.715 203.060 89.885 203.535 ;
        RECT 90.060 202.890 90.395 203.315 ;
        RECT 90.565 203.060 90.735 203.535 ;
        RECT 88.310 202.715 88.810 202.885 ;
        RECT 89.205 202.720 90.875 202.890 ;
        RECT 91.045 202.785 92.255 203.535 ;
        RECT 88.640 202.545 88.810 202.715 ;
        RECT 87.360 202.375 88.450 202.545 ;
        RECT 88.640 202.375 90.460 202.545 ;
        RECT 86.870 201.715 87.190 202.045 ;
        RECT 86.170 201.155 86.420 201.485 ;
        RECT 87.360 201.455 87.530 202.375 ;
        RECT 88.640 202.120 88.810 202.375 ;
        RECT 90.630 202.155 90.875 202.720 ;
        RECT 87.700 201.950 88.810 202.120 ;
        RECT 89.205 201.985 90.875 202.155 ;
        RECT 91.045 202.075 91.565 202.615 ;
        RECT 91.735 202.245 92.255 202.785 ;
        RECT 87.700 201.790 88.560 201.950 ;
        RECT 86.645 201.285 87.530 201.455 ;
        RECT 87.710 200.985 87.925 201.485 ;
        RECT 88.390 201.165 88.560 201.790 ;
        RECT 88.845 200.985 89.025 201.765 ;
        RECT 89.205 201.225 89.540 201.985 ;
        RECT 89.720 200.985 89.890 201.815 ;
        RECT 90.060 201.225 90.390 201.985 ;
        RECT 90.560 200.985 90.730 201.815 ;
        RECT 91.045 200.985 92.255 202.075 ;
        RECT 18.280 200.815 92.340 200.985 ;
        RECT 18.365 199.725 19.575 200.815 ;
        RECT 19.745 200.380 25.090 200.815 ;
        RECT 18.365 199.015 18.885 199.555 ;
        RECT 19.055 199.185 19.575 199.725 ;
        RECT 18.365 198.265 19.575 199.015 ;
        RECT 21.330 198.810 21.670 199.640 ;
        RECT 23.150 199.130 23.500 200.380 ;
        RECT 25.265 199.725 27.855 200.815 ;
        RECT 25.265 199.035 26.475 199.555 ;
        RECT 26.645 199.205 27.855 199.725 ;
        RECT 28.085 199.675 28.295 200.815 ;
        RECT 28.465 199.665 28.795 200.645 ;
        RECT 28.965 199.675 29.195 200.815 ;
        RECT 29.405 199.725 31.075 200.815 ;
        RECT 19.745 198.265 25.090 198.810 ;
        RECT 25.265 198.265 27.855 199.035 ;
        RECT 28.085 198.265 28.295 199.085 ;
        RECT 28.465 199.065 28.715 199.665 ;
        RECT 28.885 199.255 29.215 199.505 ;
        RECT 28.465 198.435 28.795 199.065 ;
        RECT 28.965 198.265 29.195 199.085 ;
        RECT 29.405 199.035 30.155 199.555 ;
        RECT 30.325 199.205 31.075 199.725 ;
        RECT 31.245 199.650 31.535 200.815 ;
        RECT 31.705 199.725 32.915 200.815 ;
        RECT 33.175 200.145 33.345 200.645 ;
        RECT 33.515 200.315 33.845 200.815 ;
        RECT 33.175 199.975 33.840 200.145 ;
        RECT 29.405 198.265 31.075 199.035 ;
        RECT 31.705 199.015 32.225 199.555 ;
        RECT 32.395 199.185 32.915 199.725 ;
        RECT 33.090 199.155 33.440 199.805 ;
        RECT 31.245 198.265 31.535 198.990 ;
        RECT 31.705 198.265 32.915 199.015 ;
        RECT 33.610 198.985 33.840 199.975 ;
        RECT 33.175 198.815 33.840 198.985 ;
        RECT 33.175 198.525 33.345 198.815 ;
        RECT 33.515 198.265 33.845 198.645 ;
        RECT 34.015 198.525 34.200 200.645 ;
        RECT 34.440 200.355 34.705 200.815 ;
        RECT 34.875 200.220 35.125 200.645 ;
        RECT 35.335 200.370 36.440 200.540 ;
        RECT 34.820 200.090 35.125 200.220 ;
        RECT 34.370 198.895 34.650 199.845 ;
        RECT 34.820 198.985 34.990 200.090 ;
        RECT 35.160 199.305 35.400 199.900 ;
        RECT 35.570 199.835 36.100 200.200 ;
        RECT 35.570 199.135 35.740 199.835 ;
        RECT 36.270 199.755 36.440 200.370 ;
        RECT 36.610 200.015 36.780 200.815 ;
        RECT 36.950 200.315 37.200 200.645 ;
        RECT 37.425 200.345 38.310 200.515 ;
        RECT 36.270 199.665 36.780 199.755 ;
        RECT 34.820 198.855 35.045 198.985 ;
        RECT 35.215 198.915 35.740 199.135 ;
        RECT 35.910 199.495 36.780 199.665 ;
        RECT 34.455 198.265 34.705 198.725 ;
        RECT 34.875 198.715 35.045 198.855 ;
        RECT 35.910 198.715 36.080 199.495 ;
        RECT 36.610 199.425 36.780 199.495 ;
        RECT 36.290 199.245 36.490 199.275 ;
        RECT 36.950 199.245 37.120 200.315 ;
        RECT 37.290 199.425 37.480 200.145 ;
        RECT 36.290 198.945 37.120 199.245 ;
        RECT 37.650 199.215 37.970 200.175 ;
        RECT 34.875 198.545 35.210 198.715 ;
        RECT 35.405 198.545 36.080 198.715 ;
        RECT 36.400 198.265 36.770 198.765 ;
        RECT 36.950 198.715 37.120 198.945 ;
        RECT 37.505 198.885 37.970 199.215 ;
        RECT 38.140 199.505 38.310 200.345 ;
        RECT 38.490 200.315 38.805 200.815 ;
        RECT 39.035 200.085 39.375 200.645 ;
        RECT 38.480 199.710 39.375 200.085 ;
        RECT 39.545 199.805 39.715 200.815 ;
        RECT 39.185 199.505 39.375 199.710 ;
        RECT 39.885 199.755 40.215 200.600 ;
        RECT 39.885 199.675 40.275 199.755 ;
        RECT 40.445 199.725 43.035 200.815 ;
        RECT 40.060 199.625 40.275 199.675 ;
        RECT 38.140 199.175 39.015 199.505 ;
        RECT 39.185 199.175 39.935 199.505 ;
        RECT 38.140 198.715 38.310 199.175 ;
        RECT 39.185 199.005 39.385 199.175 ;
        RECT 40.105 199.045 40.275 199.625 ;
        RECT 40.050 199.005 40.275 199.045 ;
        RECT 36.950 198.545 37.355 198.715 ;
        RECT 37.525 198.545 38.310 198.715 ;
        RECT 38.585 198.265 38.795 198.795 ;
        RECT 39.055 198.480 39.385 199.005 ;
        RECT 39.895 198.920 40.275 199.005 ;
        RECT 40.445 199.035 41.655 199.555 ;
        RECT 41.825 199.205 43.035 199.725 ;
        RECT 39.555 198.265 39.725 198.875 ;
        RECT 39.895 198.485 40.225 198.920 ;
        RECT 40.445 198.265 43.035 199.035 ;
        RECT 43.220 198.445 43.500 200.635 ;
        RECT 43.690 199.675 43.975 200.815 ;
        RECT 44.240 200.165 44.410 200.635 ;
        RECT 44.585 200.335 44.915 200.815 ;
        RECT 45.085 200.165 45.265 200.635 ;
        RECT 44.240 199.965 45.265 200.165 ;
        RECT 43.700 198.995 43.960 199.505 ;
        RECT 44.170 199.175 44.430 199.795 ;
        RECT 44.625 199.175 45.050 199.795 ;
        RECT 45.435 199.525 45.765 200.635 ;
        RECT 45.935 200.405 46.285 200.815 ;
        RECT 46.455 200.225 46.695 200.615 ;
        RECT 45.220 199.225 45.765 199.525 ;
        RECT 45.945 200.025 46.695 200.225 ;
        RECT 45.945 199.345 46.285 200.025 ;
        RECT 45.220 198.995 45.440 199.225 ;
        RECT 43.700 198.805 45.440 198.995 ;
        RECT 43.700 198.265 44.430 198.635 ;
        RECT 45.010 198.445 45.440 198.805 ;
        RECT 45.610 198.265 45.855 199.045 ;
        RECT 46.055 198.445 46.285 199.345 ;
        RECT 46.465 198.505 46.695 199.845 ;
        RECT 46.885 199.675 47.160 200.645 ;
        RECT 47.370 200.015 47.650 200.815 ;
        RECT 47.820 200.305 49.435 200.635 ;
        RECT 47.820 199.965 48.995 200.135 ;
        RECT 47.820 199.845 47.990 199.965 ;
        RECT 47.330 199.675 47.990 199.845 ;
        RECT 46.885 198.940 47.055 199.675 ;
        RECT 47.330 199.505 47.500 199.675 ;
        RECT 48.250 199.505 48.495 199.795 ;
        RECT 48.665 199.675 48.995 199.965 ;
        RECT 49.255 199.505 49.425 200.065 ;
        RECT 49.675 199.675 49.935 200.815 ;
        RECT 50.105 200.380 55.450 200.815 ;
        RECT 47.225 199.175 47.500 199.505 ;
        RECT 47.670 199.175 48.495 199.505 ;
        RECT 48.710 199.175 49.425 199.505 ;
        RECT 49.595 199.255 49.930 199.505 ;
        RECT 47.330 199.005 47.500 199.175 ;
        RECT 49.175 199.085 49.425 199.175 ;
        RECT 46.885 198.595 47.160 198.940 ;
        RECT 47.330 198.835 48.995 199.005 ;
        RECT 47.350 198.265 47.725 198.665 ;
        RECT 47.895 198.485 48.065 198.835 ;
        RECT 48.235 198.265 48.565 198.665 ;
        RECT 48.735 198.435 48.995 198.835 ;
        RECT 49.175 198.665 49.505 199.085 ;
        RECT 49.675 198.265 49.935 199.085 ;
        RECT 51.690 198.810 52.030 199.640 ;
        RECT 53.510 199.130 53.860 200.380 ;
        RECT 55.625 199.725 56.835 200.815 ;
        RECT 55.625 199.015 56.145 199.555 ;
        RECT 56.315 199.185 56.835 199.725 ;
        RECT 57.005 199.650 57.295 200.815 ;
        RECT 50.105 198.265 55.450 198.810 ;
        RECT 55.625 198.265 56.835 199.015 ;
        RECT 57.005 198.265 57.295 198.990 ;
        RECT 57.480 198.445 57.760 200.635 ;
        RECT 57.950 199.675 58.235 200.815 ;
        RECT 58.500 200.165 58.670 200.635 ;
        RECT 58.845 200.335 59.175 200.815 ;
        RECT 59.345 200.165 59.525 200.635 ;
        RECT 58.500 199.965 59.525 200.165 ;
        RECT 57.960 198.995 58.220 199.505 ;
        RECT 58.430 199.175 58.690 199.795 ;
        RECT 58.885 199.175 59.310 199.795 ;
        RECT 59.695 199.525 60.025 200.635 ;
        RECT 60.195 200.405 60.545 200.815 ;
        RECT 60.715 200.225 60.955 200.615 ;
        RECT 59.480 199.225 60.025 199.525 ;
        RECT 60.205 200.025 60.955 200.225 ;
        RECT 60.205 199.345 60.545 200.025 ;
        RECT 59.480 198.995 59.700 199.225 ;
        RECT 57.960 198.805 59.700 198.995 ;
        RECT 57.960 198.265 58.690 198.635 ;
        RECT 59.270 198.445 59.700 198.805 ;
        RECT 59.870 198.265 60.115 199.045 ;
        RECT 60.315 198.445 60.545 199.345 ;
        RECT 60.725 198.505 60.955 199.845 ;
        RECT 61.145 199.725 62.815 200.815 ;
        RECT 63.465 200.225 63.705 200.615 ;
        RECT 63.875 200.405 64.225 200.815 ;
        RECT 63.465 200.025 64.215 200.225 ;
        RECT 61.145 199.035 61.895 199.555 ;
        RECT 62.065 199.205 62.815 199.725 ;
        RECT 61.145 198.265 62.815 199.035 ;
        RECT 63.465 198.505 63.695 199.845 ;
        RECT 63.875 199.345 64.215 200.025 ;
        RECT 64.395 199.525 64.725 200.635 ;
        RECT 64.895 200.165 65.075 200.635 ;
        RECT 65.245 200.335 65.575 200.815 ;
        RECT 65.750 200.165 65.920 200.635 ;
        RECT 64.895 199.965 65.920 200.165 ;
        RECT 63.875 198.445 64.105 199.345 ;
        RECT 64.395 199.225 64.940 199.525 ;
        RECT 64.305 198.265 64.550 199.045 ;
        RECT 64.720 198.995 64.940 199.225 ;
        RECT 65.110 199.175 65.535 199.795 ;
        RECT 65.730 199.175 65.990 199.795 ;
        RECT 66.185 199.675 66.470 200.815 ;
        RECT 66.200 198.995 66.460 199.505 ;
        RECT 64.720 198.805 66.460 198.995 ;
        RECT 64.720 198.445 65.150 198.805 ;
        RECT 65.730 198.265 66.460 198.635 ;
        RECT 66.660 198.445 66.940 200.635 ;
        RECT 67.125 199.725 70.635 200.815 ;
        RECT 70.805 199.725 72.015 200.815 ;
        RECT 72.205 200.225 72.445 200.615 ;
        RECT 72.615 200.405 72.965 200.815 ;
        RECT 72.205 200.025 72.955 200.225 ;
        RECT 67.125 199.035 68.775 199.555 ;
        RECT 68.945 199.205 70.635 199.725 ;
        RECT 67.125 198.265 70.635 199.035 ;
        RECT 70.805 199.015 71.325 199.555 ;
        RECT 71.495 199.185 72.015 199.725 ;
        RECT 70.805 198.265 72.015 199.015 ;
        RECT 72.205 198.505 72.435 199.845 ;
        RECT 72.615 199.345 72.955 200.025 ;
        RECT 73.135 199.525 73.465 200.635 ;
        RECT 73.635 200.165 73.815 200.635 ;
        RECT 73.985 200.335 74.315 200.815 ;
        RECT 74.490 200.165 74.660 200.635 ;
        RECT 73.635 199.965 74.660 200.165 ;
        RECT 72.615 198.445 72.845 199.345 ;
        RECT 73.135 199.225 73.680 199.525 ;
        RECT 73.045 198.265 73.290 199.045 ;
        RECT 73.460 198.995 73.680 199.225 ;
        RECT 73.850 199.175 74.275 199.795 ;
        RECT 74.470 199.175 74.730 199.795 ;
        RECT 74.925 199.675 75.210 200.815 ;
        RECT 74.940 198.995 75.200 199.505 ;
        RECT 73.460 198.805 75.200 198.995 ;
        RECT 73.460 198.445 73.890 198.805 ;
        RECT 74.470 198.265 75.200 198.635 ;
        RECT 75.400 198.445 75.680 200.635 ;
        RECT 75.865 199.725 79.375 200.815 ;
        RECT 75.865 199.035 77.515 199.555 ;
        RECT 77.685 199.205 79.375 199.725 ;
        RECT 80.475 199.675 80.805 200.815 ;
        RECT 81.335 199.845 81.665 200.630 ;
        RECT 80.985 199.675 81.665 199.845 ;
        RECT 80.465 199.255 80.815 199.505 ;
        RECT 80.985 199.075 81.155 199.675 ;
        RECT 82.765 199.650 83.055 200.815 ;
        RECT 83.235 199.865 83.510 200.635 ;
        RECT 83.680 200.205 84.010 200.635 ;
        RECT 84.180 200.375 84.375 200.815 ;
        RECT 84.555 200.205 84.885 200.635 ;
        RECT 83.680 200.035 84.885 200.205 ;
        RECT 83.235 199.675 83.820 199.865 ;
        RECT 83.990 199.705 84.885 200.035 ;
        RECT 81.325 199.255 81.675 199.505 ;
        RECT 75.865 198.265 79.375 199.035 ;
        RECT 80.475 198.265 80.745 199.075 ;
        RECT 80.915 198.435 81.245 199.075 ;
        RECT 81.415 198.265 81.655 199.075 ;
        RECT 82.765 198.265 83.055 198.990 ;
        RECT 83.235 198.855 83.475 199.505 ;
        RECT 83.645 199.005 83.820 199.675 ;
        RECT 85.985 199.675 86.370 200.645 ;
        RECT 86.540 200.355 86.865 200.815 ;
        RECT 87.385 200.185 87.665 200.645 ;
        RECT 86.540 199.965 87.665 200.185 ;
        RECT 83.990 199.175 84.405 199.505 ;
        RECT 84.585 199.175 84.880 199.505 ;
        RECT 83.645 198.825 83.975 199.005 ;
        RECT 83.250 198.265 83.580 198.655 ;
        RECT 83.750 198.445 83.975 198.825 ;
        RECT 84.175 198.555 84.405 199.175 ;
        RECT 85.985 199.005 86.265 199.675 ;
        RECT 86.540 199.505 86.990 199.965 ;
        RECT 87.855 199.795 88.255 200.645 ;
        RECT 88.655 200.355 88.925 200.815 ;
        RECT 89.095 200.185 89.380 200.645 ;
        RECT 86.435 199.175 86.990 199.505 ;
        RECT 87.160 199.235 88.255 199.795 ;
        RECT 86.540 199.065 86.990 199.175 ;
        RECT 84.585 198.265 84.885 198.995 ;
        RECT 85.985 198.435 86.370 199.005 ;
        RECT 86.540 198.895 87.665 199.065 ;
        RECT 86.540 198.265 86.865 198.725 ;
        RECT 87.385 198.435 87.665 198.895 ;
        RECT 87.855 198.435 88.255 199.235 ;
        RECT 88.425 199.965 89.380 200.185 ;
        RECT 88.425 199.065 88.635 199.965 ;
        RECT 88.805 199.235 89.495 199.795 ;
        RECT 89.665 199.725 90.875 200.815 ;
        RECT 88.425 198.895 89.380 199.065 ;
        RECT 88.655 198.265 88.925 198.725 ;
        RECT 89.095 198.435 89.380 198.895 ;
        RECT 89.665 199.015 90.185 199.555 ;
        RECT 90.355 199.185 90.875 199.725 ;
        RECT 91.045 199.725 92.255 200.815 ;
        RECT 91.045 199.185 91.565 199.725 ;
        RECT 91.735 199.015 92.255 199.555 ;
        RECT 89.665 198.265 90.875 199.015 ;
        RECT 91.045 198.265 92.255 199.015 ;
        RECT 18.280 198.095 92.340 198.265 ;
        RECT 18.365 197.345 19.575 198.095 ;
        RECT 19.745 197.550 25.090 198.095 ;
        RECT 25.265 197.550 30.610 198.095 ;
        RECT 30.785 197.550 36.130 198.095 ;
        RECT 36.305 197.550 41.650 198.095 ;
        RECT 18.365 196.805 18.885 197.345 ;
        RECT 19.055 196.635 19.575 197.175 ;
        RECT 21.330 196.720 21.670 197.550 ;
        RECT 18.365 195.545 19.575 196.635 ;
        RECT 23.150 195.980 23.500 197.230 ;
        RECT 26.850 196.720 27.190 197.550 ;
        RECT 28.670 195.980 29.020 197.230 ;
        RECT 32.370 196.720 32.710 197.550 ;
        RECT 34.190 195.980 34.540 197.230 ;
        RECT 37.890 196.720 38.230 197.550 ;
        RECT 41.825 197.325 43.495 198.095 ;
        RECT 44.125 197.370 44.415 198.095 ;
        RECT 44.585 197.325 47.175 198.095 ;
        RECT 39.710 195.980 40.060 197.230 ;
        RECT 41.825 196.805 42.575 197.325 ;
        RECT 42.745 196.635 43.495 197.155 ;
        RECT 44.585 196.805 45.795 197.325 ;
        RECT 47.845 197.275 48.075 198.095 ;
        RECT 48.245 197.295 48.575 197.925 ;
        RECT 19.745 195.545 25.090 195.980 ;
        RECT 25.265 195.545 30.610 195.980 ;
        RECT 30.785 195.545 36.130 195.980 ;
        RECT 36.305 195.545 41.650 195.980 ;
        RECT 41.825 195.545 43.495 196.635 ;
        RECT 44.125 195.545 44.415 196.710 ;
        RECT 45.965 196.635 47.175 197.155 ;
        RECT 47.825 196.855 48.155 197.105 ;
        RECT 48.325 196.695 48.575 197.295 ;
        RECT 48.745 197.275 48.955 198.095 ;
        RECT 49.185 197.325 52.695 198.095 ;
        RECT 49.185 196.805 50.835 197.325 ;
        RECT 44.585 195.545 47.175 196.635 ;
        RECT 47.845 195.545 48.075 196.685 ;
        RECT 48.245 195.715 48.575 196.695 ;
        RECT 48.745 195.545 48.955 196.685 ;
        RECT 51.005 196.635 52.695 197.155 ;
        RECT 49.185 195.545 52.695 196.635 ;
        RECT 53.340 195.725 53.620 197.915 ;
        RECT 53.820 197.725 54.550 198.095 ;
        RECT 55.130 197.555 55.560 197.915 ;
        RECT 53.820 197.365 55.560 197.555 ;
        RECT 53.820 196.855 54.080 197.365 ;
        RECT 53.810 195.545 54.095 196.685 ;
        RECT 54.290 196.565 54.550 197.185 ;
        RECT 54.745 196.565 55.170 197.185 ;
        RECT 55.340 197.135 55.560 197.365 ;
        RECT 55.730 197.315 55.975 198.095 ;
        RECT 55.340 196.835 55.885 197.135 ;
        RECT 56.175 197.015 56.405 197.915 ;
        RECT 54.360 196.195 55.385 196.395 ;
        RECT 54.360 195.725 54.530 196.195 ;
        RECT 54.705 195.545 55.035 196.025 ;
        RECT 55.205 195.725 55.385 196.195 ;
        RECT 55.555 195.725 55.885 196.835 ;
        RECT 56.065 196.335 56.405 197.015 ;
        RECT 56.585 196.515 56.815 197.855 ;
        RECT 57.005 197.420 57.280 197.765 ;
        RECT 57.470 197.695 57.845 198.095 ;
        RECT 58.015 197.525 58.185 197.875 ;
        RECT 58.355 197.695 58.685 198.095 ;
        RECT 58.855 197.525 59.115 197.925 ;
        RECT 57.005 196.685 57.175 197.420 ;
        RECT 57.450 197.355 59.115 197.525 ;
        RECT 57.450 197.185 57.620 197.355 ;
        RECT 59.295 197.275 59.625 197.695 ;
        RECT 59.795 197.275 60.055 198.095 ;
        RECT 60.225 197.325 63.735 198.095 ;
        RECT 59.295 197.185 59.545 197.275 ;
        RECT 57.345 196.855 57.620 197.185 ;
        RECT 57.790 196.855 58.615 197.185 ;
        RECT 58.830 196.855 59.545 197.185 ;
        RECT 59.715 196.855 60.050 197.105 ;
        RECT 57.450 196.685 57.620 196.855 ;
        RECT 56.065 196.135 56.815 196.335 ;
        RECT 56.055 195.545 56.405 195.955 ;
        RECT 56.575 195.745 56.815 196.135 ;
        RECT 57.005 195.715 57.280 196.685 ;
        RECT 57.450 196.515 58.110 196.685 ;
        RECT 58.370 196.565 58.615 196.855 ;
        RECT 57.940 196.395 58.110 196.515 ;
        RECT 58.785 196.395 59.115 196.685 ;
        RECT 57.490 195.545 57.770 196.345 ;
        RECT 57.940 196.225 59.115 196.395 ;
        RECT 59.375 196.295 59.545 196.855 ;
        RECT 60.225 196.805 61.875 197.325 ;
        RECT 57.940 195.725 59.555 196.055 ;
        RECT 59.795 195.545 60.055 196.685 ;
        RECT 62.045 196.635 63.735 197.155 ;
        RECT 60.225 195.545 63.735 196.635 ;
        RECT 63.920 195.725 64.200 197.915 ;
        RECT 64.400 197.725 65.130 198.095 ;
        RECT 65.710 197.555 66.140 197.915 ;
        RECT 64.400 197.365 66.140 197.555 ;
        RECT 64.400 196.855 64.660 197.365 ;
        RECT 64.390 195.545 64.675 196.685 ;
        RECT 64.870 196.565 65.130 197.185 ;
        RECT 65.325 196.565 65.750 197.185 ;
        RECT 65.920 197.135 66.140 197.365 ;
        RECT 66.310 197.315 66.555 198.095 ;
        RECT 65.920 196.835 66.465 197.135 ;
        RECT 66.755 197.015 66.985 197.915 ;
        RECT 64.940 196.195 65.965 196.395 ;
        RECT 64.940 195.725 65.110 196.195 ;
        RECT 65.285 195.545 65.615 196.025 ;
        RECT 65.785 195.725 65.965 196.195 ;
        RECT 66.135 195.725 66.465 196.835 ;
        RECT 66.645 196.335 66.985 197.015 ;
        RECT 67.165 196.515 67.395 197.855 ;
        RECT 67.585 197.325 69.255 198.095 ;
        RECT 69.885 197.370 70.175 198.095 ;
        RECT 70.345 197.345 71.555 198.095 ;
        RECT 67.585 196.805 68.335 197.325 ;
        RECT 68.505 196.635 69.255 197.155 ;
        RECT 70.345 196.805 70.865 197.345 ;
        RECT 66.645 196.135 67.395 196.335 ;
        RECT 66.635 195.545 66.985 195.955 ;
        RECT 67.155 195.745 67.395 196.135 ;
        RECT 67.585 195.545 69.255 196.635 ;
        RECT 69.885 195.545 70.175 196.710 ;
        RECT 71.035 196.635 71.555 197.175 ;
        RECT 70.345 195.545 71.555 196.635 ;
        RECT 71.745 196.515 71.975 197.855 ;
        RECT 72.155 197.015 72.385 197.915 ;
        RECT 72.585 197.315 72.830 198.095 ;
        RECT 73.000 197.555 73.430 197.915 ;
        RECT 74.010 197.725 74.740 198.095 ;
        RECT 73.000 197.365 74.740 197.555 ;
        RECT 73.000 197.135 73.220 197.365 ;
        RECT 72.155 196.335 72.495 197.015 ;
        RECT 71.745 196.135 72.495 196.335 ;
        RECT 72.675 196.835 73.220 197.135 ;
        RECT 71.745 195.745 71.985 196.135 ;
        RECT 72.155 195.545 72.505 195.955 ;
        RECT 72.675 195.725 73.005 196.835 ;
        RECT 73.390 196.565 73.815 197.185 ;
        RECT 74.010 196.565 74.270 197.185 ;
        RECT 74.480 196.855 74.740 197.365 ;
        RECT 73.175 196.195 74.200 196.395 ;
        RECT 73.175 195.725 73.355 196.195 ;
        RECT 73.525 195.545 73.855 196.025 ;
        RECT 74.030 195.725 74.200 196.195 ;
        RECT 74.465 195.545 74.750 196.685 ;
        RECT 74.940 195.725 75.220 197.915 ;
        RECT 75.405 197.325 78.915 198.095 ;
        RECT 80.010 197.565 80.300 197.915 ;
        RECT 80.495 197.735 80.825 198.095 ;
        RECT 80.995 197.565 81.225 197.870 ;
        RECT 80.010 197.395 81.225 197.565 ;
        RECT 81.415 197.755 81.585 197.790 ;
        RECT 81.415 197.585 81.615 197.755 ;
        RECT 75.405 196.805 77.055 197.325 ;
        RECT 81.415 197.225 81.585 197.585 ;
        RECT 82.050 197.315 82.550 197.925 ;
        RECT 77.225 196.635 78.915 197.155 ;
        RECT 80.070 197.075 80.330 197.185 ;
        RECT 80.065 196.905 80.330 197.075 ;
        RECT 80.070 196.855 80.330 196.905 ;
        RECT 80.510 196.855 80.895 197.185 ;
        RECT 81.065 197.055 81.585 197.225 ;
        RECT 75.405 195.545 78.915 196.635 ;
        RECT 80.010 195.545 80.330 196.685 ;
        RECT 80.510 195.805 80.705 196.855 ;
        RECT 81.065 196.675 81.235 197.055 ;
        RECT 80.885 196.395 81.235 196.675 ;
        RECT 81.425 196.525 81.670 196.885 ;
        RECT 81.845 196.855 82.195 197.105 ;
        RECT 82.380 196.685 82.550 197.315 ;
        RECT 83.180 197.445 83.510 197.925 ;
        RECT 83.680 197.635 83.905 198.095 ;
        RECT 84.075 197.445 84.405 197.925 ;
        RECT 83.180 197.275 84.405 197.445 ;
        RECT 84.595 197.295 84.845 198.095 ;
        RECT 85.015 197.295 85.355 197.925 ;
        RECT 82.720 196.905 83.050 197.105 ;
        RECT 83.220 196.905 83.550 197.105 ;
        RECT 83.720 196.905 84.140 197.105 ;
        RECT 84.315 196.935 85.010 197.105 ;
        RECT 84.315 196.685 84.485 196.935 ;
        RECT 85.180 196.685 85.355 197.295 ;
        RECT 85.725 197.465 86.055 197.825 ;
        RECT 86.675 197.635 86.925 198.095 ;
        RECT 87.095 197.635 87.655 197.925 ;
        RECT 85.725 197.275 87.115 197.465 ;
        RECT 86.945 197.185 87.115 197.275 ;
        RECT 82.050 196.515 84.485 196.685 ;
        RECT 80.885 195.715 81.215 196.395 ;
        RECT 81.415 195.545 81.670 196.345 ;
        RECT 82.050 195.715 82.380 196.515 ;
        RECT 82.550 195.545 82.880 196.345 ;
        RECT 83.180 195.715 83.510 196.515 ;
        RECT 84.155 195.545 84.405 196.345 ;
        RECT 84.675 195.545 84.845 196.685 ;
        RECT 85.015 195.715 85.355 196.685 ;
        RECT 85.540 196.855 86.215 197.105 ;
        RECT 86.435 196.855 86.775 197.105 ;
        RECT 86.945 196.855 87.235 197.185 ;
        RECT 85.540 196.495 85.805 196.855 ;
        RECT 86.945 196.605 87.115 196.855 ;
        RECT 86.175 196.435 87.115 196.605 ;
        RECT 85.725 195.545 86.005 196.215 ;
        RECT 86.175 195.885 86.475 196.435 ;
        RECT 87.405 196.265 87.655 197.635 ;
        RECT 87.825 197.325 90.415 198.095 ;
        RECT 91.045 197.345 92.255 198.095 ;
        RECT 87.825 196.805 89.035 197.325 ;
        RECT 89.205 196.635 90.415 197.155 ;
        RECT 86.675 195.545 87.005 196.265 ;
        RECT 87.195 195.715 87.655 196.265 ;
        RECT 87.825 195.545 90.415 196.635 ;
        RECT 91.045 196.635 91.565 197.175 ;
        RECT 91.735 196.805 92.255 197.345 ;
        RECT 91.045 195.545 92.255 196.635 ;
        RECT 18.280 195.375 92.340 195.545 ;
        RECT 18.365 194.285 19.575 195.375 ;
        RECT 19.745 194.940 25.090 195.375 ;
        RECT 25.265 194.940 30.610 195.375 ;
        RECT 18.365 193.575 18.885 194.115 ;
        RECT 19.055 193.745 19.575 194.285 ;
        RECT 18.365 192.825 19.575 193.575 ;
        RECT 21.330 193.370 21.670 194.200 ;
        RECT 23.150 193.690 23.500 194.940 ;
        RECT 26.850 193.370 27.190 194.200 ;
        RECT 28.670 193.690 29.020 194.940 ;
        RECT 31.245 194.210 31.535 195.375 ;
        RECT 32.715 194.705 32.885 195.205 ;
        RECT 33.055 194.875 33.385 195.375 ;
        RECT 32.715 194.535 33.380 194.705 ;
        RECT 32.630 193.715 32.980 194.365 ;
        RECT 19.745 192.825 25.090 193.370 ;
        RECT 25.265 192.825 30.610 193.370 ;
        RECT 31.245 192.825 31.535 193.550 ;
        RECT 33.150 193.545 33.380 194.535 ;
        RECT 32.715 193.375 33.380 193.545 ;
        RECT 32.715 193.085 32.885 193.375 ;
        RECT 33.055 192.825 33.385 193.205 ;
        RECT 33.555 193.085 33.740 195.205 ;
        RECT 33.980 194.915 34.245 195.375 ;
        RECT 34.415 194.780 34.665 195.205 ;
        RECT 34.875 194.930 35.980 195.100 ;
        RECT 34.360 194.650 34.665 194.780 ;
        RECT 33.910 193.455 34.190 194.405 ;
        RECT 34.360 193.545 34.530 194.650 ;
        RECT 34.700 193.865 34.940 194.460 ;
        RECT 35.110 194.395 35.640 194.760 ;
        RECT 35.110 193.695 35.280 194.395 ;
        RECT 35.810 194.315 35.980 194.930 ;
        RECT 36.150 194.575 36.320 195.375 ;
        RECT 36.490 194.875 36.740 195.205 ;
        RECT 36.965 194.905 37.850 195.075 ;
        RECT 35.810 194.225 36.320 194.315 ;
        RECT 34.360 193.415 34.585 193.545 ;
        RECT 34.755 193.475 35.280 193.695 ;
        RECT 35.450 194.055 36.320 194.225 ;
        RECT 33.995 192.825 34.245 193.285 ;
        RECT 34.415 193.275 34.585 193.415 ;
        RECT 35.450 193.275 35.620 194.055 ;
        RECT 36.150 193.985 36.320 194.055 ;
        RECT 35.830 193.805 36.030 193.835 ;
        RECT 36.490 193.805 36.660 194.875 ;
        RECT 36.830 193.985 37.020 194.705 ;
        RECT 35.830 193.505 36.660 193.805 ;
        RECT 37.190 193.775 37.510 194.735 ;
        RECT 34.415 193.105 34.750 193.275 ;
        RECT 34.945 193.105 35.620 193.275 ;
        RECT 35.940 192.825 36.310 193.325 ;
        RECT 36.490 193.275 36.660 193.505 ;
        RECT 37.045 193.445 37.510 193.775 ;
        RECT 37.680 194.065 37.850 194.905 ;
        RECT 38.030 194.875 38.345 195.375 ;
        RECT 38.575 194.645 38.915 195.205 ;
        RECT 38.020 194.270 38.915 194.645 ;
        RECT 39.085 194.365 39.255 195.375 ;
        RECT 38.725 194.065 38.915 194.270 ;
        RECT 39.425 194.315 39.755 195.160 ;
        RECT 39.425 194.235 39.815 194.315 ;
        RECT 39.985 194.285 41.655 195.375 ;
        RECT 39.600 194.185 39.815 194.235 ;
        RECT 37.680 193.735 38.555 194.065 ;
        RECT 38.725 193.735 39.475 194.065 ;
        RECT 37.680 193.275 37.850 193.735 ;
        RECT 38.725 193.565 38.925 193.735 ;
        RECT 39.645 193.605 39.815 194.185 ;
        RECT 39.590 193.565 39.815 193.605 ;
        RECT 36.490 193.105 36.895 193.275 ;
        RECT 37.065 193.105 37.850 193.275 ;
        RECT 38.125 192.825 38.335 193.355 ;
        RECT 38.595 193.040 38.925 193.565 ;
        RECT 39.435 193.480 39.815 193.565 ;
        RECT 39.985 193.595 40.735 194.115 ;
        RECT 40.905 193.765 41.655 194.285 ;
        RECT 41.830 194.235 42.085 195.375 ;
        RECT 42.280 194.825 43.475 195.155 ;
        RECT 42.335 194.065 42.505 194.625 ;
        RECT 42.730 194.405 43.150 194.655 ;
        RECT 43.655 194.575 43.935 195.375 ;
        RECT 42.730 194.235 43.975 194.405 ;
        RECT 44.145 194.235 44.415 195.205 ;
        RECT 44.675 194.755 44.845 195.185 ;
        RECT 45.015 194.925 45.345 195.375 ;
        RECT 44.675 194.525 45.350 194.755 ;
        RECT 43.805 194.065 43.975 194.235 ;
        RECT 41.830 193.815 42.165 194.065 ;
        RECT 42.335 193.735 43.075 194.065 ;
        RECT 43.805 193.735 44.035 194.065 ;
        RECT 42.335 193.645 42.585 193.735 ;
        RECT 39.095 192.825 39.265 193.435 ;
        RECT 39.435 193.045 39.765 193.480 ;
        RECT 39.985 192.825 41.655 193.595 ;
        RECT 41.850 193.475 42.585 193.645 ;
        RECT 43.805 193.565 43.975 193.735 ;
        RECT 41.850 193.005 42.160 193.475 ;
        RECT 43.235 193.395 43.975 193.565 ;
        RECT 44.245 193.500 44.415 194.235 ;
        RECT 44.645 193.505 44.945 194.355 ;
        RECT 45.115 193.875 45.350 194.525 ;
        RECT 45.520 194.215 45.805 195.160 ;
        RECT 45.985 194.905 46.670 195.375 ;
        RECT 45.980 194.385 46.675 194.695 ;
        RECT 46.850 194.320 47.155 195.105 ;
        RECT 45.520 194.065 46.380 194.215 ;
        RECT 45.520 194.045 46.805 194.065 ;
        RECT 45.115 193.545 45.650 193.875 ;
        RECT 45.820 193.685 46.805 194.045 ;
        RECT 42.330 192.825 43.065 193.305 ;
        RECT 43.235 193.045 43.405 193.395 ;
        RECT 43.575 192.825 43.955 193.225 ;
        RECT 44.145 193.155 44.415 193.500 ;
        RECT 45.115 193.395 45.335 193.545 ;
        RECT 44.590 192.825 44.925 193.330 ;
        RECT 45.095 193.020 45.335 193.395 ;
        RECT 45.820 193.350 45.990 193.685 ;
        RECT 46.980 193.515 47.155 194.320 ;
        RECT 48.325 194.315 48.655 195.160 ;
        RECT 48.825 194.365 48.995 195.375 ;
        RECT 49.165 194.645 49.505 195.205 ;
        RECT 49.735 194.875 50.050 195.375 ;
        RECT 50.230 194.905 51.115 195.075 ;
        RECT 45.615 193.155 45.990 193.350 ;
        RECT 45.615 193.010 45.785 193.155 ;
        RECT 46.350 192.825 46.745 193.320 ;
        RECT 46.915 192.995 47.155 193.515 ;
        RECT 48.265 194.235 48.655 194.315 ;
        RECT 49.165 194.270 50.060 194.645 ;
        RECT 48.265 194.185 48.480 194.235 ;
        RECT 48.265 193.605 48.435 194.185 ;
        RECT 49.165 194.065 49.355 194.270 ;
        RECT 50.230 194.065 50.400 194.905 ;
        RECT 51.340 194.875 51.590 195.205 ;
        RECT 48.605 193.735 49.355 194.065 ;
        RECT 49.525 193.735 50.400 194.065 ;
        RECT 48.265 193.565 48.490 193.605 ;
        RECT 49.155 193.565 49.355 193.735 ;
        RECT 48.265 193.480 48.645 193.565 ;
        RECT 48.315 193.045 48.645 193.480 ;
        RECT 48.815 192.825 48.985 193.435 ;
        RECT 49.155 193.040 49.485 193.565 ;
        RECT 49.745 192.825 49.955 193.355 ;
        RECT 50.230 193.275 50.400 193.735 ;
        RECT 50.570 193.775 50.890 194.735 ;
        RECT 51.060 193.985 51.250 194.705 ;
        RECT 51.420 193.805 51.590 194.875 ;
        RECT 51.760 194.575 51.930 195.375 ;
        RECT 52.100 194.930 53.205 195.100 ;
        RECT 52.100 194.315 52.270 194.930 ;
        RECT 53.415 194.780 53.665 195.205 ;
        RECT 53.835 194.915 54.100 195.375 ;
        RECT 52.440 194.395 52.970 194.760 ;
        RECT 53.415 194.650 53.720 194.780 ;
        RECT 51.760 194.225 52.270 194.315 ;
        RECT 51.760 194.055 52.630 194.225 ;
        RECT 51.760 193.985 51.930 194.055 ;
        RECT 52.050 193.805 52.250 193.835 ;
        RECT 50.570 193.445 51.035 193.775 ;
        RECT 51.420 193.505 52.250 193.805 ;
        RECT 51.420 193.275 51.590 193.505 ;
        RECT 50.230 193.105 51.015 193.275 ;
        RECT 51.185 193.105 51.590 193.275 ;
        RECT 51.770 192.825 52.140 193.325 ;
        RECT 52.460 193.275 52.630 194.055 ;
        RECT 52.800 193.695 52.970 194.395 ;
        RECT 53.140 193.865 53.380 194.460 ;
        RECT 52.800 193.475 53.325 193.695 ;
        RECT 53.550 193.545 53.720 194.650 ;
        RECT 53.495 193.415 53.720 193.545 ;
        RECT 53.890 193.455 54.170 194.405 ;
        RECT 53.495 193.275 53.665 193.415 ;
        RECT 52.460 193.105 53.135 193.275 ;
        RECT 53.330 193.105 53.665 193.275 ;
        RECT 53.835 192.825 54.085 193.285 ;
        RECT 54.340 193.085 54.525 195.205 ;
        RECT 54.695 194.875 55.025 195.375 ;
        RECT 55.195 194.705 55.365 195.205 ;
        RECT 54.700 194.535 55.365 194.705 ;
        RECT 54.700 193.545 54.930 194.535 ;
        RECT 55.100 193.715 55.450 194.365 ;
        RECT 55.625 194.285 56.835 195.375 ;
        RECT 55.625 193.575 56.145 194.115 ;
        RECT 56.315 193.745 56.835 194.285 ;
        RECT 57.005 194.210 57.295 195.375 ;
        RECT 57.465 194.285 58.675 195.375 ;
        RECT 57.465 193.575 57.985 194.115 ;
        RECT 58.155 193.745 58.675 194.285 ;
        RECT 58.905 194.235 59.115 195.375 ;
        RECT 59.285 194.225 59.615 195.205 ;
        RECT 59.785 194.235 60.015 195.375 ;
        RECT 60.285 194.315 60.615 195.160 ;
        RECT 60.785 194.365 60.955 195.375 ;
        RECT 61.125 194.645 61.465 195.205 ;
        RECT 61.695 194.875 62.010 195.375 ;
        RECT 62.190 194.905 63.075 195.075 ;
        RECT 60.225 194.235 60.615 194.315 ;
        RECT 61.125 194.270 62.020 194.645 ;
        RECT 54.700 193.375 55.365 193.545 ;
        RECT 54.695 192.825 55.025 193.205 ;
        RECT 55.195 193.085 55.365 193.375 ;
        RECT 55.625 192.825 56.835 193.575 ;
        RECT 57.005 192.825 57.295 193.550 ;
        RECT 57.465 192.825 58.675 193.575 ;
        RECT 58.905 192.825 59.115 193.645 ;
        RECT 59.285 193.625 59.535 194.225 ;
        RECT 60.225 194.185 60.440 194.235 ;
        RECT 59.705 193.815 60.035 194.065 ;
        RECT 59.285 192.995 59.615 193.625 ;
        RECT 59.785 192.825 60.015 193.645 ;
        RECT 60.225 193.605 60.395 194.185 ;
        RECT 61.125 194.065 61.315 194.270 ;
        RECT 62.190 194.065 62.360 194.905 ;
        RECT 63.300 194.875 63.550 195.205 ;
        RECT 60.565 193.735 61.315 194.065 ;
        RECT 61.485 193.735 62.360 194.065 ;
        RECT 60.225 193.565 60.450 193.605 ;
        RECT 61.115 193.565 61.315 193.735 ;
        RECT 60.225 193.480 60.605 193.565 ;
        RECT 60.275 193.045 60.605 193.480 ;
        RECT 60.775 192.825 60.945 193.435 ;
        RECT 61.115 193.040 61.445 193.565 ;
        RECT 61.705 192.825 61.915 193.355 ;
        RECT 62.190 193.275 62.360 193.735 ;
        RECT 62.530 193.775 62.850 194.735 ;
        RECT 63.020 193.985 63.210 194.705 ;
        RECT 63.380 193.805 63.550 194.875 ;
        RECT 63.720 194.575 63.890 195.375 ;
        RECT 64.060 194.930 65.165 195.100 ;
        RECT 64.060 194.315 64.230 194.930 ;
        RECT 65.375 194.780 65.625 195.205 ;
        RECT 65.795 194.915 66.060 195.375 ;
        RECT 64.400 194.395 64.930 194.760 ;
        RECT 65.375 194.650 65.680 194.780 ;
        RECT 63.720 194.225 64.230 194.315 ;
        RECT 63.720 194.055 64.590 194.225 ;
        RECT 63.720 193.985 63.890 194.055 ;
        RECT 64.010 193.805 64.210 193.835 ;
        RECT 62.530 193.445 62.995 193.775 ;
        RECT 63.380 193.505 64.210 193.805 ;
        RECT 63.380 193.275 63.550 193.505 ;
        RECT 62.190 193.105 62.975 193.275 ;
        RECT 63.145 193.105 63.550 193.275 ;
        RECT 63.730 192.825 64.100 193.325 ;
        RECT 64.420 193.275 64.590 194.055 ;
        RECT 64.760 193.695 64.930 194.395 ;
        RECT 65.100 193.865 65.340 194.460 ;
        RECT 64.760 193.475 65.285 193.695 ;
        RECT 65.510 193.545 65.680 194.650 ;
        RECT 65.455 193.415 65.680 193.545 ;
        RECT 65.850 193.455 66.130 194.405 ;
        RECT 65.455 193.275 65.625 193.415 ;
        RECT 64.420 193.105 65.095 193.275 ;
        RECT 65.290 193.105 65.625 193.275 ;
        RECT 65.795 192.825 66.045 193.285 ;
        RECT 66.300 193.085 66.485 195.205 ;
        RECT 66.655 194.875 66.985 195.375 ;
        RECT 67.155 194.705 67.325 195.205 ;
        RECT 66.660 194.535 67.325 194.705 ;
        RECT 66.660 193.545 66.890 194.535 ;
        RECT 67.060 193.715 67.410 194.365 ;
        RECT 67.585 194.285 69.255 195.375 ;
        RECT 69.485 194.315 69.815 195.160 ;
        RECT 69.985 194.365 70.155 195.375 ;
        RECT 70.325 194.645 70.665 195.205 ;
        RECT 70.895 194.875 71.210 195.375 ;
        RECT 71.390 194.905 72.275 195.075 ;
        RECT 67.585 193.595 68.335 194.115 ;
        RECT 68.505 193.765 69.255 194.285 ;
        RECT 69.425 194.235 69.815 194.315 ;
        RECT 70.325 194.270 71.220 194.645 ;
        RECT 69.425 194.185 69.640 194.235 ;
        RECT 69.425 193.605 69.595 194.185 ;
        RECT 70.325 194.065 70.515 194.270 ;
        RECT 71.390 194.065 71.560 194.905 ;
        RECT 72.500 194.875 72.750 195.205 ;
        RECT 69.765 193.735 70.515 194.065 ;
        RECT 70.685 193.735 71.560 194.065 ;
        RECT 66.660 193.375 67.325 193.545 ;
        RECT 66.655 192.825 66.985 193.205 ;
        RECT 67.155 193.085 67.325 193.375 ;
        RECT 67.585 192.825 69.255 193.595 ;
        RECT 69.425 193.565 69.650 193.605 ;
        RECT 70.315 193.565 70.515 193.735 ;
        RECT 69.425 193.480 69.805 193.565 ;
        RECT 69.475 193.045 69.805 193.480 ;
        RECT 69.975 192.825 70.145 193.435 ;
        RECT 70.315 193.040 70.645 193.565 ;
        RECT 70.905 192.825 71.115 193.355 ;
        RECT 71.390 193.275 71.560 193.735 ;
        RECT 71.730 193.775 72.050 194.735 ;
        RECT 72.220 193.985 72.410 194.705 ;
        RECT 72.580 193.805 72.750 194.875 ;
        RECT 72.920 194.575 73.090 195.375 ;
        RECT 73.260 194.930 74.365 195.100 ;
        RECT 73.260 194.315 73.430 194.930 ;
        RECT 74.575 194.780 74.825 195.205 ;
        RECT 74.995 194.915 75.260 195.375 ;
        RECT 73.600 194.395 74.130 194.760 ;
        RECT 74.575 194.650 74.880 194.780 ;
        RECT 72.920 194.225 73.430 194.315 ;
        RECT 72.920 194.055 73.790 194.225 ;
        RECT 72.920 193.985 73.090 194.055 ;
        RECT 73.210 193.805 73.410 193.835 ;
        RECT 71.730 193.445 72.195 193.775 ;
        RECT 72.580 193.505 73.410 193.805 ;
        RECT 72.580 193.275 72.750 193.505 ;
        RECT 71.390 193.105 72.175 193.275 ;
        RECT 72.345 193.105 72.750 193.275 ;
        RECT 72.930 192.825 73.300 193.325 ;
        RECT 73.620 193.275 73.790 194.055 ;
        RECT 73.960 193.695 74.130 194.395 ;
        RECT 74.300 193.865 74.540 194.460 ;
        RECT 73.960 193.475 74.485 193.695 ;
        RECT 74.710 193.545 74.880 194.650 ;
        RECT 74.655 193.415 74.880 193.545 ;
        RECT 75.050 193.455 75.330 194.405 ;
        RECT 74.655 193.275 74.825 193.415 ;
        RECT 73.620 193.105 74.295 193.275 ;
        RECT 74.490 193.105 74.825 193.275 ;
        RECT 74.995 192.825 75.245 193.285 ;
        RECT 75.500 193.085 75.685 195.205 ;
        RECT 75.855 194.875 76.185 195.375 ;
        RECT 76.355 194.705 76.525 195.205 ;
        RECT 75.860 194.535 76.525 194.705 ;
        RECT 75.860 193.545 76.090 194.535 ;
        RECT 76.260 193.715 76.610 194.365 ;
        RECT 76.785 194.285 77.995 195.375 ;
        RECT 76.785 193.575 77.305 194.115 ;
        RECT 77.475 193.745 77.995 194.285 ;
        RECT 78.350 194.405 78.740 194.580 ;
        RECT 79.225 194.575 79.555 195.375 ;
        RECT 79.725 194.585 80.260 195.205 ;
        RECT 78.350 194.235 79.775 194.405 ;
        RECT 75.860 193.375 76.525 193.545 ;
        RECT 75.855 192.825 76.185 193.205 ;
        RECT 76.355 193.085 76.525 193.375 ;
        RECT 76.785 192.825 77.995 193.575 ;
        RECT 78.225 193.505 78.580 194.065 ;
        RECT 78.750 193.335 78.920 194.235 ;
        RECT 79.090 193.505 79.355 194.065 ;
        RECT 79.605 193.735 79.775 194.235 ;
        RECT 79.945 193.565 80.260 194.585 ;
        RECT 78.330 192.825 78.570 193.335 ;
        RECT 78.750 193.005 79.030 193.335 ;
        RECT 79.260 192.825 79.475 193.335 ;
        RECT 79.645 192.995 80.260 193.565 ;
        RECT 80.465 194.655 80.925 195.205 ;
        RECT 81.115 194.655 81.445 195.375 ;
        RECT 80.465 193.285 80.715 194.655 ;
        RECT 81.645 194.485 81.945 195.035 ;
        RECT 82.115 194.705 82.395 195.375 ;
        RECT 81.005 194.315 81.945 194.485 ;
        RECT 81.005 194.065 81.175 194.315 ;
        RECT 82.315 194.065 82.580 194.425 ;
        RECT 82.765 194.210 83.055 195.375 ;
        RECT 83.225 194.525 83.565 195.165 ;
        RECT 83.735 194.915 83.980 195.375 ;
        RECT 84.155 194.745 84.405 195.205 ;
        RECT 84.595 194.995 85.265 195.375 ;
        RECT 85.465 194.745 85.715 195.205 ;
        RECT 84.155 194.575 85.715 194.745 ;
        RECT 80.885 193.735 81.175 194.065 ;
        RECT 81.345 193.815 81.685 194.065 ;
        RECT 81.905 193.815 82.580 194.065 ;
        RECT 81.005 193.645 81.175 193.735 ;
        RECT 81.005 193.455 82.395 193.645 ;
        RECT 80.465 192.995 81.025 193.285 ;
        RECT 81.195 192.825 81.445 193.285 ;
        RECT 82.065 193.095 82.395 193.455 ;
        RECT 82.765 192.825 83.055 193.550 ;
        RECT 83.225 193.410 83.395 194.525 ;
        RECT 86.475 194.405 86.645 195.205 ;
        RECT 83.705 194.235 86.645 194.405 ;
        RECT 86.905 194.235 87.185 195.375 ;
        RECT 83.705 194.065 83.875 194.235 ;
        RECT 87.355 194.225 87.685 195.205 ;
        RECT 87.855 194.235 88.115 195.375 ;
        RECT 88.285 194.285 90.875 195.375 ;
        RECT 83.565 193.735 83.875 194.065 ;
        RECT 84.045 193.735 84.380 194.065 ;
        RECT 83.705 193.565 83.875 193.735 ;
        RECT 83.225 192.995 83.535 193.410 ;
        RECT 83.705 193.395 84.400 193.565 ;
        RECT 84.650 193.490 84.845 194.065 ;
        RECT 85.105 193.735 85.450 194.065 ;
        RECT 85.760 193.735 86.235 194.065 ;
        RECT 86.490 193.735 86.675 194.065 ;
        RECT 86.915 193.795 87.250 194.065 ;
        RECT 85.105 193.505 85.295 193.735 ;
        RECT 87.420 193.625 87.590 194.225 ;
        RECT 87.760 193.815 88.095 194.065 ;
        RECT 83.730 192.825 84.060 193.205 ;
        RECT 84.230 193.165 84.400 193.395 ;
        RECT 85.465 193.395 86.645 193.565 ;
        RECT 85.465 193.165 85.635 193.395 ;
        RECT 84.230 192.995 85.635 193.165 ;
        RECT 85.905 192.825 86.235 193.225 ;
        RECT 86.475 192.995 86.645 193.395 ;
        RECT 86.905 192.825 87.215 193.625 ;
        RECT 87.420 192.995 88.115 193.625 ;
        RECT 88.285 193.595 89.495 194.115 ;
        RECT 89.665 193.765 90.875 194.285 ;
        RECT 91.045 194.285 92.255 195.375 ;
        RECT 91.045 193.745 91.565 194.285 ;
        RECT 88.285 192.825 90.875 193.595 ;
        RECT 91.735 193.575 92.255 194.115 ;
        RECT 91.045 192.825 92.255 193.575 ;
        RECT 18.280 192.655 92.340 192.825 ;
        RECT 18.365 191.905 19.575 192.655 ;
        RECT 19.745 192.110 25.090 192.655 ;
        RECT 18.365 191.365 18.885 191.905 ;
        RECT 19.055 191.195 19.575 191.735 ;
        RECT 21.330 191.280 21.670 192.110 ;
        RECT 26.275 192.105 26.445 192.395 ;
        RECT 26.615 192.275 26.945 192.655 ;
        RECT 26.275 191.935 26.940 192.105 ;
        RECT 18.365 190.105 19.575 191.195 ;
        RECT 23.150 190.540 23.500 191.790 ;
        RECT 26.190 191.115 26.540 191.765 ;
        RECT 26.710 190.945 26.940 191.935 ;
        RECT 26.275 190.775 26.940 190.945 ;
        RECT 19.745 190.105 25.090 190.540 ;
        RECT 26.275 190.275 26.445 190.775 ;
        RECT 26.615 190.105 26.945 190.605 ;
        RECT 27.115 190.275 27.300 192.395 ;
        RECT 27.555 192.195 27.805 192.655 ;
        RECT 27.975 192.205 28.310 192.375 ;
        RECT 28.505 192.205 29.180 192.375 ;
        RECT 27.975 192.065 28.145 192.205 ;
        RECT 27.470 191.075 27.750 192.025 ;
        RECT 27.920 191.935 28.145 192.065 ;
        RECT 27.920 190.830 28.090 191.935 ;
        RECT 28.315 191.785 28.840 192.005 ;
        RECT 28.260 191.020 28.500 191.615 ;
        RECT 28.670 191.085 28.840 191.785 ;
        RECT 29.010 191.425 29.180 192.205 ;
        RECT 29.500 192.155 29.870 192.655 ;
        RECT 30.050 192.205 30.455 192.375 ;
        RECT 30.625 192.205 31.410 192.375 ;
        RECT 30.050 191.975 30.220 192.205 ;
        RECT 29.390 191.675 30.220 191.975 ;
        RECT 30.605 191.705 31.070 192.035 ;
        RECT 29.390 191.645 29.590 191.675 ;
        RECT 29.710 191.425 29.880 191.495 ;
        RECT 29.010 191.255 29.880 191.425 ;
        RECT 29.370 191.165 29.880 191.255 ;
        RECT 27.920 190.700 28.225 190.830 ;
        RECT 28.670 190.720 29.200 191.085 ;
        RECT 27.540 190.105 27.805 190.565 ;
        RECT 27.975 190.275 28.225 190.700 ;
        RECT 29.370 190.550 29.540 191.165 ;
        RECT 28.435 190.380 29.540 190.550 ;
        RECT 29.710 190.105 29.880 190.905 ;
        RECT 30.050 190.605 30.220 191.675 ;
        RECT 30.390 190.775 30.580 191.495 ;
        RECT 30.750 190.745 31.070 191.705 ;
        RECT 31.240 191.745 31.410 192.205 ;
        RECT 31.685 192.125 31.895 192.655 ;
        RECT 32.155 191.915 32.485 192.440 ;
        RECT 32.655 192.045 32.825 192.655 ;
        RECT 32.995 192.000 33.325 192.435 ;
        RECT 32.995 191.915 33.375 192.000 ;
        RECT 32.285 191.745 32.485 191.915 ;
        RECT 33.150 191.875 33.375 191.915 ;
        RECT 31.240 191.415 32.115 191.745 ;
        RECT 32.285 191.415 33.035 191.745 ;
        RECT 30.050 190.275 30.300 190.605 ;
        RECT 31.240 190.575 31.410 191.415 ;
        RECT 32.285 191.210 32.475 191.415 ;
        RECT 33.205 191.295 33.375 191.875 ;
        RECT 34.015 191.845 34.285 192.655 ;
        RECT 34.455 191.845 34.785 192.485 ;
        RECT 34.955 191.845 35.195 192.655 ;
        RECT 35.385 191.905 36.595 192.655 ;
        RECT 34.005 191.415 34.355 191.665 ;
        RECT 33.160 191.245 33.375 191.295 ;
        RECT 34.525 191.245 34.695 191.845 ;
        RECT 34.865 191.415 35.215 191.665 ;
        RECT 35.385 191.365 35.905 191.905 ;
        RECT 36.805 191.835 37.035 192.655 ;
        RECT 37.205 191.855 37.535 192.485 ;
        RECT 31.580 190.835 32.475 191.210 ;
        RECT 32.985 191.165 33.375 191.245 ;
        RECT 30.525 190.405 31.410 190.575 ;
        RECT 31.590 190.105 31.905 190.605 ;
        RECT 32.135 190.275 32.475 190.835 ;
        RECT 32.645 190.105 32.815 191.115 ;
        RECT 32.985 190.320 33.315 191.165 ;
        RECT 34.015 190.105 34.345 191.245 ;
        RECT 34.525 191.075 35.205 191.245 ;
        RECT 36.075 191.195 36.595 191.735 ;
        RECT 36.785 191.415 37.115 191.665 ;
        RECT 37.285 191.255 37.535 191.855 ;
        RECT 37.705 191.835 37.915 192.655 ;
        RECT 38.145 191.885 39.815 192.655 ;
        RECT 40.100 192.025 40.385 192.485 ;
        RECT 40.555 192.195 40.825 192.655 ;
        RECT 38.145 191.365 38.895 191.885 ;
        RECT 40.100 191.855 41.055 192.025 ;
        RECT 34.875 190.290 35.205 191.075 ;
        RECT 35.385 190.105 36.595 191.195 ;
        RECT 36.805 190.105 37.035 191.245 ;
        RECT 37.205 190.275 37.535 191.255 ;
        RECT 37.705 190.105 37.915 191.245 ;
        RECT 39.065 191.195 39.815 191.715 ;
        RECT 38.145 190.105 39.815 191.195 ;
        RECT 39.985 191.125 40.675 191.685 ;
        RECT 40.845 190.955 41.055 191.855 ;
        RECT 40.100 190.735 41.055 190.955 ;
        RECT 41.225 191.685 41.625 192.485 ;
        RECT 41.815 192.025 42.095 192.485 ;
        RECT 42.615 192.195 42.940 192.655 ;
        RECT 41.815 191.855 42.940 192.025 ;
        RECT 43.110 191.915 43.495 192.485 ;
        RECT 44.125 191.930 44.415 192.655 ;
        RECT 45.135 192.005 45.305 192.485 ;
        RECT 45.475 192.175 45.805 192.655 ;
        RECT 46.030 192.235 47.565 192.485 ;
        RECT 46.030 192.005 46.200 192.235 ;
        RECT 42.490 191.745 42.940 191.855 ;
        RECT 41.225 191.125 42.320 191.685 ;
        RECT 42.490 191.415 43.045 191.745 ;
        RECT 40.100 190.275 40.385 190.735 ;
        RECT 40.555 190.105 40.825 190.565 ;
        RECT 41.225 190.275 41.625 191.125 ;
        RECT 42.490 190.955 42.940 191.415 ;
        RECT 43.215 191.245 43.495 191.915 ;
        RECT 45.135 191.835 46.200 192.005 ;
        RECT 46.380 191.665 46.660 192.065 ;
        RECT 45.050 191.455 45.400 191.665 ;
        RECT 45.570 191.465 46.015 191.665 ;
        RECT 46.185 191.465 46.660 191.665 ;
        RECT 46.930 191.665 47.215 192.065 ;
        RECT 47.395 192.005 47.565 192.235 ;
        RECT 47.735 192.175 48.065 192.655 ;
        RECT 48.280 192.155 48.535 192.485 ;
        RECT 48.350 192.075 48.535 192.155 ;
        RECT 47.395 191.835 48.195 192.005 ;
        RECT 46.930 191.465 47.260 191.665 ;
        RECT 47.430 191.635 47.795 191.665 ;
        RECT 47.430 191.465 47.805 191.635 ;
        RECT 48.025 191.285 48.195 191.835 ;
        RECT 41.815 190.735 42.940 190.955 ;
        RECT 41.815 190.275 42.095 190.735 ;
        RECT 42.615 190.105 42.940 190.565 ;
        RECT 43.110 190.275 43.495 191.245 ;
        RECT 44.125 190.105 44.415 191.270 ;
        RECT 45.135 191.115 48.195 191.285 ;
        RECT 45.135 190.275 45.305 191.115 ;
        RECT 48.365 190.945 48.535 192.075 ;
        RECT 48.725 191.885 51.315 192.655 ;
        RECT 51.485 192.045 51.825 192.460 ;
        RECT 51.995 192.215 52.165 192.655 ;
        RECT 52.335 192.265 53.585 192.445 ;
        RECT 52.335 192.045 52.665 192.265 ;
        RECT 53.855 192.195 54.025 192.655 ;
        RECT 48.725 191.365 49.935 191.885 ;
        RECT 51.485 191.875 52.665 192.045 ;
        RECT 52.835 192.025 53.200 192.095 ;
        RECT 52.835 191.845 54.085 192.025 ;
        RECT 50.105 191.195 51.315 191.715 ;
        RECT 51.485 191.465 51.950 191.665 ;
        RECT 52.125 191.415 52.455 191.665 ;
        RECT 52.625 191.635 53.090 191.665 ;
        RECT 52.625 191.465 53.095 191.635 ;
        RECT 52.625 191.415 53.090 191.465 ;
        RECT 53.285 191.415 53.640 191.665 ;
        RECT 52.125 191.295 52.305 191.415 ;
        RECT 45.475 190.445 45.805 190.945 ;
        RECT 45.975 190.705 47.610 190.945 ;
        RECT 45.975 190.615 46.205 190.705 ;
        RECT 46.315 190.445 46.645 190.485 ;
        RECT 45.475 190.275 46.645 190.445 ;
        RECT 46.835 190.105 47.190 190.525 ;
        RECT 47.360 190.275 47.610 190.705 ;
        RECT 47.780 190.105 48.110 190.865 ;
        RECT 48.280 190.275 48.535 190.945 ;
        RECT 48.725 190.105 51.315 191.195 ;
        RECT 51.485 190.105 51.805 191.285 ;
        RECT 51.975 191.125 52.305 191.295 ;
        RECT 53.810 191.245 54.085 191.845 ;
        RECT 51.975 190.335 52.175 191.125 ;
        RECT 52.475 191.035 54.085 191.245 ;
        RECT 52.475 190.935 52.885 191.035 ;
        RECT 52.500 190.275 52.885 190.935 ;
        RECT 53.280 190.105 54.065 190.865 ;
        RECT 54.255 190.275 54.535 192.375 ;
        RECT 54.705 192.110 60.050 192.655 ;
        RECT 56.290 191.280 56.630 192.110 ;
        RECT 60.225 191.885 62.815 192.655 ;
        RECT 63.000 192.085 63.255 192.435 ;
        RECT 63.425 192.255 63.755 192.655 ;
        RECT 63.925 192.085 64.095 192.435 ;
        RECT 64.265 192.255 64.645 192.655 ;
        RECT 63.000 191.915 64.665 192.085 ;
        RECT 64.835 191.980 65.110 192.325 ;
        RECT 58.110 190.540 58.460 191.790 ;
        RECT 60.225 191.365 61.435 191.885 ;
        RECT 64.495 191.745 64.665 191.915 ;
        RECT 61.605 191.195 62.815 191.715 ;
        RECT 62.985 191.415 63.330 191.745 ;
        RECT 63.500 191.415 64.325 191.745 ;
        RECT 64.495 191.415 64.770 191.745 ;
        RECT 54.705 190.105 60.050 190.540 ;
        RECT 60.225 190.105 62.815 191.195 ;
        RECT 63.005 190.955 63.330 191.245 ;
        RECT 63.500 191.125 63.695 191.415 ;
        RECT 64.495 191.245 64.665 191.415 ;
        RECT 64.940 191.245 65.110 191.980 ;
        RECT 65.285 191.885 68.795 192.655 ;
        RECT 69.885 191.930 70.175 192.655 ;
        RECT 71.265 191.980 71.540 192.325 ;
        RECT 71.730 192.255 72.105 192.655 ;
        RECT 72.275 192.085 72.445 192.435 ;
        RECT 72.615 192.255 72.945 192.655 ;
        RECT 73.115 192.085 73.375 192.485 ;
        RECT 65.285 191.365 66.935 191.885 ;
        RECT 64.005 191.075 64.665 191.245 ;
        RECT 64.005 190.955 64.175 191.075 ;
        RECT 63.005 190.785 64.175 190.955 ;
        RECT 62.985 190.325 64.175 190.615 ;
        RECT 64.345 190.105 64.625 190.905 ;
        RECT 64.835 190.275 65.110 191.245 ;
        RECT 67.105 191.195 68.795 191.715 ;
        RECT 65.285 190.105 68.795 191.195 ;
        RECT 69.885 190.105 70.175 191.270 ;
        RECT 71.265 191.245 71.435 191.980 ;
        RECT 71.710 191.915 73.375 192.085 ;
        RECT 71.710 191.745 71.880 191.915 ;
        RECT 73.555 191.835 73.885 192.255 ;
        RECT 74.055 191.835 74.315 192.655 ;
        RECT 74.485 192.110 79.830 192.655 ;
        RECT 73.555 191.745 73.805 191.835 ;
        RECT 71.605 191.415 71.880 191.745 ;
        RECT 72.050 191.415 72.875 191.745 ;
        RECT 73.090 191.415 73.805 191.745 ;
        RECT 73.975 191.415 74.310 191.665 ;
        RECT 71.710 191.245 71.880 191.415 ;
        RECT 71.265 190.275 71.540 191.245 ;
        RECT 71.710 191.075 72.370 191.245 ;
        RECT 72.630 191.125 72.875 191.415 ;
        RECT 72.200 190.955 72.370 191.075 ;
        RECT 73.045 190.955 73.375 191.245 ;
        RECT 71.750 190.105 72.030 190.905 ;
        RECT 72.200 190.785 73.375 190.955 ;
        RECT 73.635 190.855 73.805 191.415 ;
        RECT 76.070 191.280 76.410 192.110 ;
        RECT 80.005 191.885 81.675 192.655 ;
        RECT 82.395 192.105 82.565 192.395 ;
        RECT 82.735 192.275 83.065 192.655 ;
        RECT 82.395 191.935 83.060 192.105 ;
        RECT 72.200 190.285 73.815 190.615 ;
        RECT 74.055 190.105 74.315 191.245 ;
        RECT 77.890 190.540 78.240 191.790 ;
        RECT 80.005 191.365 80.755 191.885 ;
        RECT 80.925 191.195 81.675 191.715 ;
        RECT 74.485 190.105 79.830 190.540 ;
        RECT 80.005 190.105 81.675 191.195 ;
        RECT 82.310 191.115 82.660 191.765 ;
        RECT 82.830 190.945 83.060 191.935 ;
        RECT 82.395 190.775 83.060 190.945 ;
        RECT 82.395 190.275 82.565 190.775 ;
        RECT 82.735 190.105 83.065 190.605 ;
        RECT 83.235 190.275 83.460 192.395 ;
        RECT 83.675 192.195 83.925 192.655 ;
        RECT 84.110 192.205 84.440 192.375 ;
        RECT 84.620 192.205 85.370 192.375 ;
        RECT 83.660 191.075 83.940 191.675 ;
        RECT 84.110 190.675 84.280 192.205 ;
        RECT 84.450 191.705 85.030 192.035 ;
        RECT 84.450 190.835 84.690 191.705 ;
        RECT 85.200 191.425 85.370 192.205 ;
        RECT 85.620 192.155 85.990 192.655 ;
        RECT 86.170 192.205 86.630 192.375 ;
        RECT 86.860 192.205 87.530 192.375 ;
        RECT 86.170 191.975 86.340 192.205 ;
        RECT 85.540 191.675 86.340 191.975 ;
        RECT 86.510 191.705 87.060 192.035 ;
        RECT 85.540 191.645 85.710 191.675 ;
        RECT 85.830 191.425 86.000 191.495 ;
        RECT 85.200 191.255 86.000 191.425 ;
        RECT 85.490 191.165 86.000 191.255 ;
        RECT 84.880 190.730 85.320 191.085 ;
        RECT 83.660 190.105 83.925 190.565 ;
        RECT 84.110 190.300 84.345 190.675 ;
        RECT 85.490 190.550 85.660 191.165 ;
        RECT 84.590 190.380 85.660 190.550 ;
        RECT 85.830 190.105 86.000 190.905 ;
        RECT 86.170 190.605 86.340 191.675 ;
        RECT 86.510 190.775 86.700 191.495 ;
        RECT 86.870 191.165 87.060 191.705 ;
        RECT 87.360 191.665 87.530 192.205 ;
        RECT 87.845 192.125 88.015 192.655 ;
        RECT 88.310 192.005 88.670 192.445 ;
        RECT 88.845 192.175 89.015 192.655 ;
        RECT 89.205 192.010 89.540 192.435 ;
        RECT 89.715 192.180 89.885 192.655 ;
        RECT 90.060 192.010 90.395 192.435 ;
        RECT 90.565 192.180 90.735 192.655 ;
        RECT 88.310 191.835 88.810 192.005 ;
        RECT 89.205 191.840 90.875 192.010 ;
        RECT 91.045 191.905 92.255 192.655 ;
        RECT 88.640 191.665 88.810 191.835 ;
        RECT 87.360 191.495 88.450 191.665 ;
        RECT 88.640 191.495 90.460 191.665 ;
        RECT 86.870 190.835 87.190 191.165 ;
        RECT 86.170 190.275 86.420 190.605 ;
        RECT 87.360 190.575 87.530 191.495 ;
        RECT 88.640 191.240 88.810 191.495 ;
        RECT 90.630 191.275 90.875 191.840 ;
        RECT 87.700 191.070 88.810 191.240 ;
        RECT 89.205 191.105 90.875 191.275 ;
        RECT 91.045 191.195 91.565 191.735 ;
        RECT 91.735 191.365 92.255 191.905 ;
        RECT 87.700 190.910 88.560 191.070 ;
        RECT 86.645 190.405 87.530 190.575 ;
        RECT 87.710 190.105 87.925 190.605 ;
        RECT 88.390 190.285 88.560 190.910 ;
        RECT 88.845 190.105 89.025 190.885 ;
        RECT 89.205 190.345 89.540 191.105 ;
        RECT 89.720 190.105 89.890 190.935 ;
        RECT 90.060 190.345 90.390 191.105 ;
        RECT 90.560 190.105 90.730 190.935 ;
        RECT 91.045 190.105 92.255 191.195 ;
        RECT 18.280 189.935 92.340 190.105 ;
        RECT 18.365 188.845 19.575 189.935 ;
        RECT 19.745 189.500 25.090 189.935 ;
        RECT 18.365 188.135 18.885 188.675 ;
        RECT 19.055 188.305 19.575 188.845 ;
        RECT 18.365 187.385 19.575 188.135 ;
        RECT 21.330 187.930 21.670 188.760 ;
        RECT 23.150 188.250 23.500 189.500 ;
        RECT 25.265 188.845 27.855 189.935 ;
        RECT 25.265 188.155 26.475 188.675 ;
        RECT 26.645 188.325 27.855 188.845 ;
        RECT 28.035 188.965 28.365 189.750 ;
        RECT 28.035 188.795 28.715 188.965 ;
        RECT 28.895 188.795 29.225 189.935 ;
        RECT 29.405 188.845 31.075 189.935 ;
        RECT 28.025 188.375 28.375 188.625 ;
        RECT 28.545 188.195 28.715 188.795 ;
        RECT 28.885 188.375 29.235 188.625 ;
        RECT 19.745 187.385 25.090 187.930 ;
        RECT 25.265 187.385 27.855 188.155 ;
        RECT 28.045 187.385 28.285 188.195 ;
        RECT 28.455 187.555 28.785 188.195 ;
        RECT 28.955 187.385 29.225 188.195 ;
        RECT 29.405 188.155 30.155 188.675 ;
        RECT 30.325 188.325 31.075 188.845 ;
        RECT 31.245 188.770 31.535 189.935 ;
        RECT 31.705 188.845 32.915 189.935 ;
        RECT 29.405 187.385 31.075 188.155 ;
        RECT 31.705 188.135 32.225 188.675 ;
        RECT 32.395 188.305 32.915 188.845 ;
        RECT 33.085 188.795 33.470 189.755 ;
        RECT 33.685 189.135 33.975 189.935 ;
        RECT 34.145 189.595 35.510 189.765 ;
        RECT 34.145 188.965 34.315 189.595 ;
        RECT 33.640 188.795 34.315 188.965 ;
        RECT 33.085 188.745 33.315 188.795 ;
        RECT 31.245 187.385 31.535 188.110 ;
        RECT 31.705 187.385 32.915 188.135 ;
        RECT 33.085 188.125 33.260 188.745 ;
        RECT 33.640 188.625 33.810 188.795 ;
        RECT 34.485 188.625 34.810 189.425 ;
        RECT 35.180 189.385 35.510 189.595 ;
        RECT 35.180 189.135 36.135 189.385 ;
        RECT 33.445 188.375 33.810 188.625 ;
        RECT 34.005 188.375 34.255 188.625 ;
        RECT 33.445 188.295 33.635 188.375 ;
        RECT 34.005 188.295 34.175 188.375 ;
        RECT 34.465 188.295 34.810 188.625 ;
        RECT 34.980 188.295 35.255 188.960 ;
        RECT 35.440 188.295 35.795 188.960 ;
        RECT 35.965 188.125 36.135 189.135 ;
        RECT 36.305 188.795 36.595 189.935 ;
        RECT 37.690 189.555 38.025 189.935 ;
        RECT 36.320 188.295 36.595 188.625 ;
        RECT 33.085 187.555 33.595 188.125 ;
        RECT 34.140 187.955 35.540 188.125 ;
        RECT 33.765 187.385 33.935 187.945 ;
        RECT 34.140 187.555 34.470 187.955 ;
        RECT 34.645 187.385 34.975 187.785 ;
        RECT 35.210 187.765 35.540 187.955 ;
        RECT 35.710 187.935 36.135 188.125 ;
        RECT 37.685 188.065 37.925 189.375 ;
        RECT 38.195 188.965 38.445 189.765 ;
        RECT 38.665 189.215 38.995 189.935 ;
        RECT 39.180 188.965 39.430 189.765 ;
        RECT 39.895 189.135 40.225 189.935 ;
        RECT 40.395 189.505 40.735 189.765 ;
        RECT 38.095 188.795 40.285 188.965 ;
        RECT 36.305 187.765 36.595 188.035 ;
        RECT 38.095 187.885 38.265 188.795 ;
        RECT 39.970 188.625 40.285 188.795 ;
        RECT 35.210 187.555 36.595 187.765 ;
        RECT 37.770 187.555 38.265 187.885 ;
        RECT 38.485 187.660 38.835 188.625 ;
        RECT 39.015 187.655 39.315 188.625 ;
        RECT 39.495 187.655 39.775 188.625 ;
        RECT 39.970 188.375 40.300 188.625 ;
        RECT 39.955 187.385 40.225 188.185 ;
        RECT 40.475 188.105 40.735 189.505 ;
        RECT 41.455 189.315 41.625 189.745 ;
        RECT 41.795 189.485 42.125 189.935 ;
        RECT 41.455 189.085 42.130 189.315 ;
        RECT 40.395 187.595 40.735 188.105 ;
        RECT 41.425 188.065 41.725 188.915 ;
        RECT 41.895 188.435 42.130 189.085 ;
        RECT 42.300 188.775 42.585 189.720 ;
        RECT 42.765 189.465 43.450 189.935 ;
        RECT 42.760 188.945 43.455 189.255 ;
        RECT 43.630 188.880 43.935 189.665 ;
        RECT 42.300 188.625 43.160 188.775 ;
        RECT 42.300 188.605 43.585 188.625 ;
        RECT 41.895 188.105 42.430 188.435 ;
        RECT 42.600 188.245 43.585 188.605 ;
        RECT 41.895 187.955 42.115 188.105 ;
        RECT 41.370 187.385 41.705 187.890 ;
        RECT 41.875 187.580 42.115 187.955 ;
        RECT 42.600 187.910 42.770 188.245 ;
        RECT 43.760 188.075 43.935 188.880 ;
        RECT 44.165 188.795 44.395 189.935 ;
        RECT 44.565 188.785 44.895 189.765 ;
        RECT 45.065 188.795 45.275 189.935 ;
        RECT 45.505 188.845 47.175 189.935 ;
        RECT 44.145 188.375 44.475 188.625 ;
        RECT 42.395 187.715 42.770 187.910 ;
        RECT 42.395 187.570 42.565 187.715 ;
        RECT 43.130 187.385 43.525 187.880 ;
        RECT 43.695 187.555 43.935 188.075 ;
        RECT 44.165 187.385 44.395 188.205 ;
        RECT 44.645 188.185 44.895 188.785 ;
        RECT 44.565 187.555 44.895 188.185 ;
        RECT 45.065 187.385 45.275 188.205 ;
        RECT 45.505 188.155 46.255 188.675 ;
        RECT 46.425 188.325 47.175 188.845 ;
        RECT 47.345 188.860 47.615 189.765 ;
        RECT 47.785 189.175 48.115 189.935 ;
        RECT 48.295 189.005 48.465 189.765 ;
        RECT 45.505 187.385 47.175 188.155 ;
        RECT 47.345 188.060 47.515 188.860 ;
        RECT 47.800 188.835 48.465 189.005 ;
        RECT 48.725 188.845 52.235 189.935 ;
        RECT 47.800 188.690 47.970 188.835 ;
        RECT 47.685 188.360 47.970 188.690 ;
        RECT 47.800 188.105 47.970 188.360 ;
        RECT 48.205 188.285 48.535 188.655 ;
        RECT 48.725 188.155 50.375 188.675 ;
        RECT 50.545 188.325 52.235 188.845 ;
        RECT 53.415 188.925 53.585 189.765 ;
        RECT 53.755 189.595 54.925 189.765 ;
        RECT 53.755 189.095 54.085 189.595 ;
        RECT 54.595 189.555 54.925 189.595 ;
        RECT 55.115 189.515 55.470 189.935 ;
        RECT 54.255 189.335 54.485 189.425 ;
        RECT 55.640 189.335 55.890 189.765 ;
        RECT 54.255 189.095 55.890 189.335 ;
        RECT 56.060 189.175 56.390 189.935 ;
        RECT 56.560 189.095 56.815 189.765 ;
        RECT 53.415 188.755 56.475 188.925 ;
        RECT 53.330 188.375 53.680 188.585 ;
        RECT 53.850 188.375 54.295 188.575 ;
        RECT 54.465 188.375 54.940 188.575 ;
        RECT 47.345 187.555 47.605 188.060 ;
        RECT 47.800 187.935 48.465 188.105 ;
        RECT 47.785 187.385 48.115 187.765 ;
        RECT 48.295 187.555 48.465 187.935 ;
        RECT 48.725 187.385 52.235 188.155 ;
        RECT 53.415 188.035 54.480 188.205 ;
        RECT 53.415 187.555 53.585 188.035 ;
        RECT 53.755 187.385 54.085 187.865 ;
        RECT 54.310 187.805 54.480 188.035 ;
        RECT 54.660 187.975 54.940 188.375 ;
        RECT 55.210 188.375 55.540 188.575 ;
        RECT 55.710 188.405 56.085 188.575 ;
        RECT 55.710 188.375 56.075 188.405 ;
        RECT 55.210 187.975 55.495 188.375 ;
        RECT 56.305 188.205 56.475 188.755 ;
        RECT 55.675 188.035 56.475 188.205 ;
        RECT 55.675 187.805 55.845 188.035 ;
        RECT 56.645 187.965 56.815 189.095 ;
        RECT 57.005 188.770 57.295 189.935 ;
        RECT 57.530 188.965 57.800 189.760 ;
        RECT 57.980 189.135 58.195 189.935 ;
        RECT 58.375 188.965 58.660 189.760 ;
        RECT 57.530 188.795 58.660 188.965 ;
        RECT 57.510 188.325 58.010 188.590 ;
        RECT 58.230 188.295 58.615 188.625 ;
        RECT 58.840 188.295 59.120 189.765 ;
        RECT 59.300 188.350 59.630 189.765 ;
        RECT 59.800 188.590 60.005 189.765 ;
        RECT 60.175 188.945 60.385 189.760 ;
        RECT 60.625 189.115 60.955 189.935 ;
        RECT 60.175 188.765 60.825 188.945 ;
        RECT 61.130 188.920 61.385 189.760 ;
        RECT 59.800 188.350 60.230 188.590 ;
        RECT 58.230 188.145 58.535 188.295 ;
        RECT 56.630 187.885 56.815 187.965 ;
        RECT 54.310 187.555 55.845 187.805 ;
        RECT 56.015 187.385 56.345 187.865 ;
        RECT 56.560 187.555 56.815 187.885 ;
        RECT 57.005 187.385 57.295 188.110 ;
        RECT 57.565 187.385 57.805 188.060 ;
        RECT 57.980 187.585 58.535 188.145 ;
        RECT 60.605 188.125 60.825 188.765 ;
        RECT 58.715 187.955 60.825 188.125 ;
        RECT 58.715 187.560 58.920 187.955 ;
        RECT 59.605 187.950 60.825 187.955 ;
        RECT 59.090 187.385 59.435 187.785 ;
        RECT 59.605 187.560 59.935 187.950 ;
        RECT 60.210 187.385 60.885 187.770 ;
        RECT 61.055 187.555 61.385 188.920 ;
        RECT 61.605 188.825 61.865 189.765 ;
        RECT 62.035 189.535 62.365 189.935 ;
        RECT 63.510 189.670 63.765 189.765 ;
        RECT 62.625 189.500 63.765 189.670 ;
        RECT 63.935 189.555 64.265 189.725 ;
        RECT 62.625 189.275 62.795 189.500 ;
        RECT 62.035 189.105 62.795 189.275 ;
        RECT 63.510 189.365 63.765 189.500 ;
        RECT 61.605 188.110 61.780 188.825 ;
        RECT 62.035 188.625 62.205 189.105 ;
        RECT 63.060 189.015 63.230 189.205 ;
        RECT 63.510 189.195 63.920 189.365 ;
        RECT 61.950 188.295 62.205 188.625 ;
        RECT 62.430 188.295 62.760 188.915 ;
        RECT 63.060 188.845 63.580 189.015 ;
        RECT 62.930 188.295 63.220 188.675 ;
        RECT 63.410 188.125 63.580 188.845 ;
        RECT 61.605 187.555 61.865 188.110 ;
        RECT 62.700 187.955 63.580 188.125 ;
        RECT 63.750 188.170 63.920 189.195 ;
        RECT 64.095 189.305 64.265 189.555 ;
        RECT 64.435 189.475 64.685 189.935 ;
        RECT 64.855 189.305 65.035 189.765 ;
        RECT 64.095 189.135 65.035 189.305 ;
        RECT 64.120 188.655 64.600 188.955 ;
        RECT 63.750 188.000 64.100 188.170 ;
        RECT 64.340 188.065 64.600 188.655 ;
        RECT 64.800 188.065 65.060 188.955 ;
        RECT 65.305 188.880 65.610 189.665 ;
        RECT 65.790 189.465 66.475 189.935 ;
        RECT 65.785 188.945 66.480 189.255 ;
        RECT 65.305 188.075 65.480 188.880 ;
        RECT 66.655 188.775 66.940 189.720 ;
        RECT 67.115 189.485 67.445 189.935 ;
        RECT 67.615 189.315 67.785 189.745 ;
        RECT 66.080 188.625 66.940 188.775 ;
        RECT 65.655 188.605 66.940 188.625 ;
        RECT 67.110 189.085 67.785 189.315 ;
        RECT 69.055 189.315 69.225 189.745 ;
        RECT 69.395 189.485 69.725 189.935 ;
        RECT 69.055 189.085 69.730 189.315 ;
        RECT 65.655 188.245 66.640 188.605 ;
        RECT 67.110 188.435 67.345 189.085 ;
        RECT 62.035 187.385 62.465 187.830 ;
        RECT 62.700 187.555 62.870 187.955 ;
        RECT 63.040 187.385 63.760 187.785 ;
        RECT 63.930 187.555 64.100 188.000 ;
        RECT 64.675 187.385 65.075 187.895 ;
        RECT 65.305 187.555 65.545 188.075 ;
        RECT 66.470 187.910 66.640 188.245 ;
        RECT 66.810 188.105 67.345 188.435 ;
        RECT 67.125 187.955 67.345 188.105 ;
        RECT 67.515 188.065 67.815 188.915 ;
        RECT 69.025 188.065 69.325 188.915 ;
        RECT 69.495 188.435 69.730 189.085 ;
        RECT 69.900 188.775 70.185 189.720 ;
        RECT 70.365 189.465 71.050 189.935 ;
        RECT 70.360 188.945 71.055 189.255 ;
        RECT 71.230 188.880 71.535 189.665 ;
        RECT 69.900 188.625 70.760 188.775 ;
        RECT 69.900 188.605 71.185 188.625 ;
        RECT 69.495 188.105 70.030 188.435 ;
        RECT 70.200 188.245 71.185 188.605 ;
        RECT 69.495 187.955 69.715 188.105 ;
        RECT 65.715 187.385 66.110 187.880 ;
        RECT 66.470 187.715 66.845 187.910 ;
        RECT 66.675 187.570 66.845 187.715 ;
        RECT 67.125 187.580 67.365 187.955 ;
        RECT 67.535 187.385 67.870 187.890 ;
        RECT 68.970 187.385 69.305 187.890 ;
        RECT 69.475 187.580 69.715 187.955 ;
        RECT 70.200 187.910 70.370 188.245 ;
        RECT 71.360 188.075 71.535 188.880 ;
        RECT 71.785 188.795 71.995 189.935 ;
        RECT 72.165 188.785 72.495 189.765 ;
        RECT 72.665 188.795 72.895 189.935 ;
        RECT 73.565 188.795 73.835 189.765 ;
        RECT 74.045 189.135 74.325 189.935 ;
        RECT 74.505 189.385 75.700 189.715 ;
        RECT 74.830 188.965 75.250 189.215 ;
        RECT 74.005 188.795 75.250 188.965 ;
        RECT 69.995 187.715 70.370 187.910 ;
        RECT 69.995 187.570 70.165 187.715 ;
        RECT 70.730 187.385 71.125 187.880 ;
        RECT 71.295 187.555 71.535 188.075 ;
        RECT 71.785 187.385 71.995 188.205 ;
        RECT 72.165 188.185 72.415 188.785 ;
        RECT 72.585 188.375 72.915 188.625 ;
        RECT 72.165 187.555 72.495 188.185 ;
        RECT 72.665 187.385 72.895 188.205 ;
        RECT 73.565 188.060 73.735 188.795 ;
        RECT 74.005 188.625 74.175 188.795 ;
        RECT 75.475 188.625 75.645 189.185 ;
        RECT 75.895 188.795 76.150 189.935 ;
        RECT 76.325 189.500 81.670 189.935 ;
        RECT 73.945 188.295 74.175 188.625 ;
        RECT 74.905 188.295 75.645 188.625 ;
        RECT 75.815 188.375 76.150 188.625 ;
        RECT 74.005 188.125 74.175 188.295 ;
        RECT 75.395 188.205 75.645 188.295 ;
        RECT 73.565 187.715 73.835 188.060 ;
        RECT 74.005 187.955 74.745 188.125 ;
        RECT 75.395 188.035 76.130 188.205 ;
        RECT 74.025 187.385 74.405 187.785 ;
        RECT 74.575 187.605 74.745 187.955 ;
        RECT 74.915 187.385 75.650 187.865 ;
        RECT 75.820 187.565 76.130 188.035 ;
        RECT 77.910 187.930 78.250 188.760 ;
        RECT 79.730 188.250 80.080 189.500 ;
        RECT 82.765 188.770 83.055 189.935 ;
        RECT 83.225 189.500 88.570 189.935 ;
        RECT 76.325 187.385 81.670 187.930 ;
        RECT 82.765 187.385 83.055 188.110 ;
        RECT 84.810 187.930 85.150 188.760 ;
        RECT 86.630 188.250 86.980 189.500 ;
        RECT 88.745 188.845 90.415 189.935 ;
        RECT 88.745 188.155 89.495 188.675 ;
        RECT 89.665 188.325 90.415 188.845 ;
        RECT 91.045 188.845 92.255 189.935 ;
        RECT 91.045 188.305 91.565 188.845 ;
        RECT 83.225 187.385 88.570 187.930 ;
        RECT 88.745 187.385 90.415 188.155 ;
        RECT 91.735 188.135 92.255 188.675 ;
        RECT 91.045 187.385 92.255 188.135 ;
        RECT 18.280 187.215 92.340 187.385 ;
        RECT 18.365 186.465 19.575 187.215 ;
        RECT 20.715 186.560 21.045 186.995 ;
        RECT 21.215 186.605 21.385 187.215 ;
        RECT 20.665 186.475 21.045 186.560 ;
        RECT 21.555 186.475 21.885 187.000 ;
        RECT 22.145 186.685 22.355 187.215 ;
        RECT 22.630 186.765 23.415 186.935 ;
        RECT 23.585 186.765 23.990 186.935 ;
        RECT 18.365 185.925 18.885 186.465 ;
        RECT 20.665 186.435 20.890 186.475 ;
        RECT 19.055 185.755 19.575 186.295 ;
        RECT 18.365 184.665 19.575 185.755 ;
        RECT 20.665 185.855 20.835 186.435 ;
        RECT 21.555 186.305 21.755 186.475 ;
        RECT 22.630 186.305 22.800 186.765 ;
        RECT 21.005 185.975 21.755 186.305 ;
        RECT 21.925 185.975 22.800 186.305 ;
        RECT 20.665 185.805 20.880 185.855 ;
        RECT 20.665 185.725 21.055 185.805 ;
        RECT 20.725 184.880 21.055 185.725 ;
        RECT 21.565 185.770 21.755 185.975 ;
        RECT 21.225 184.665 21.395 185.675 ;
        RECT 21.565 185.395 22.460 185.770 ;
        RECT 21.565 184.835 21.905 185.395 ;
        RECT 22.135 184.665 22.450 185.165 ;
        RECT 22.630 185.135 22.800 185.975 ;
        RECT 22.970 186.265 23.435 186.595 ;
        RECT 23.820 186.535 23.990 186.765 ;
        RECT 24.170 186.715 24.540 187.215 ;
        RECT 24.860 186.765 25.535 186.935 ;
        RECT 25.730 186.765 26.065 186.935 ;
        RECT 22.970 185.305 23.290 186.265 ;
        RECT 23.820 186.235 24.650 186.535 ;
        RECT 23.460 185.335 23.650 186.055 ;
        RECT 23.820 185.165 23.990 186.235 ;
        RECT 24.450 186.205 24.650 186.235 ;
        RECT 24.160 185.985 24.330 186.055 ;
        RECT 24.860 185.985 25.030 186.765 ;
        RECT 25.895 186.625 26.065 186.765 ;
        RECT 26.235 186.755 26.485 187.215 ;
        RECT 24.160 185.815 25.030 185.985 ;
        RECT 25.200 186.345 25.725 186.565 ;
        RECT 25.895 186.495 26.120 186.625 ;
        RECT 24.160 185.725 24.670 185.815 ;
        RECT 22.630 184.965 23.515 185.135 ;
        RECT 23.740 184.835 23.990 185.165 ;
        RECT 24.160 184.665 24.330 185.465 ;
        RECT 24.500 185.110 24.670 185.725 ;
        RECT 25.200 185.645 25.370 186.345 ;
        RECT 24.840 185.280 25.370 185.645 ;
        RECT 25.540 185.580 25.780 186.175 ;
        RECT 25.950 185.390 26.120 186.495 ;
        RECT 26.290 185.635 26.570 186.585 ;
        RECT 25.815 185.260 26.120 185.390 ;
        RECT 24.500 184.940 25.605 185.110 ;
        RECT 25.815 184.835 26.065 185.260 ;
        RECT 26.235 184.665 26.500 185.125 ;
        RECT 26.740 184.835 26.925 186.955 ;
        RECT 27.095 186.835 27.425 187.215 ;
        RECT 27.595 186.665 27.765 186.955 ;
        RECT 27.100 186.495 27.765 186.665 ;
        RECT 27.100 185.505 27.330 186.495 ;
        RECT 28.025 186.475 28.410 187.045 ;
        RECT 28.580 186.755 28.905 187.215 ;
        RECT 29.425 186.585 29.705 187.045 ;
        RECT 27.500 185.675 27.850 186.325 ;
        RECT 28.025 185.805 28.305 186.475 ;
        RECT 28.580 186.415 29.705 186.585 ;
        RECT 28.580 186.305 29.030 186.415 ;
        RECT 28.475 185.975 29.030 186.305 ;
        RECT 29.895 186.245 30.295 187.045 ;
        RECT 30.695 186.755 30.965 187.215 ;
        RECT 31.135 186.585 31.420 187.045 ;
        RECT 27.100 185.335 27.765 185.505 ;
        RECT 27.095 184.665 27.425 185.165 ;
        RECT 27.595 184.835 27.765 185.335 ;
        RECT 28.025 184.835 28.410 185.805 ;
        RECT 28.580 185.515 29.030 185.975 ;
        RECT 29.200 185.685 30.295 186.245 ;
        RECT 28.580 185.295 29.705 185.515 ;
        RECT 28.580 184.665 28.905 185.125 ;
        RECT 29.425 184.835 29.705 185.295 ;
        RECT 29.895 184.835 30.295 185.685 ;
        RECT 30.465 186.415 31.420 186.585 ;
        RECT 30.465 185.515 30.675 186.415 ;
        RECT 30.845 185.685 31.535 186.245 ;
        RECT 31.710 185.615 32.045 187.035 ;
        RECT 32.225 186.845 32.970 187.215 ;
        RECT 33.535 186.675 33.790 187.035 ;
        RECT 33.970 186.845 34.300 187.215 ;
        RECT 34.480 186.675 34.705 187.035 ;
        RECT 32.220 186.485 34.705 186.675 ;
        RECT 32.220 185.795 32.445 186.485 ;
        RECT 34.945 186.405 35.185 187.215 ;
        RECT 35.355 186.405 35.685 187.045 ;
        RECT 35.855 186.405 36.125 187.215 ;
        RECT 36.305 186.475 36.815 187.045 ;
        RECT 36.985 186.655 37.155 187.215 ;
        RECT 37.360 186.645 37.690 187.045 ;
        RECT 37.865 186.815 38.195 187.215 ;
        RECT 38.430 186.835 39.815 187.045 ;
        RECT 38.430 186.645 38.760 186.835 ;
        RECT 37.360 186.475 38.760 186.645 ;
        RECT 38.930 186.475 39.355 186.665 ;
        RECT 39.525 186.565 39.815 186.835 ;
        RECT 40.010 186.825 40.340 187.215 ;
        RECT 40.510 186.655 40.735 187.035 ;
        RECT 32.645 185.975 32.925 186.305 ;
        RECT 33.105 185.975 33.680 186.305 ;
        RECT 33.860 185.975 34.295 186.305 ;
        RECT 34.475 185.975 34.745 186.305 ;
        RECT 34.925 185.975 35.275 186.225 ;
        RECT 35.445 185.805 35.615 186.405 ;
        RECT 35.785 185.975 36.135 186.225 ;
        RECT 36.305 185.805 36.480 186.475 ;
        RECT 36.665 186.225 36.855 186.305 ;
        RECT 37.225 186.225 37.395 186.305 ;
        RECT 36.665 185.975 37.030 186.225 ;
        RECT 37.225 185.975 37.475 186.225 ;
        RECT 37.685 185.975 38.030 186.305 ;
        RECT 36.860 185.805 37.030 185.975 ;
        RECT 32.220 185.615 34.715 185.795 ;
        RECT 30.465 185.295 31.420 185.515 ;
        RECT 30.695 184.665 30.965 185.125 ;
        RECT 31.135 184.835 31.420 185.295 ;
        RECT 31.710 184.845 31.975 185.615 ;
        RECT 32.145 184.665 32.475 185.385 ;
        RECT 32.665 185.205 33.855 185.435 ;
        RECT 32.665 184.845 32.925 185.205 ;
        RECT 33.095 184.665 33.425 185.035 ;
        RECT 33.595 184.845 33.855 185.205 ;
        RECT 34.425 184.845 34.715 185.615 ;
        RECT 34.935 185.635 35.615 185.805 ;
        RECT 34.935 184.850 35.265 185.635 ;
        RECT 35.795 184.665 36.125 185.805 ;
        RECT 36.305 184.845 36.690 185.805 ;
        RECT 36.860 185.635 37.535 185.805 ;
        RECT 36.905 184.665 37.195 185.465 ;
        RECT 37.365 185.005 37.535 185.635 ;
        RECT 37.705 185.175 38.030 185.975 ;
        RECT 38.200 185.640 38.475 186.305 ;
        RECT 38.660 185.640 39.015 186.305 ;
        RECT 39.185 185.465 39.355 186.475 ;
        RECT 39.540 185.975 39.815 186.305 ;
        RECT 39.995 185.975 40.235 186.625 ;
        RECT 40.405 186.475 40.735 186.655 ;
        RECT 40.405 185.805 40.580 186.475 ;
        RECT 40.935 186.305 41.165 186.925 ;
        RECT 41.345 186.485 41.645 187.215 ;
        RECT 41.885 186.395 42.095 187.215 ;
        RECT 42.265 186.415 42.595 187.045 ;
        RECT 40.750 185.975 41.165 186.305 ;
        RECT 41.345 185.975 41.640 186.305 ;
        RECT 42.265 185.815 42.515 186.415 ;
        RECT 42.765 186.395 42.995 187.215 ;
        RECT 44.125 186.490 44.415 187.215 ;
        RECT 45.595 186.665 45.765 186.955 ;
        RECT 45.935 186.835 46.265 187.215 ;
        RECT 45.595 186.495 46.260 186.665 ;
        RECT 42.685 185.975 43.015 186.225 ;
        RECT 38.400 185.215 39.355 185.465 ;
        RECT 38.400 185.005 38.730 185.215 ;
        RECT 37.365 184.835 38.730 185.005 ;
        RECT 39.525 184.665 39.815 185.805 ;
        RECT 39.995 185.615 40.580 185.805 ;
        RECT 39.995 184.845 40.270 185.615 ;
        RECT 40.750 185.445 41.645 185.775 ;
        RECT 40.440 185.275 41.645 185.445 ;
        RECT 40.440 184.845 40.770 185.275 ;
        RECT 40.940 184.665 41.135 185.105 ;
        RECT 41.315 184.845 41.645 185.275 ;
        RECT 41.885 184.665 42.095 185.805 ;
        RECT 42.265 184.835 42.595 185.815 ;
        RECT 42.765 184.665 42.995 185.805 ;
        RECT 44.125 184.665 44.415 185.830 ;
        RECT 45.510 185.675 45.860 186.325 ;
        RECT 46.030 185.505 46.260 186.495 ;
        RECT 45.595 185.335 46.260 185.505 ;
        RECT 45.595 184.835 45.765 185.335 ;
        RECT 45.935 184.665 46.265 185.165 ;
        RECT 46.435 184.835 46.620 186.955 ;
        RECT 46.875 186.755 47.125 187.215 ;
        RECT 47.295 186.765 47.630 186.935 ;
        RECT 47.825 186.765 48.500 186.935 ;
        RECT 47.295 186.625 47.465 186.765 ;
        RECT 46.790 185.635 47.070 186.585 ;
        RECT 47.240 186.495 47.465 186.625 ;
        RECT 47.240 185.390 47.410 186.495 ;
        RECT 47.635 186.345 48.160 186.565 ;
        RECT 47.580 185.580 47.820 186.175 ;
        RECT 47.990 185.645 48.160 186.345 ;
        RECT 48.330 185.985 48.500 186.765 ;
        RECT 48.820 186.715 49.190 187.215 ;
        RECT 49.370 186.765 49.775 186.935 ;
        RECT 49.945 186.765 50.730 186.935 ;
        RECT 49.370 186.535 49.540 186.765 ;
        RECT 48.710 186.235 49.540 186.535 ;
        RECT 49.925 186.265 50.390 186.595 ;
        RECT 48.710 186.205 48.910 186.235 ;
        RECT 49.030 185.985 49.200 186.055 ;
        RECT 48.330 185.815 49.200 185.985 ;
        RECT 48.690 185.725 49.200 185.815 ;
        RECT 47.240 185.260 47.545 185.390 ;
        RECT 47.990 185.280 48.520 185.645 ;
        RECT 46.860 184.665 47.125 185.125 ;
        RECT 47.295 184.835 47.545 185.260 ;
        RECT 48.690 185.110 48.860 185.725 ;
        RECT 47.755 184.940 48.860 185.110 ;
        RECT 49.030 184.665 49.200 185.465 ;
        RECT 49.370 185.165 49.540 186.235 ;
        RECT 49.710 185.335 49.900 186.055 ;
        RECT 50.070 185.305 50.390 186.265 ;
        RECT 50.560 186.305 50.730 186.765 ;
        RECT 51.005 186.685 51.215 187.215 ;
        RECT 51.475 186.475 51.805 187.000 ;
        RECT 51.975 186.605 52.145 187.215 ;
        RECT 52.315 186.560 52.645 186.995 ;
        RECT 52.865 186.670 58.210 187.215 ;
        RECT 52.315 186.475 52.695 186.560 ;
        RECT 51.605 186.305 51.805 186.475 ;
        RECT 52.470 186.435 52.695 186.475 ;
        RECT 50.560 185.975 51.435 186.305 ;
        RECT 51.605 185.975 52.355 186.305 ;
        RECT 49.370 184.835 49.620 185.165 ;
        RECT 50.560 185.135 50.730 185.975 ;
        RECT 51.605 185.770 51.795 185.975 ;
        RECT 52.525 185.855 52.695 186.435 ;
        RECT 52.480 185.805 52.695 185.855 ;
        RECT 54.450 185.840 54.790 186.670 ;
        RECT 58.385 186.445 60.055 187.215 ;
        RECT 60.225 186.605 60.565 187.020 ;
        RECT 60.735 186.775 60.905 187.215 ;
        RECT 61.075 186.825 62.325 187.005 ;
        RECT 61.075 186.605 61.405 186.825 ;
        RECT 62.595 186.755 62.765 187.215 ;
        RECT 50.900 185.395 51.795 185.770 ;
        RECT 52.305 185.725 52.695 185.805 ;
        RECT 49.845 184.965 50.730 185.135 ;
        RECT 50.910 184.665 51.225 185.165 ;
        RECT 51.455 184.835 51.795 185.395 ;
        RECT 51.965 184.665 52.135 185.675 ;
        RECT 52.305 184.880 52.635 185.725 ;
        RECT 56.270 185.100 56.620 186.350 ;
        RECT 58.385 185.925 59.135 186.445 ;
        RECT 60.225 186.435 61.405 186.605 ;
        RECT 61.575 186.585 61.940 186.655 ;
        RECT 61.575 186.405 62.825 186.585 ;
        RECT 59.305 185.755 60.055 186.275 ;
        RECT 60.225 186.025 60.690 186.225 ;
        RECT 60.865 185.975 61.195 186.225 ;
        RECT 61.365 186.195 61.830 186.225 ;
        RECT 61.365 186.025 61.835 186.195 ;
        RECT 61.365 185.975 61.830 186.025 ;
        RECT 62.025 185.975 62.380 186.225 ;
        RECT 60.865 185.855 61.045 185.975 ;
        RECT 52.865 184.665 58.210 185.100 ;
        RECT 58.385 184.665 60.055 185.755 ;
        RECT 60.225 184.665 60.545 185.845 ;
        RECT 60.715 185.685 61.045 185.855 ;
        RECT 62.550 185.805 62.825 186.405 ;
        RECT 60.715 184.895 60.915 185.685 ;
        RECT 61.215 185.595 62.825 185.805 ;
        RECT 61.215 185.495 61.625 185.595 ;
        RECT 61.240 184.835 61.625 185.495 ;
        RECT 62.020 184.665 62.805 185.425 ;
        RECT 62.995 184.835 63.275 186.935 ;
        RECT 63.445 186.475 63.885 187.035 ;
        RECT 64.055 186.475 64.505 187.215 ;
        RECT 64.675 186.645 64.845 187.045 ;
        RECT 65.015 186.815 65.435 187.215 ;
        RECT 65.605 186.645 65.835 187.045 ;
        RECT 64.675 186.475 65.835 186.645 ;
        RECT 66.005 186.475 66.495 187.045 ;
        RECT 63.445 185.465 63.755 186.475 ;
        RECT 63.925 185.855 64.095 186.305 ;
        RECT 64.265 186.025 64.655 186.305 ;
        RECT 64.840 185.975 65.085 186.305 ;
        RECT 63.925 185.685 64.715 185.855 ;
        RECT 63.445 184.835 63.885 185.465 ;
        RECT 64.060 184.665 64.375 185.515 ;
        RECT 64.545 185.005 64.715 185.685 ;
        RECT 64.885 185.175 65.085 185.975 ;
        RECT 65.285 185.175 65.535 186.305 ;
        RECT 65.750 185.975 66.155 186.305 ;
        RECT 66.325 185.805 66.495 186.475 ;
        RECT 67.150 186.565 67.460 187.035 ;
        RECT 67.630 186.735 68.365 187.215 ;
        RECT 68.535 186.645 68.705 186.995 ;
        RECT 68.875 186.815 69.255 187.215 ;
        RECT 67.150 186.395 67.885 186.565 ;
        RECT 68.535 186.475 69.275 186.645 ;
        RECT 69.445 186.540 69.715 186.885 ;
        RECT 67.635 186.305 67.885 186.395 ;
        RECT 69.105 186.305 69.275 186.475 ;
        RECT 67.130 185.975 67.465 186.225 ;
        RECT 67.635 185.975 68.375 186.305 ;
        RECT 69.105 185.975 69.335 186.305 ;
        RECT 65.725 185.635 66.495 185.805 ;
        RECT 65.725 185.005 65.975 185.635 ;
        RECT 64.545 184.835 65.975 185.005 ;
        RECT 66.155 184.665 66.485 185.465 ;
        RECT 67.130 184.665 67.385 185.805 ;
        RECT 67.635 185.415 67.805 185.975 ;
        RECT 69.105 185.805 69.275 185.975 ;
        RECT 69.545 185.855 69.715 186.540 ;
        RECT 69.885 186.490 70.175 187.215 ;
        RECT 70.345 186.540 70.620 186.885 ;
        RECT 70.810 186.815 71.185 187.215 ;
        RECT 71.355 186.645 71.525 186.995 ;
        RECT 71.695 186.815 72.025 187.215 ;
        RECT 72.195 186.645 72.455 187.045 ;
        RECT 69.485 185.805 69.715 185.855 ;
        RECT 68.030 185.635 69.275 185.805 ;
        RECT 68.030 185.385 68.450 185.635 ;
        RECT 67.580 184.885 68.775 185.215 ;
        RECT 68.955 184.665 69.235 185.465 ;
        RECT 69.445 184.835 69.715 185.805 ;
        RECT 69.885 184.665 70.175 185.830 ;
        RECT 70.345 185.805 70.515 186.540 ;
        RECT 70.790 186.475 72.455 186.645 ;
        RECT 70.790 186.305 70.960 186.475 ;
        RECT 72.635 186.395 72.965 186.815 ;
        RECT 73.135 186.395 73.395 187.215 ;
        RECT 72.635 186.305 72.885 186.395 ;
        RECT 73.565 186.380 73.855 187.215 ;
        RECT 74.025 186.815 74.980 186.985 ;
        RECT 75.395 186.825 75.725 187.215 ;
        RECT 70.685 185.975 70.960 186.305 ;
        RECT 71.130 185.975 71.955 186.305 ;
        RECT 72.170 185.975 72.885 186.305 ;
        RECT 73.055 185.975 73.390 186.225 ;
        RECT 70.790 185.805 70.960 185.975 ;
        RECT 70.345 184.835 70.620 185.805 ;
        RECT 70.790 185.635 71.450 185.805 ;
        RECT 71.710 185.685 71.955 185.975 ;
        RECT 71.280 185.515 71.450 185.635 ;
        RECT 72.125 185.515 72.455 185.805 ;
        RECT 70.830 184.665 71.110 185.465 ;
        RECT 71.280 185.345 72.455 185.515 ;
        RECT 72.715 185.415 72.885 185.975 ;
        RECT 74.025 185.935 74.195 186.815 ;
        RECT 75.895 186.645 76.065 186.965 ;
        RECT 76.235 186.825 76.565 187.215 ;
        RECT 74.365 186.475 76.615 186.645 ;
        RECT 74.365 185.975 74.595 186.475 ;
        RECT 74.765 186.055 75.140 186.225 ;
        RECT 71.280 184.845 72.895 185.175 ;
        RECT 73.135 184.665 73.395 185.805 ;
        RECT 73.565 185.765 74.195 185.935 ;
        RECT 74.970 185.855 75.140 186.055 ;
        RECT 75.310 186.025 75.860 186.225 ;
        RECT 76.030 185.855 76.275 186.305 ;
        RECT 73.565 184.835 73.885 185.765 ;
        RECT 74.970 185.685 76.275 185.855 ;
        RECT 76.445 185.515 76.615 186.475 ;
        RECT 77.255 186.405 77.525 187.215 ;
        RECT 77.695 186.405 78.025 187.045 ;
        RECT 78.195 186.405 78.435 187.215 ;
        RECT 78.715 186.565 78.885 187.045 ;
        RECT 79.055 186.735 79.385 187.215 ;
        RECT 79.610 186.795 81.145 187.045 ;
        RECT 79.610 186.565 79.780 186.795 ;
        RECT 77.245 185.975 77.595 186.225 ;
        RECT 77.765 185.805 77.935 186.405 ;
        RECT 78.715 186.395 79.780 186.565 ;
        RECT 79.960 186.225 80.240 186.625 ;
        RECT 78.105 185.975 78.455 186.225 ;
        RECT 78.630 186.015 78.980 186.225 ;
        RECT 79.150 186.025 79.595 186.225 ;
        RECT 79.765 186.025 80.240 186.225 ;
        RECT 80.510 186.225 80.795 186.625 ;
        RECT 80.975 186.565 81.145 186.795 ;
        RECT 81.315 186.735 81.645 187.215 ;
        RECT 81.860 186.715 82.115 187.045 ;
        RECT 81.930 186.635 82.115 186.715 ;
        RECT 80.975 186.395 81.775 186.565 ;
        RECT 80.510 186.025 80.840 186.225 ;
        RECT 81.010 186.025 81.375 186.225 ;
        RECT 81.605 185.845 81.775 186.395 ;
        RECT 74.065 185.345 75.305 185.515 ;
        RECT 74.065 184.835 74.465 185.345 ;
        RECT 74.635 184.665 74.805 185.175 ;
        RECT 74.975 184.835 75.305 185.345 ;
        RECT 75.475 184.665 75.645 185.515 ;
        RECT 76.235 184.835 76.615 185.515 ;
        RECT 77.255 184.665 77.585 185.805 ;
        RECT 77.765 185.635 78.445 185.805 ;
        RECT 78.115 184.850 78.445 185.635 ;
        RECT 78.715 185.675 81.775 185.845 ;
        RECT 78.715 184.835 78.885 185.675 ;
        RECT 81.945 185.505 82.115 186.635 ;
        RECT 82.395 186.665 82.565 186.955 ;
        RECT 82.735 186.835 83.065 187.215 ;
        RECT 82.395 186.495 83.060 186.665 ;
        RECT 82.310 185.675 82.660 186.325 ;
        RECT 82.830 185.505 83.060 186.495 ;
        RECT 79.055 185.005 79.385 185.505 ;
        RECT 79.555 185.265 81.190 185.505 ;
        RECT 79.555 185.175 79.785 185.265 ;
        RECT 79.895 185.005 80.225 185.045 ;
        RECT 79.055 184.835 80.225 185.005 ;
        RECT 80.415 184.665 80.770 185.085 ;
        RECT 80.940 184.835 81.190 185.265 ;
        RECT 81.360 184.665 81.690 185.425 ;
        RECT 81.860 184.835 82.115 185.505 ;
        RECT 82.395 185.335 83.060 185.505 ;
        RECT 82.395 184.835 82.565 185.335 ;
        RECT 82.735 184.665 83.065 185.165 ;
        RECT 83.235 184.835 83.460 186.955 ;
        RECT 83.675 186.755 83.925 187.215 ;
        RECT 84.110 186.765 84.440 186.935 ;
        RECT 84.620 186.765 85.370 186.935 ;
        RECT 83.660 185.635 83.940 186.235 ;
        RECT 84.110 185.235 84.280 186.765 ;
        RECT 84.450 186.265 85.030 186.595 ;
        RECT 84.450 185.395 84.690 186.265 ;
        RECT 85.200 185.985 85.370 186.765 ;
        RECT 85.620 186.715 85.990 187.215 ;
        RECT 86.170 186.765 86.630 186.935 ;
        RECT 86.860 186.765 87.530 186.935 ;
        RECT 86.170 186.535 86.340 186.765 ;
        RECT 85.540 186.235 86.340 186.535 ;
        RECT 86.510 186.265 87.060 186.595 ;
        RECT 85.540 186.205 85.710 186.235 ;
        RECT 85.830 185.985 86.000 186.055 ;
        RECT 85.200 185.815 86.000 185.985 ;
        RECT 85.490 185.725 86.000 185.815 ;
        RECT 84.880 185.290 85.320 185.645 ;
        RECT 83.660 184.665 83.925 185.125 ;
        RECT 84.110 184.860 84.345 185.235 ;
        RECT 85.490 185.110 85.660 185.725 ;
        RECT 84.590 184.940 85.660 185.110 ;
        RECT 85.830 184.665 86.000 185.465 ;
        RECT 86.170 185.165 86.340 186.235 ;
        RECT 86.510 185.335 86.700 186.055 ;
        RECT 86.870 185.725 87.060 186.265 ;
        RECT 87.360 186.225 87.530 186.765 ;
        RECT 87.845 186.685 88.015 187.215 ;
        RECT 88.310 186.565 88.670 187.005 ;
        RECT 88.845 186.735 89.015 187.215 ;
        RECT 89.205 186.570 89.540 186.995 ;
        RECT 89.715 186.740 89.885 187.215 ;
        RECT 90.060 186.570 90.395 186.995 ;
        RECT 90.565 186.740 90.735 187.215 ;
        RECT 88.310 186.395 88.810 186.565 ;
        RECT 89.205 186.400 90.875 186.570 ;
        RECT 91.045 186.465 92.255 187.215 ;
        RECT 88.640 186.225 88.810 186.395 ;
        RECT 87.360 186.055 88.450 186.225 ;
        RECT 88.640 186.055 90.460 186.225 ;
        RECT 86.870 185.395 87.190 185.725 ;
        RECT 86.170 184.835 86.420 185.165 ;
        RECT 87.360 185.135 87.530 186.055 ;
        RECT 88.640 185.800 88.810 186.055 ;
        RECT 90.630 185.835 90.875 186.400 ;
        RECT 87.700 185.630 88.810 185.800 ;
        RECT 89.205 185.665 90.875 185.835 ;
        RECT 91.045 185.755 91.565 186.295 ;
        RECT 91.735 185.925 92.255 186.465 ;
        RECT 87.700 185.470 88.560 185.630 ;
        RECT 86.645 184.965 87.530 185.135 ;
        RECT 87.710 184.665 87.925 185.165 ;
        RECT 88.390 184.845 88.560 185.470 ;
        RECT 88.845 184.665 89.025 185.445 ;
        RECT 89.205 184.905 89.540 185.665 ;
        RECT 89.720 184.665 89.890 185.495 ;
        RECT 90.060 184.905 90.390 185.665 ;
        RECT 90.560 184.665 90.730 185.495 ;
        RECT 91.045 184.665 92.255 185.755 ;
        RECT 18.280 184.495 92.340 184.665 ;
        RECT 18.365 183.405 19.575 184.495 ;
        RECT 19.745 184.060 25.090 184.495 ;
        RECT 18.365 182.695 18.885 183.235 ;
        RECT 19.055 182.865 19.575 183.405 ;
        RECT 18.365 181.945 19.575 182.695 ;
        RECT 21.330 182.490 21.670 183.320 ;
        RECT 23.150 182.810 23.500 184.060 ;
        RECT 25.265 183.405 26.935 184.495 ;
        RECT 25.265 182.715 26.015 183.235 ;
        RECT 26.185 182.885 26.935 183.405 ;
        RECT 27.115 183.545 27.390 184.315 ;
        RECT 27.560 183.885 27.890 184.315 ;
        RECT 28.060 184.055 28.255 184.495 ;
        RECT 28.435 183.885 28.765 184.315 ;
        RECT 27.560 183.715 28.765 183.885 ;
        RECT 27.115 183.355 27.700 183.545 ;
        RECT 27.870 183.385 28.765 183.715 ;
        RECT 28.945 183.355 29.225 184.495 ;
        RECT 19.745 181.945 25.090 182.490 ;
        RECT 25.265 181.945 26.935 182.715 ;
        RECT 27.115 182.535 27.355 183.185 ;
        RECT 27.525 182.685 27.700 183.355 ;
        RECT 29.395 183.345 29.725 184.325 ;
        RECT 29.895 183.355 30.155 184.495 ;
        RECT 27.870 182.855 28.285 183.185 ;
        RECT 28.465 182.855 28.760 183.185 ;
        RECT 28.955 182.915 29.290 183.185 ;
        RECT 27.525 182.505 27.855 182.685 ;
        RECT 27.130 181.945 27.460 182.335 ;
        RECT 27.630 182.125 27.855 182.505 ;
        RECT 28.055 182.235 28.285 182.855 ;
        RECT 29.460 182.745 29.630 183.345 ;
        RECT 31.245 183.330 31.535 184.495 ;
        RECT 31.795 183.750 32.065 184.495 ;
        RECT 32.695 184.490 38.970 184.495 ;
        RECT 32.235 183.580 32.525 184.320 ;
        RECT 32.695 183.765 32.950 184.490 ;
        RECT 33.135 183.595 33.395 184.320 ;
        RECT 33.565 183.765 33.810 184.490 ;
        RECT 33.995 183.595 34.255 184.320 ;
        RECT 34.425 183.765 34.670 184.490 ;
        RECT 34.855 183.595 35.115 184.320 ;
        RECT 35.285 183.765 35.530 184.490 ;
        RECT 35.700 183.595 35.960 184.320 ;
        RECT 36.130 183.765 36.390 184.490 ;
        RECT 36.560 183.595 36.820 184.320 ;
        RECT 36.990 183.765 37.250 184.490 ;
        RECT 37.420 183.595 37.680 184.320 ;
        RECT 37.850 183.765 38.110 184.490 ;
        RECT 38.280 183.595 38.540 184.320 ;
        RECT 38.710 183.695 38.970 184.490 ;
        RECT 33.135 183.580 38.540 183.595 ;
        RECT 31.795 183.355 38.540 183.580 ;
        RECT 29.800 182.935 30.135 183.185 ;
        RECT 31.795 182.765 32.960 183.355 ;
        RECT 39.140 183.185 39.390 184.320 ;
        RECT 39.570 183.685 39.830 184.495 ;
        RECT 40.005 183.185 40.250 184.325 ;
        RECT 40.430 183.685 40.725 184.495 ;
        RECT 40.905 183.775 41.365 184.325 ;
        RECT 41.555 183.775 41.885 184.495 ;
        RECT 33.130 182.935 40.250 183.185 ;
        RECT 28.465 181.945 28.765 182.675 ;
        RECT 28.945 181.945 29.255 182.745 ;
        RECT 29.460 182.115 30.155 182.745 ;
        RECT 31.245 181.945 31.535 182.670 ;
        RECT 31.795 182.595 38.540 182.765 ;
        RECT 31.795 181.945 32.095 182.425 ;
        RECT 32.265 182.140 32.525 182.595 ;
        RECT 32.695 181.945 32.955 182.425 ;
        RECT 33.135 182.140 33.395 182.595 ;
        RECT 33.565 181.945 33.815 182.425 ;
        RECT 33.995 182.140 34.255 182.595 ;
        RECT 34.425 181.945 34.675 182.425 ;
        RECT 34.855 182.140 35.115 182.595 ;
        RECT 35.285 181.945 35.530 182.425 ;
        RECT 35.700 182.140 35.975 182.595 ;
        RECT 36.145 181.945 36.390 182.425 ;
        RECT 36.560 182.140 36.820 182.595 ;
        RECT 36.990 181.945 37.250 182.425 ;
        RECT 37.420 182.140 37.680 182.595 ;
        RECT 37.850 181.945 38.110 182.425 ;
        RECT 38.280 182.140 38.540 182.595 ;
        RECT 38.710 181.945 38.970 182.505 ;
        RECT 39.140 182.125 39.390 182.935 ;
        RECT 39.570 181.945 39.830 182.470 ;
        RECT 40.000 182.125 40.250 182.935 ;
        RECT 40.420 182.625 40.735 183.185 ;
        RECT 40.430 181.945 40.735 182.455 ;
        RECT 40.905 182.405 41.155 183.775 ;
        RECT 42.085 183.605 42.385 184.155 ;
        RECT 42.555 183.825 42.835 184.495 ;
        RECT 41.445 183.435 42.385 183.605 ;
        RECT 41.445 183.185 41.615 183.435 ;
        RECT 42.755 183.185 43.020 183.545 ;
        RECT 43.390 183.525 43.780 183.700 ;
        RECT 44.265 183.695 44.595 184.495 ;
        RECT 44.765 183.705 45.300 184.325 ;
        RECT 45.705 183.825 45.985 184.495 ;
        RECT 43.390 183.355 44.815 183.525 ;
        RECT 41.325 182.855 41.615 183.185 ;
        RECT 41.785 182.935 42.125 183.185 ;
        RECT 42.345 182.935 43.020 183.185 ;
        RECT 41.445 182.765 41.615 182.855 ;
        RECT 41.445 182.575 42.835 182.765 ;
        RECT 43.265 182.625 43.620 183.185 ;
        RECT 40.905 182.115 41.465 182.405 ;
        RECT 41.635 181.945 41.885 182.405 ;
        RECT 42.505 182.215 42.835 182.575 ;
        RECT 43.790 182.455 43.960 183.355 ;
        RECT 44.130 182.625 44.395 183.185 ;
        RECT 44.645 182.855 44.815 183.355 ;
        RECT 44.985 182.685 45.300 183.705 ;
        RECT 46.155 183.605 46.455 184.155 ;
        RECT 46.655 183.775 46.985 184.495 ;
        RECT 47.175 183.775 47.635 184.325 ;
        RECT 45.520 183.185 45.785 183.545 ;
        RECT 46.155 183.435 47.095 183.605 ;
        RECT 46.925 183.185 47.095 183.435 ;
        RECT 45.520 182.935 46.195 183.185 ;
        RECT 46.415 182.935 46.755 183.185 ;
        RECT 46.925 182.855 47.215 183.185 ;
        RECT 46.925 182.765 47.095 182.855 ;
        RECT 43.370 181.945 43.610 182.455 ;
        RECT 43.790 182.125 44.070 182.455 ;
        RECT 44.300 181.945 44.515 182.455 ;
        RECT 44.685 182.115 45.300 182.685 ;
        RECT 45.705 182.575 47.095 182.765 ;
        RECT 45.705 182.215 46.035 182.575 ;
        RECT 47.385 182.405 47.635 183.775 ;
        RECT 46.655 181.945 46.905 182.405 ;
        RECT 47.075 182.115 47.635 182.405 ;
        RECT 47.810 183.775 48.145 184.285 ;
        RECT 47.810 182.420 48.065 183.775 ;
        RECT 48.395 183.695 48.725 184.495 ;
        RECT 48.970 183.905 49.255 184.325 ;
        RECT 49.510 184.075 49.840 184.495 ;
        RECT 50.065 184.155 51.225 184.325 ;
        RECT 50.065 183.905 50.395 184.155 ;
        RECT 48.970 183.735 50.395 183.905 ;
        RECT 50.625 183.525 50.795 183.985 ;
        RECT 51.055 183.655 51.225 184.155 ;
        RECT 48.425 183.355 50.795 183.525 ;
        RECT 48.425 183.185 48.595 183.355 ;
        RECT 51.045 183.185 51.250 183.475 ;
        RECT 51.485 183.405 54.995 184.495 ;
        RECT 48.290 182.855 48.595 183.185 ;
        RECT 48.790 183.135 49.040 183.185 ;
        RECT 48.785 182.965 49.040 183.135 ;
        RECT 48.790 182.855 49.040 182.965 ;
        RECT 48.425 182.685 48.595 182.855 ;
        RECT 49.250 182.795 49.520 183.185 ;
        RECT 49.710 182.795 50.000 183.185 ;
        RECT 48.425 182.515 48.985 182.685 ;
        RECT 49.245 182.625 49.520 182.795 ;
        RECT 49.705 182.625 50.000 182.795 ;
        RECT 49.250 182.525 49.520 182.625 ;
        RECT 49.710 182.525 50.000 182.625 ;
        RECT 50.170 182.520 50.590 183.185 ;
        RECT 50.900 183.135 51.250 183.185 ;
        RECT 50.900 182.965 51.255 183.135 ;
        RECT 50.900 182.855 51.250 182.965 ;
        RECT 51.485 182.715 53.135 183.235 ;
        RECT 53.305 182.885 54.995 183.405 ;
        RECT 55.685 183.355 55.895 184.495 ;
        RECT 56.065 183.345 56.395 184.325 ;
        RECT 56.565 183.355 56.795 184.495 ;
        RECT 47.810 182.160 48.145 182.420 ;
        RECT 48.815 182.345 48.985 182.515 ;
        RECT 48.315 181.945 48.645 182.345 ;
        RECT 48.815 182.175 50.430 182.345 ;
        RECT 50.975 181.945 51.305 182.665 ;
        RECT 51.485 181.945 54.995 182.715 ;
        RECT 55.685 181.945 55.895 182.765 ;
        RECT 56.065 182.745 56.315 183.345 ;
        RECT 57.005 183.330 57.295 184.495 ;
        RECT 57.475 183.685 57.770 184.495 ;
        RECT 57.950 183.185 58.195 184.325 ;
        RECT 58.370 183.685 58.630 184.495 ;
        RECT 59.230 184.490 65.505 184.495 ;
        RECT 58.810 183.185 59.060 184.320 ;
        RECT 59.230 183.695 59.490 184.490 ;
        RECT 59.660 183.595 59.920 184.320 ;
        RECT 60.090 183.765 60.350 184.490 ;
        RECT 60.520 183.595 60.780 184.320 ;
        RECT 60.950 183.765 61.210 184.490 ;
        RECT 61.380 183.595 61.640 184.320 ;
        RECT 61.810 183.765 62.070 184.490 ;
        RECT 62.240 183.595 62.500 184.320 ;
        RECT 62.670 183.765 62.915 184.490 ;
        RECT 63.085 183.595 63.345 184.320 ;
        RECT 63.530 183.765 63.775 184.490 ;
        RECT 63.945 183.595 64.205 184.320 ;
        RECT 64.390 183.765 64.635 184.490 ;
        RECT 64.805 183.595 65.065 184.320 ;
        RECT 65.250 183.765 65.505 184.490 ;
        RECT 59.660 183.580 65.065 183.595 ;
        RECT 65.675 183.580 65.965 184.320 ;
        RECT 66.135 183.750 66.405 184.495 ;
        RECT 59.660 183.355 66.405 183.580 ;
        RECT 66.665 183.405 67.875 184.495 ;
        RECT 56.485 182.935 56.815 183.185 ;
        RECT 56.065 182.115 56.395 182.745 ;
        RECT 56.565 181.945 56.795 182.765 ;
        RECT 57.005 181.945 57.295 182.670 ;
        RECT 57.465 182.625 57.780 183.185 ;
        RECT 57.950 182.935 65.070 183.185 ;
        RECT 57.465 181.945 57.770 182.455 ;
        RECT 57.950 182.125 58.200 182.935 ;
        RECT 58.370 181.945 58.630 182.470 ;
        RECT 58.810 182.125 59.060 182.935 ;
        RECT 65.240 182.765 66.405 183.355 ;
        RECT 59.660 182.595 66.405 182.765 ;
        RECT 66.665 182.695 67.185 183.235 ;
        RECT 67.355 182.865 67.875 183.405 ;
        RECT 68.045 183.355 68.385 184.325 ;
        RECT 68.555 183.355 68.725 184.495 ;
        RECT 68.995 183.695 69.245 184.495 ;
        RECT 69.890 183.525 70.220 184.325 ;
        RECT 70.520 183.695 70.850 184.495 ;
        RECT 71.020 183.525 71.350 184.325 ;
        RECT 68.915 183.355 71.350 183.525 ;
        RECT 71.725 183.525 72.035 184.325 ;
        RECT 72.205 183.695 72.515 184.495 ;
        RECT 72.685 183.865 72.945 184.325 ;
        RECT 73.115 184.035 73.370 184.495 ;
        RECT 73.545 183.865 73.805 184.325 ;
        RECT 72.685 183.695 73.805 183.865 ;
        RECT 71.725 183.355 72.755 183.525 ;
        RECT 68.045 182.745 68.220 183.355 ;
        RECT 68.915 183.105 69.085 183.355 ;
        RECT 68.390 182.935 69.085 183.105 ;
        RECT 69.260 182.935 69.680 183.135 ;
        RECT 69.850 182.935 70.180 183.135 ;
        RECT 70.350 182.935 70.680 183.135 ;
        RECT 59.230 181.945 59.490 182.505 ;
        RECT 59.660 182.140 59.920 182.595 ;
        RECT 60.090 181.945 60.350 182.425 ;
        RECT 60.520 182.140 60.780 182.595 ;
        RECT 60.950 181.945 61.210 182.425 ;
        RECT 61.380 182.140 61.640 182.595 ;
        RECT 61.810 181.945 62.055 182.425 ;
        RECT 62.225 182.140 62.500 182.595 ;
        RECT 62.670 181.945 62.915 182.425 ;
        RECT 63.085 182.140 63.345 182.595 ;
        RECT 63.525 181.945 63.775 182.425 ;
        RECT 63.945 182.140 64.205 182.595 ;
        RECT 64.385 181.945 64.635 182.425 ;
        RECT 64.805 182.140 65.065 182.595 ;
        RECT 65.245 181.945 65.505 182.425 ;
        RECT 65.675 182.140 65.935 182.595 ;
        RECT 66.105 181.945 66.405 182.425 ;
        RECT 66.665 181.945 67.875 182.695 ;
        RECT 68.045 182.115 68.385 182.745 ;
        RECT 68.555 181.945 68.805 182.745 ;
        RECT 68.995 182.595 70.220 182.765 ;
        RECT 68.995 182.115 69.325 182.595 ;
        RECT 69.495 181.945 69.720 182.405 ;
        RECT 69.890 182.115 70.220 182.595 ;
        RECT 70.850 182.725 71.020 183.355 ;
        RECT 71.205 182.935 71.555 183.185 ;
        RECT 70.850 182.115 71.350 182.725 ;
        RECT 71.725 182.445 71.895 183.355 ;
        RECT 72.065 182.615 72.415 183.185 ;
        RECT 72.585 183.105 72.755 183.355 ;
        RECT 73.545 183.445 73.805 183.695 ;
        RECT 73.975 183.625 74.260 184.495 ;
        RECT 74.485 184.060 79.830 184.495 ;
        RECT 73.545 183.275 74.300 183.445 ;
        RECT 72.585 182.935 73.725 183.105 ;
        RECT 73.895 182.765 74.300 183.275 ;
        RECT 72.650 182.595 74.300 182.765 ;
        RECT 71.725 182.115 72.025 182.445 ;
        RECT 72.195 181.945 72.470 182.425 ;
        RECT 72.650 182.205 72.945 182.595 ;
        RECT 73.115 181.945 73.370 182.425 ;
        RECT 73.545 182.205 73.805 182.595 ;
        RECT 76.070 182.490 76.410 183.320 ;
        RECT 77.890 182.810 78.240 184.060 ;
        RECT 73.975 181.945 74.255 182.425 ;
        RECT 74.485 181.945 79.830 182.490 ;
        RECT 80.015 182.125 80.275 184.315 ;
        RECT 80.445 183.765 80.785 184.495 ;
        RECT 80.965 183.585 81.235 184.315 ;
        RECT 80.465 183.365 81.235 183.585 ;
        RECT 81.415 183.605 81.645 184.315 ;
        RECT 81.815 183.785 82.145 184.495 ;
        RECT 82.315 183.605 82.575 184.315 ;
        RECT 81.415 183.365 82.575 183.605 ;
        RECT 80.465 182.695 80.755 183.365 ;
        RECT 82.765 183.330 83.055 184.495 ;
        RECT 83.225 183.355 83.565 184.325 ;
        RECT 83.735 183.355 83.905 184.495 ;
        RECT 84.175 183.695 84.425 184.495 ;
        RECT 85.070 183.525 85.400 184.325 ;
        RECT 85.700 183.695 86.030 184.495 ;
        RECT 86.200 183.525 86.530 184.325 ;
        RECT 84.095 183.355 86.530 183.525 ;
        RECT 86.905 183.625 87.180 184.325 ;
        RECT 87.350 183.950 87.605 184.495 ;
        RECT 87.775 183.985 88.255 184.325 ;
        RECT 88.430 183.940 89.035 184.495 ;
        RECT 88.420 183.840 89.035 183.940 ;
        RECT 88.420 183.815 88.605 183.840 ;
        RECT 80.935 182.875 81.400 183.185 ;
        RECT 81.580 182.875 82.105 183.185 ;
        RECT 80.465 182.495 81.695 182.695 ;
        RECT 80.535 181.945 81.205 182.315 ;
        RECT 81.385 182.125 81.695 182.495 ;
        RECT 81.875 182.235 82.105 182.875 ;
        RECT 82.285 182.855 82.585 183.185 ;
        RECT 83.225 182.745 83.400 183.355 ;
        RECT 84.095 183.105 84.265 183.355 ;
        RECT 83.570 182.935 84.265 183.105 ;
        RECT 84.440 182.935 84.860 183.135 ;
        RECT 85.030 182.935 85.360 183.135 ;
        RECT 85.530 182.935 85.860 183.135 ;
        RECT 82.285 181.945 82.575 182.675 ;
        RECT 82.765 181.945 83.055 182.670 ;
        RECT 83.225 182.115 83.565 182.745 ;
        RECT 83.735 181.945 83.985 182.745 ;
        RECT 84.175 182.595 85.400 182.765 ;
        RECT 84.175 182.115 84.505 182.595 ;
        RECT 84.675 181.945 84.900 182.405 ;
        RECT 85.070 182.115 85.400 182.595 ;
        RECT 86.030 182.725 86.200 183.355 ;
        RECT 86.385 182.935 86.735 183.185 ;
        RECT 86.030 182.115 86.530 182.725 ;
        RECT 86.905 182.595 87.075 183.625 ;
        RECT 87.350 183.495 88.105 183.745 ;
        RECT 88.275 183.570 88.605 183.815 ;
        RECT 87.350 183.460 88.120 183.495 ;
        RECT 87.350 183.450 88.135 183.460 ;
        RECT 87.245 183.435 88.140 183.450 ;
        RECT 87.245 183.420 88.160 183.435 ;
        RECT 87.245 183.410 88.180 183.420 ;
        RECT 87.245 183.400 88.205 183.410 ;
        RECT 87.245 183.370 88.275 183.400 ;
        RECT 87.245 183.340 88.295 183.370 ;
        RECT 87.245 183.310 88.315 183.340 ;
        RECT 87.245 183.285 88.345 183.310 ;
        RECT 87.245 183.250 88.380 183.285 ;
        RECT 87.245 183.245 88.410 183.250 ;
        RECT 87.245 182.850 87.475 183.245 ;
        RECT 88.020 183.240 88.410 183.245 ;
        RECT 88.045 183.230 88.410 183.240 ;
        RECT 88.060 183.225 88.410 183.230 ;
        RECT 88.075 183.220 88.410 183.225 ;
        RECT 88.775 183.220 89.035 183.670 ;
        RECT 89.205 183.405 90.875 184.495 ;
        RECT 88.075 183.215 89.035 183.220 ;
        RECT 88.085 183.205 89.035 183.215 ;
        RECT 88.095 183.200 89.035 183.205 ;
        RECT 88.105 183.190 89.035 183.200 ;
        RECT 88.110 183.180 89.035 183.190 ;
        RECT 88.115 183.175 89.035 183.180 ;
        RECT 88.125 183.160 89.035 183.175 ;
        RECT 88.130 183.145 89.035 183.160 ;
        RECT 88.140 183.120 89.035 183.145 ;
        RECT 87.645 182.650 87.975 183.075 ;
        RECT 86.905 182.115 87.165 182.595 ;
        RECT 87.335 181.945 87.585 182.485 ;
        RECT 87.755 182.165 87.975 182.650 ;
        RECT 88.145 183.050 89.035 183.120 ;
        RECT 88.145 182.325 88.315 183.050 ;
        RECT 88.485 182.495 89.035 182.880 ;
        RECT 89.205 182.715 89.955 183.235 ;
        RECT 90.125 182.885 90.875 183.405 ;
        RECT 91.045 183.405 92.255 184.495 ;
        RECT 91.045 182.865 91.565 183.405 ;
        RECT 88.145 182.155 89.035 182.325 ;
        RECT 89.205 181.945 90.875 182.715 ;
        RECT 91.735 182.695 92.255 183.235 ;
        RECT 91.045 181.945 92.255 182.695 ;
        RECT 18.280 181.775 92.340 181.945 ;
        RECT 18.365 181.025 19.575 181.775 ;
        RECT 19.745 181.230 25.090 181.775 ;
        RECT 25.265 181.230 30.610 181.775 ;
        RECT 30.785 181.230 36.130 181.775 ;
        RECT 18.365 180.485 18.885 181.025 ;
        RECT 19.055 180.315 19.575 180.855 ;
        RECT 21.330 180.400 21.670 181.230 ;
        RECT 18.365 179.225 19.575 180.315 ;
        RECT 23.150 179.660 23.500 180.910 ;
        RECT 26.850 180.400 27.190 181.230 ;
        RECT 28.670 179.660 29.020 180.910 ;
        RECT 32.370 180.400 32.710 181.230 ;
        RECT 37.225 181.125 37.485 181.605 ;
        RECT 37.655 181.235 37.905 181.775 ;
        RECT 34.190 179.660 34.540 180.910 ;
        RECT 37.225 180.095 37.395 181.125 ;
        RECT 38.075 181.070 38.295 181.555 ;
        RECT 37.565 180.475 37.795 180.870 ;
        RECT 37.965 180.645 38.295 181.070 ;
        RECT 38.465 181.395 39.355 181.565 ;
        RECT 38.465 180.670 38.635 181.395 ;
        RECT 38.805 180.840 39.355 181.225 ;
        RECT 39.525 181.005 41.195 181.775 ;
        RECT 38.465 180.600 39.355 180.670 ;
        RECT 38.460 180.575 39.355 180.600 ;
        RECT 38.450 180.560 39.355 180.575 ;
        RECT 38.445 180.545 39.355 180.560 ;
        RECT 38.435 180.540 39.355 180.545 ;
        RECT 38.430 180.530 39.355 180.540 ;
        RECT 38.425 180.520 39.355 180.530 ;
        RECT 38.415 180.515 39.355 180.520 ;
        RECT 38.405 180.505 39.355 180.515 ;
        RECT 38.395 180.500 39.355 180.505 ;
        RECT 38.395 180.495 38.730 180.500 ;
        RECT 38.380 180.490 38.730 180.495 ;
        RECT 38.365 180.480 38.730 180.490 ;
        RECT 38.340 180.475 38.730 180.480 ;
        RECT 37.565 180.470 38.730 180.475 ;
        RECT 37.565 180.435 38.700 180.470 ;
        RECT 37.565 180.410 38.665 180.435 ;
        RECT 37.565 180.380 38.635 180.410 ;
        RECT 37.565 180.350 38.615 180.380 ;
        RECT 37.565 180.320 38.595 180.350 ;
        RECT 37.565 180.310 38.525 180.320 ;
        RECT 37.565 180.300 38.500 180.310 ;
        RECT 37.565 180.285 38.480 180.300 ;
        RECT 37.565 180.270 38.460 180.285 ;
        RECT 37.670 180.260 38.455 180.270 ;
        RECT 37.670 180.225 38.440 180.260 ;
        RECT 19.745 179.225 25.090 179.660 ;
        RECT 25.265 179.225 30.610 179.660 ;
        RECT 30.785 179.225 36.130 179.660 ;
        RECT 37.225 179.395 37.500 180.095 ;
        RECT 37.670 179.975 38.425 180.225 ;
        RECT 38.595 179.905 38.925 180.150 ;
        RECT 39.095 180.050 39.355 180.500 ;
        RECT 39.525 180.485 40.275 181.005 ;
        RECT 41.825 180.975 42.520 181.605 ;
        RECT 42.725 180.975 43.035 181.775 ;
        RECT 44.125 181.050 44.415 181.775 ;
        RECT 44.585 181.230 49.930 181.775 ;
        RECT 50.105 181.230 55.450 181.775 ;
        RECT 40.445 180.315 41.195 180.835 ;
        RECT 41.845 180.535 42.180 180.785 ;
        RECT 42.350 180.375 42.520 180.975 ;
        RECT 42.690 180.535 43.025 180.805 ;
        RECT 46.170 180.400 46.510 181.230 ;
        RECT 38.740 179.880 38.925 179.905 ;
        RECT 38.740 179.780 39.355 179.880 ;
        RECT 37.670 179.225 37.925 179.770 ;
        RECT 38.095 179.395 38.575 179.735 ;
        RECT 38.750 179.225 39.355 179.780 ;
        RECT 39.525 179.225 41.195 180.315 ;
        RECT 41.825 179.225 42.085 180.365 ;
        RECT 42.255 179.395 42.585 180.375 ;
        RECT 42.755 179.225 43.035 180.365 ;
        RECT 44.125 179.225 44.415 180.390 ;
        RECT 47.990 179.660 48.340 180.910 ;
        RECT 51.690 180.400 52.030 181.230 ;
        RECT 55.625 181.005 58.215 181.775 ;
        RECT 58.385 181.315 58.945 181.605 ;
        RECT 59.115 181.315 59.365 181.775 ;
        RECT 53.510 179.660 53.860 180.910 ;
        RECT 55.625 180.485 56.835 181.005 ;
        RECT 57.005 180.315 58.215 180.835 ;
        RECT 44.585 179.225 49.930 179.660 ;
        RECT 50.105 179.225 55.450 179.660 ;
        RECT 55.625 179.225 58.215 180.315 ;
        RECT 58.385 179.945 58.635 181.315 ;
        RECT 59.985 181.145 60.315 181.505 ;
        RECT 58.925 180.955 60.315 181.145 ;
        RECT 60.685 180.975 61.380 181.605 ;
        RECT 61.585 180.975 61.895 181.775 ;
        RECT 62.065 181.275 62.365 181.605 ;
        RECT 62.535 181.295 62.810 181.775 ;
        RECT 58.925 180.865 59.095 180.955 ;
        RECT 58.805 180.535 59.095 180.865 ;
        RECT 59.265 180.535 59.605 180.785 ;
        RECT 59.825 180.535 60.500 180.785 ;
        RECT 60.705 180.535 61.040 180.785 ;
        RECT 58.925 180.285 59.095 180.535 ;
        RECT 58.925 180.115 59.865 180.285 ;
        RECT 60.235 180.175 60.500 180.535 ;
        RECT 61.210 180.375 61.380 180.975 ;
        RECT 61.550 180.535 61.885 180.805 ;
        RECT 58.385 179.395 58.845 179.945 ;
        RECT 59.035 179.225 59.365 179.945 ;
        RECT 59.565 179.565 59.865 180.115 ;
        RECT 60.035 179.225 60.315 179.895 ;
        RECT 60.685 179.225 60.945 180.365 ;
        RECT 61.115 179.395 61.445 180.375 ;
        RECT 62.065 180.365 62.235 181.275 ;
        RECT 62.990 181.125 63.285 181.515 ;
        RECT 63.455 181.295 63.710 181.775 ;
        RECT 63.885 181.125 64.145 181.515 ;
        RECT 64.315 181.295 64.595 181.775 ;
        RECT 62.405 180.535 62.755 181.105 ;
        RECT 62.990 180.955 64.640 181.125 ;
        RECT 62.925 180.615 64.065 180.785 ;
        RECT 62.925 180.365 63.095 180.615 ;
        RECT 64.235 180.445 64.640 180.955 ;
        RECT 64.825 181.005 68.335 181.775 ;
        RECT 68.505 181.025 69.715 181.775 ;
        RECT 69.885 181.050 70.175 181.775 ;
        RECT 71.595 181.375 71.925 181.775 ;
        RECT 72.095 181.205 72.425 181.545 ;
        RECT 73.475 181.375 73.805 181.775 ;
        RECT 71.440 181.035 73.805 181.205 ;
        RECT 73.975 181.050 74.305 181.560 ;
        RECT 74.485 181.230 79.830 181.775 ;
        RECT 80.005 181.230 85.350 181.775 ;
        RECT 85.525 181.230 90.870 181.775 ;
        RECT 64.825 180.485 66.475 181.005 ;
        RECT 61.615 179.225 61.895 180.365 ;
        RECT 62.065 180.195 63.095 180.365 ;
        RECT 63.885 180.275 64.640 180.445 ;
        RECT 66.645 180.315 68.335 180.835 ;
        RECT 68.505 180.485 69.025 181.025 ;
        RECT 69.195 180.315 69.715 180.855 ;
        RECT 62.065 179.395 62.375 180.195 ;
        RECT 63.885 180.025 64.145 180.275 ;
        RECT 62.545 179.225 62.855 180.025 ;
        RECT 63.025 179.855 64.145 180.025 ;
        RECT 63.025 179.395 63.285 179.855 ;
        RECT 63.455 179.225 63.710 179.685 ;
        RECT 63.885 179.395 64.145 179.855 ;
        RECT 64.315 179.225 64.600 180.095 ;
        RECT 64.825 179.225 68.335 180.315 ;
        RECT 68.505 179.225 69.715 180.315 ;
        RECT 69.885 179.225 70.175 180.390 ;
        RECT 71.440 180.035 71.610 181.035 ;
        RECT 73.635 180.865 73.805 181.035 ;
        RECT 71.780 180.205 72.025 180.865 ;
        RECT 72.240 180.205 72.505 180.865 ;
        RECT 72.700 180.205 72.985 180.865 ;
        RECT 73.160 180.535 73.465 180.865 ;
        RECT 73.635 180.535 73.945 180.865 ;
        RECT 73.160 180.205 73.375 180.535 ;
        RECT 71.440 179.865 71.895 180.035 ;
        RECT 71.565 179.435 71.895 179.865 ;
        RECT 72.075 179.865 73.365 180.035 ;
        RECT 72.075 179.445 72.325 179.865 ;
        RECT 72.555 179.225 72.885 179.695 ;
        RECT 73.115 179.445 73.365 179.865 ;
        RECT 73.555 179.225 73.805 180.365 ;
        RECT 74.115 180.285 74.305 181.050 ;
        RECT 76.070 180.400 76.410 181.230 ;
        RECT 73.975 179.435 74.305 180.285 ;
        RECT 77.890 179.660 78.240 180.910 ;
        RECT 81.590 180.400 81.930 181.230 ;
        RECT 83.410 179.660 83.760 180.910 ;
        RECT 87.110 180.400 87.450 181.230 ;
        RECT 91.045 181.025 92.255 181.775 ;
        RECT 88.930 179.660 89.280 180.910 ;
        RECT 91.045 180.315 91.565 180.855 ;
        RECT 91.735 180.485 92.255 181.025 ;
        RECT 74.485 179.225 79.830 179.660 ;
        RECT 80.005 179.225 85.350 179.660 ;
        RECT 85.525 179.225 90.870 179.660 ;
        RECT 91.045 179.225 92.255 180.315 ;
        RECT 18.280 179.055 92.340 179.225 ;
        RECT 18.365 177.965 19.575 179.055 ;
        RECT 19.745 177.965 23.255 179.055 ;
        RECT 23.975 178.385 24.145 178.885 ;
        RECT 24.315 178.555 24.645 179.055 ;
        RECT 23.975 178.215 24.640 178.385 ;
        RECT 18.365 177.255 18.885 177.795 ;
        RECT 19.055 177.425 19.575 177.965 ;
        RECT 19.745 177.275 21.395 177.795 ;
        RECT 21.565 177.445 23.255 177.965 ;
        RECT 23.890 177.395 24.240 178.045 ;
        RECT 18.365 176.505 19.575 177.255 ;
        RECT 19.745 176.505 23.255 177.275 ;
        RECT 24.410 177.225 24.640 178.215 ;
        RECT 23.975 177.055 24.640 177.225 ;
        RECT 23.975 176.765 24.145 177.055 ;
        RECT 24.315 176.505 24.645 176.885 ;
        RECT 24.815 176.765 25.000 178.885 ;
        RECT 25.240 178.595 25.505 179.055 ;
        RECT 25.675 178.460 25.925 178.885 ;
        RECT 26.135 178.610 27.240 178.780 ;
        RECT 25.620 178.330 25.925 178.460 ;
        RECT 25.170 177.135 25.450 178.085 ;
        RECT 25.620 177.225 25.790 178.330 ;
        RECT 25.960 177.545 26.200 178.140 ;
        RECT 26.370 178.075 26.900 178.440 ;
        RECT 26.370 177.375 26.540 178.075 ;
        RECT 27.070 177.995 27.240 178.610 ;
        RECT 27.410 178.255 27.580 179.055 ;
        RECT 27.750 178.555 28.000 178.885 ;
        RECT 28.225 178.585 29.110 178.755 ;
        RECT 27.070 177.905 27.580 177.995 ;
        RECT 25.620 177.095 25.845 177.225 ;
        RECT 26.015 177.155 26.540 177.375 ;
        RECT 26.710 177.735 27.580 177.905 ;
        RECT 25.255 176.505 25.505 176.965 ;
        RECT 25.675 176.955 25.845 177.095 ;
        RECT 26.710 176.955 26.880 177.735 ;
        RECT 27.410 177.665 27.580 177.735 ;
        RECT 27.090 177.485 27.290 177.515 ;
        RECT 27.750 177.485 27.920 178.555 ;
        RECT 28.090 177.665 28.280 178.385 ;
        RECT 27.090 177.185 27.920 177.485 ;
        RECT 28.450 177.455 28.770 178.415 ;
        RECT 25.675 176.785 26.010 176.955 ;
        RECT 26.205 176.785 26.880 176.955 ;
        RECT 27.200 176.505 27.570 177.005 ;
        RECT 27.750 176.955 27.920 177.185 ;
        RECT 28.305 177.125 28.770 177.455 ;
        RECT 28.940 177.745 29.110 178.585 ;
        RECT 29.290 178.555 29.605 179.055 ;
        RECT 29.835 178.325 30.175 178.885 ;
        RECT 29.280 177.950 30.175 178.325 ;
        RECT 30.345 178.045 30.515 179.055 ;
        RECT 29.985 177.745 30.175 177.950 ;
        RECT 30.685 177.995 31.015 178.840 ;
        RECT 30.685 177.915 31.075 177.995 ;
        RECT 30.860 177.865 31.075 177.915 ;
        RECT 31.245 177.890 31.535 179.055 ;
        RECT 31.705 177.915 32.090 178.875 ;
        RECT 32.305 178.255 32.595 179.055 ;
        RECT 32.765 178.715 34.130 178.885 ;
        RECT 32.765 178.085 32.935 178.715 ;
        RECT 32.260 177.915 32.935 178.085 ;
        RECT 28.940 177.415 29.815 177.745 ;
        RECT 29.985 177.415 30.735 177.745 ;
        RECT 28.940 176.955 29.110 177.415 ;
        RECT 29.985 177.245 30.185 177.415 ;
        RECT 30.905 177.285 31.075 177.865 ;
        RECT 30.850 177.245 31.075 177.285 ;
        RECT 27.750 176.785 28.155 176.955 ;
        RECT 28.325 176.785 29.110 176.955 ;
        RECT 29.385 176.505 29.595 177.035 ;
        RECT 29.855 176.720 30.185 177.245 ;
        RECT 30.695 177.160 31.075 177.245 ;
        RECT 31.705 177.245 31.880 177.915 ;
        RECT 32.260 177.745 32.430 177.915 ;
        RECT 33.105 177.745 33.430 178.545 ;
        RECT 33.800 178.505 34.130 178.715 ;
        RECT 33.800 178.255 34.755 178.505 ;
        RECT 32.065 177.495 32.430 177.745 ;
        RECT 32.625 177.495 32.875 177.745 ;
        RECT 32.065 177.415 32.255 177.495 ;
        RECT 32.625 177.415 32.795 177.495 ;
        RECT 33.085 177.415 33.430 177.745 ;
        RECT 33.600 177.415 33.875 178.080 ;
        RECT 34.060 177.415 34.415 178.080 ;
        RECT 34.585 177.245 34.755 178.255 ;
        RECT 34.925 177.915 35.215 179.055 ;
        RECT 35.500 178.425 35.785 178.885 ;
        RECT 35.955 178.595 36.225 179.055 ;
        RECT 35.500 178.205 36.455 178.425 ;
        RECT 34.940 177.415 35.215 177.745 ;
        RECT 35.385 177.475 36.075 178.035 ;
        RECT 36.245 177.305 36.455 178.205 ;
        RECT 30.355 176.505 30.525 177.115 ;
        RECT 30.695 176.725 31.025 177.160 ;
        RECT 31.245 176.505 31.535 177.230 ;
        RECT 31.705 176.675 32.215 177.245 ;
        RECT 32.760 177.075 34.160 177.245 ;
        RECT 32.385 176.505 32.555 177.065 ;
        RECT 32.760 176.675 33.090 177.075 ;
        RECT 33.265 176.505 33.595 176.905 ;
        RECT 33.830 176.885 34.160 177.075 ;
        RECT 34.330 177.055 34.755 177.245 ;
        RECT 34.925 176.885 35.215 177.155 ;
        RECT 33.830 176.675 35.215 176.885 ;
        RECT 35.500 177.135 36.455 177.305 ;
        RECT 36.625 178.035 37.025 178.885 ;
        RECT 37.215 178.425 37.495 178.885 ;
        RECT 38.015 178.595 38.340 179.055 ;
        RECT 37.215 178.205 38.340 178.425 ;
        RECT 36.625 177.475 37.720 178.035 ;
        RECT 37.890 177.745 38.340 178.205 ;
        RECT 38.510 177.915 38.895 178.885 ;
        RECT 39.065 178.500 39.670 179.055 ;
        RECT 39.845 178.545 40.325 178.885 ;
        RECT 40.495 178.510 40.750 179.055 ;
        RECT 39.065 178.400 39.680 178.500 ;
        RECT 39.495 178.375 39.680 178.400 ;
        RECT 35.500 176.675 35.785 177.135 ;
        RECT 35.955 176.505 36.225 176.965 ;
        RECT 36.625 176.675 37.025 177.475 ;
        RECT 37.890 177.415 38.445 177.745 ;
        RECT 37.890 177.305 38.340 177.415 ;
        RECT 37.215 177.135 38.340 177.305 ;
        RECT 38.615 177.245 38.895 177.915 ;
        RECT 39.065 177.780 39.325 178.230 ;
        RECT 39.495 178.130 39.825 178.375 ;
        RECT 39.995 178.055 40.750 178.305 ;
        RECT 40.920 178.185 41.195 178.885 ;
        RECT 42.025 178.385 42.305 179.055 ;
        RECT 39.980 178.020 40.750 178.055 ;
        RECT 39.965 178.010 40.750 178.020 ;
        RECT 39.960 177.995 40.855 178.010 ;
        RECT 39.940 177.980 40.855 177.995 ;
        RECT 39.920 177.970 40.855 177.980 ;
        RECT 39.895 177.960 40.855 177.970 ;
        RECT 39.825 177.930 40.855 177.960 ;
        RECT 39.805 177.900 40.855 177.930 ;
        RECT 39.785 177.870 40.855 177.900 ;
        RECT 39.755 177.845 40.855 177.870 ;
        RECT 39.720 177.810 40.855 177.845 ;
        RECT 39.690 177.805 40.855 177.810 ;
        RECT 39.690 177.800 40.080 177.805 ;
        RECT 39.690 177.790 40.055 177.800 ;
        RECT 39.690 177.785 40.040 177.790 ;
        RECT 39.690 177.780 40.025 177.785 ;
        RECT 39.065 177.775 40.025 177.780 ;
        RECT 39.065 177.765 40.015 177.775 ;
        RECT 39.065 177.760 40.005 177.765 ;
        RECT 39.065 177.750 39.995 177.760 ;
        RECT 39.065 177.740 39.990 177.750 ;
        RECT 39.065 177.735 39.985 177.740 ;
        RECT 39.065 177.720 39.975 177.735 ;
        RECT 39.065 177.705 39.970 177.720 ;
        RECT 39.065 177.680 39.960 177.705 ;
        RECT 39.065 177.610 39.955 177.680 ;
        RECT 37.215 176.675 37.495 177.135 ;
        RECT 38.015 176.505 38.340 176.965 ;
        RECT 38.510 176.675 38.895 177.245 ;
        RECT 39.065 177.055 39.615 177.440 ;
        RECT 39.785 176.885 39.955 177.610 ;
        RECT 39.065 176.715 39.955 176.885 ;
        RECT 40.125 177.210 40.455 177.635 ;
        RECT 40.625 177.410 40.855 177.805 ;
        RECT 40.125 176.725 40.345 177.210 ;
        RECT 41.025 177.155 41.195 178.185 ;
        RECT 42.475 178.165 42.775 178.715 ;
        RECT 42.975 178.335 43.305 179.055 ;
        RECT 43.495 178.335 43.955 178.885 ;
        RECT 41.840 177.745 42.105 178.105 ;
        RECT 42.475 177.995 43.415 178.165 ;
        RECT 43.245 177.745 43.415 177.995 ;
        RECT 41.840 177.495 42.515 177.745 ;
        RECT 42.735 177.495 43.075 177.745 ;
        RECT 43.245 177.415 43.535 177.745 ;
        RECT 43.245 177.325 43.415 177.415 ;
        RECT 40.515 176.505 40.765 177.045 ;
        RECT 40.935 176.675 41.195 177.155 ;
        RECT 42.025 177.135 43.415 177.325 ;
        RECT 42.025 176.775 42.355 177.135 ;
        RECT 43.705 176.965 43.955 178.335 ;
        RECT 44.215 178.125 44.385 178.885 ;
        RECT 44.600 178.295 44.930 179.055 ;
        RECT 44.215 177.955 44.930 178.125 ;
        RECT 45.100 177.980 45.355 178.885 ;
        RECT 44.125 177.405 44.480 177.775 ;
        RECT 44.760 177.745 44.930 177.955 ;
        RECT 44.760 177.415 45.015 177.745 ;
        RECT 44.760 177.225 44.930 177.415 ;
        RECT 45.185 177.250 45.355 177.980 ;
        RECT 45.530 177.905 45.790 179.055 ;
        RECT 46.885 177.980 47.155 178.885 ;
        RECT 47.325 178.295 47.655 179.055 ;
        RECT 47.835 178.125 48.005 178.885 ;
        RECT 42.975 176.505 43.225 176.965 ;
        RECT 43.395 176.675 43.955 176.965 ;
        RECT 44.215 177.055 44.930 177.225 ;
        RECT 44.215 176.675 44.385 177.055 ;
        RECT 44.600 176.505 44.930 176.885 ;
        RECT 45.100 176.675 45.355 177.250 ;
        RECT 45.530 176.505 45.790 177.345 ;
        RECT 46.885 177.180 47.055 177.980 ;
        RECT 47.340 177.955 48.005 178.125 ;
        RECT 49.190 178.335 49.525 178.845 ;
        RECT 47.340 177.810 47.510 177.955 ;
        RECT 47.225 177.480 47.510 177.810 ;
        RECT 47.340 177.225 47.510 177.480 ;
        RECT 47.745 177.405 48.075 177.775 ;
        RECT 46.885 176.675 47.145 177.180 ;
        RECT 47.340 177.055 48.005 177.225 ;
        RECT 47.325 176.505 47.655 176.885 ;
        RECT 47.835 176.675 48.005 177.055 ;
        RECT 49.190 176.980 49.445 178.335 ;
        RECT 49.775 178.255 50.105 179.055 ;
        RECT 50.350 178.465 50.635 178.885 ;
        RECT 50.890 178.635 51.220 179.055 ;
        RECT 51.445 178.715 52.605 178.885 ;
        RECT 51.445 178.465 51.775 178.715 ;
        RECT 50.350 178.295 51.775 178.465 ;
        RECT 52.005 178.085 52.175 178.545 ;
        RECT 52.435 178.215 52.605 178.715 ;
        RECT 52.900 178.265 53.435 178.885 ;
        RECT 49.805 177.915 52.175 178.085 ;
        RECT 49.805 177.745 49.975 177.915 ;
        RECT 52.425 177.745 52.630 178.035 ;
        RECT 49.670 177.415 49.975 177.745 ;
        RECT 50.170 177.695 50.420 177.745 ;
        RECT 50.165 177.525 50.420 177.695 ;
        RECT 50.170 177.415 50.420 177.525 ;
        RECT 49.805 177.245 49.975 177.415 ;
        RECT 50.630 177.355 50.900 177.745 ;
        RECT 51.090 177.695 51.380 177.745 ;
        RECT 51.085 177.525 51.380 177.695 ;
        RECT 49.805 177.075 50.365 177.245 ;
        RECT 50.625 177.185 50.900 177.355 ;
        RECT 50.630 177.085 50.900 177.185 ;
        RECT 51.090 177.085 51.380 177.525 ;
        RECT 51.550 177.080 51.970 177.745 ;
        RECT 52.280 177.695 52.630 177.745 ;
        RECT 52.280 177.525 52.635 177.695 ;
        RECT 52.280 177.415 52.630 177.525 ;
        RECT 52.900 177.245 53.215 178.265 ;
        RECT 53.605 178.255 53.935 179.055 ;
        RECT 54.420 178.085 54.810 178.260 ;
        RECT 53.385 177.915 54.810 178.085 ;
        RECT 55.165 177.915 55.425 179.055 ;
        RECT 53.385 177.415 53.555 177.915 ;
        RECT 49.190 176.720 49.525 176.980 ;
        RECT 50.195 176.905 50.365 177.075 ;
        RECT 49.695 176.505 50.025 176.905 ;
        RECT 50.195 176.735 51.810 176.905 ;
        RECT 52.355 176.505 52.685 177.225 ;
        RECT 52.900 176.675 53.515 177.245 ;
        RECT 53.805 177.185 54.070 177.745 ;
        RECT 54.240 177.015 54.410 177.915 ;
        RECT 55.595 177.905 55.925 178.885 ;
        RECT 56.095 177.915 56.375 179.055 ;
        RECT 55.685 177.865 55.860 177.905 ;
        RECT 57.005 177.890 57.295 179.055 ;
        RECT 57.465 178.500 58.070 179.055 ;
        RECT 58.245 178.545 58.725 178.885 ;
        RECT 58.895 178.510 59.150 179.055 ;
        RECT 57.465 178.400 58.080 178.500 ;
        RECT 57.895 178.375 58.080 178.400 ;
        RECT 54.580 177.185 54.935 177.745 ;
        RECT 55.185 177.495 55.520 177.745 ;
        RECT 55.690 177.305 55.860 177.865 ;
        RECT 57.465 177.780 57.725 178.230 ;
        RECT 57.895 178.130 58.225 178.375 ;
        RECT 58.395 178.055 59.150 178.305 ;
        RECT 59.320 178.185 59.595 178.885 ;
        RECT 59.765 178.500 60.370 179.055 ;
        RECT 60.545 178.545 61.025 178.885 ;
        RECT 61.195 178.510 61.450 179.055 ;
        RECT 59.765 178.400 60.380 178.500 ;
        RECT 60.195 178.375 60.380 178.400 ;
        RECT 58.380 178.020 59.150 178.055 ;
        RECT 58.365 178.010 59.150 178.020 ;
        RECT 58.360 177.995 59.255 178.010 ;
        RECT 58.340 177.980 59.255 177.995 ;
        RECT 58.320 177.970 59.255 177.980 ;
        RECT 58.295 177.960 59.255 177.970 ;
        RECT 58.225 177.930 59.255 177.960 ;
        RECT 58.205 177.900 59.255 177.930 ;
        RECT 58.185 177.870 59.255 177.900 ;
        RECT 58.155 177.845 59.255 177.870 ;
        RECT 58.120 177.810 59.255 177.845 ;
        RECT 58.090 177.805 59.255 177.810 ;
        RECT 58.090 177.800 58.480 177.805 ;
        RECT 58.090 177.790 58.455 177.800 ;
        RECT 58.090 177.785 58.440 177.790 ;
        RECT 58.090 177.780 58.425 177.785 ;
        RECT 57.465 177.775 58.425 177.780 ;
        RECT 57.465 177.765 58.415 177.775 ;
        RECT 57.465 177.760 58.405 177.765 ;
        RECT 57.465 177.750 58.395 177.760 ;
        RECT 56.030 177.475 56.365 177.745 ;
        RECT 57.465 177.740 58.390 177.750 ;
        RECT 57.465 177.735 58.385 177.740 ;
        RECT 57.465 177.720 58.375 177.735 ;
        RECT 57.465 177.705 58.370 177.720 ;
        RECT 57.465 177.680 58.360 177.705 ;
        RECT 57.465 177.610 58.355 177.680 ;
        RECT 53.685 176.505 53.900 177.015 ;
        RECT 54.130 176.685 54.410 177.015 ;
        RECT 54.590 176.505 54.830 177.015 ;
        RECT 55.165 176.675 55.860 177.305 ;
        RECT 56.065 176.505 56.375 177.305 ;
        RECT 57.005 176.505 57.295 177.230 ;
        RECT 57.465 177.055 58.015 177.440 ;
        RECT 58.185 176.885 58.355 177.610 ;
        RECT 57.465 176.715 58.355 176.885 ;
        RECT 58.525 177.210 58.855 177.635 ;
        RECT 59.025 177.410 59.255 177.805 ;
        RECT 58.525 176.725 58.745 177.210 ;
        RECT 59.425 177.155 59.595 178.185 ;
        RECT 59.765 177.780 60.025 178.230 ;
        RECT 60.195 178.130 60.525 178.375 ;
        RECT 60.695 178.055 61.450 178.305 ;
        RECT 61.620 178.185 61.895 178.885 ;
        RECT 60.680 178.020 61.450 178.055 ;
        RECT 60.665 178.010 61.450 178.020 ;
        RECT 60.660 177.995 61.555 178.010 ;
        RECT 60.640 177.980 61.555 177.995 ;
        RECT 60.620 177.970 61.555 177.980 ;
        RECT 60.595 177.960 61.555 177.970 ;
        RECT 60.525 177.930 61.555 177.960 ;
        RECT 60.505 177.900 61.555 177.930 ;
        RECT 60.485 177.870 61.555 177.900 ;
        RECT 60.455 177.845 61.555 177.870 ;
        RECT 60.420 177.810 61.555 177.845 ;
        RECT 60.390 177.805 61.555 177.810 ;
        RECT 60.390 177.800 60.780 177.805 ;
        RECT 60.390 177.790 60.755 177.800 ;
        RECT 60.390 177.785 60.740 177.790 ;
        RECT 60.390 177.780 60.725 177.785 ;
        RECT 59.765 177.775 60.725 177.780 ;
        RECT 59.765 177.765 60.715 177.775 ;
        RECT 59.765 177.760 60.705 177.765 ;
        RECT 59.765 177.750 60.695 177.760 ;
        RECT 59.765 177.740 60.690 177.750 ;
        RECT 59.765 177.735 60.685 177.740 ;
        RECT 59.765 177.720 60.675 177.735 ;
        RECT 59.765 177.705 60.670 177.720 ;
        RECT 59.765 177.680 60.660 177.705 ;
        RECT 59.765 177.610 60.655 177.680 ;
        RECT 58.915 176.505 59.165 177.045 ;
        RECT 59.335 176.675 59.595 177.155 ;
        RECT 59.765 177.055 60.315 177.440 ;
        RECT 60.485 176.885 60.655 177.610 ;
        RECT 59.765 176.715 60.655 176.885 ;
        RECT 60.825 177.210 61.155 177.635 ;
        RECT 61.325 177.410 61.555 177.805 ;
        RECT 60.825 176.725 61.045 177.210 ;
        RECT 61.725 177.155 61.895 178.185 ;
        RECT 61.215 176.505 61.465 177.045 ;
        RECT 61.635 176.675 61.895 177.155 ;
        RECT 62.065 178.085 62.375 178.885 ;
        RECT 62.545 178.255 62.855 179.055 ;
        RECT 63.025 178.425 63.285 178.885 ;
        RECT 63.455 178.595 63.710 179.055 ;
        RECT 63.885 178.425 64.145 178.885 ;
        RECT 63.025 178.255 64.145 178.425 ;
        RECT 62.065 177.915 63.095 178.085 ;
        RECT 62.065 177.005 62.235 177.915 ;
        RECT 62.405 177.175 62.755 177.745 ;
        RECT 62.925 177.665 63.095 177.915 ;
        RECT 63.885 178.005 64.145 178.255 ;
        RECT 64.315 178.185 64.600 179.055 ;
        RECT 63.885 177.835 64.640 178.005 ;
        RECT 64.825 177.965 68.335 179.055 ;
        RECT 62.925 177.495 64.065 177.665 ;
        RECT 64.235 177.325 64.640 177.835 ;
        RECT 62.990 177.155 64.640 177.325 ;
        RECT 64.825 177.275 66.475 177.795 ;
        RECT 66.645 177.445 68.335 177.965 ;
        RECT 69.485 177.915 69.695 179.055 ;
        RECT 69.865 177.905 70.195 178.885 ;
        RECT 70.365 177.915 70.595 179.055 ;
        RECT 70.895 178.385 71.065 178.885 ;
        RECT 71.235 178.555 71.565 179.055 ;
        RECT 70.895 178.215 71.560 178.385 ;
        RECT 62.065 176.675 62.365 177.005 ;
        RECT 62.535 176.505 62.810 176.985 ;
        RECT 62.990 176.765 63.285 177.155 ;
        RECT 63.455 176.505 63.710 176.985 ;
        RECT 63.885 176.765 64.145 177.155 ;
        RECT 64.315 176.505 64.595 176.985 ;
        RECT 64.825 176.505 68.335 177.275 ;
        RECT 69.485 176.505 69.695 177.325 ;
        RECT 69.865 177.305 70.115 177.905 ;
        RECT 70.285 177.495 70.615 177.745 ;
        RECT 70.810 177.395 71.160 178.045 ;
        RECT 69.865 176.675 70.195 177.305 ;
        RECT 70.365 176.505 70.595 177.325 ;
        RECT 71.330 177.225 71.560 178.215 ;
        RECT 70.895 177.055 71.560 177.225 ;
        RECT 70.895 176.765 71.065 177.055 ;
        RECT 71.235 176.505 71.565 176.885 ;
        RECT 71.735 176.765 71.920 178.885 ;
        RECT 72.160 178.595 72.425 179.055 ;
        RECT 72.595 178.460 72.845 178.885 ;
        RECT 73.055 178.610 74.160 178.780 ;
        RECT 72.540 178.330 72.845 178.460 ;
        RECT 72.090 177.135 72.370 178.085 ;
        RECT 72.540 177.225 72.710 178.330 ;
        RECT 72.880 177.545 73.120 178.140 ;
        RECT 73.290 178.075 73.820 178.440 ;
        RECT 73.290 177.375 73.460 178.075 ;
        RECT 73.990 177.995 74.160 178.610 ;
        RECT 74.330 178.255 74.500 179.055 ;
        RECT 74.670 178.555 74.920 178.885 ;
        RECT 75.145 178.585 76.030 178.755 ;
        RECT 73.990 177.905 74.500 177.995 ;
        RECT 72.540 177.095 72.765 177.225 ;
        RECT 72.935 177.155 73.460 177.375 ;
        RECT 73.630 177.735 74.500 177.905 ;
        RECT 72.175 176.505 72.425 176.965 ;
        RECT 72.595 176.955 72.765 177.095 ;
        RECT 73.630 176.955 73.800 177.735 ;
        RECT 74.330 177.665 74.500 177.735 ;
        RECT 74.010 177.485 74.210 177.515 ;
        RECT 74.670 177.485 74.840 178.555 ;
        RECT 75.010 177.665 75.200 178.385 ;
        RECT 74.010 177.185 74.840 177.485 ;
        RECT 75.370 177.455 75.690 178.415 ;
        RECT 72.595 176.785 72.930 176.955 ;
        RECT 73.125 176.785 73.800 176.955 ;
        RECT 74.120 176.505 74.490 177.005 ;
        RECT 74.670 176.955 74.840 177.185 ;
        RECT 75.225 177.125 75.690 177.455 ;
        RECT 75.860 177.745 76.030 178.585 ;
        RECT 76.210 178.555 76.525 179.055 ;
        RECT 76.755 178.325 77.095 178.885 ;
        RECT 76.200 177.950 77.095 178.325 ;
        RECT 77.265 178.045 77.435 179.055 ;
        RECT 76.905 177.745 77.095 177.950 ;
        RECT 77.605 177.995 77.935 178.840 ;
        RECT 77.605 177.915 77.995 177.995 ;
        RECT 77.780 177.865 77.995 177.915 ;
        RECT 75.860 177.415 76.735 177.745 ;
        RECT 76.905 177.415 77.655 177.745 ;
        RECT 75.860 176.955 76.030 177.415 ;
        RECT 76.905 177.245 77.105 177.415 ;
        RECT 77.825 177.285 77.995 177.865 ;
        RECT 77.770 177.245 77.995 177.285 ;
        RECT 74.670 176.785 75.075 176.955 ;
        RECT 75.245 176.785 76.030 176.955 ;
        RECT 76.305 176.505 76.515 177.035 ;
        RECT 76.775 176.720 77.105 177.245 ;
        RECT 77.615 177.160 77.995 177.245 ;
        RECT 78.165 177.915 78.550 178.885 ;
        RECT 78.720 178.595 79.045 179.055 ;
        RECT 79.565 178.425 79.845 178.885 ;
        RECT 78.720 178.205 79.845 178.425 ;
        RECT 78.165 177.245 78.445 177.915 ;
        RECT 78.720 177.745 79.170 178.205 ;
        RECT 80.035 178.035 80.435 178.885 ;
        RECT 80.835 178.595 81.105 179.055 ;
        RECT 81.275 178.425 81.560 178.885 ;
        RECT 78.615 177.415 79.170 177.745 ;
        RECT 79.340 177.475 80.435 178.035 ;
        RECT 78.720 177.305 79.170 177.415 ;
        RECT 77.275 176.505 77.445 177.115 ;
        RECT 77.615 176.725 77.945 177.160 ;
        RECT 78.165 176.675 78.550 177.245 ;
        RECT 78.720 177.135 79.845 177.305 ;
        RECT 78.720 176.505 79.045 176.965 ;
        RECT 79.565 176.675 79.845 177.135 ;
        RECT 80.035 176.675 80.435 177.475 ;
        RECT 80.605 178.205 81.560 178.425 ;
        RECT 80.605 177.305 80.815 178.205 ;
        RECT 80.985 177.475 81.675 178.035 ;
        RECT 82.765 177.890 83.055 179.055 ;
        RECT 83.230 177.915 83.565 178.885 ;
        RECT 83.735 177.915 83.905 179.055 ;
        RECT 84.075 178.715 86.105 178.885 ;
        RECT 80.605 177.135 81.560 177.305 ;
        RECT 83.230 177.245 83.400 177.915 ;
        RECT 84.075 177.745 84.245 178.715 ;
        RECT 83.570 177.415 83.825 177.745 ;
        RECT 84.050 177.415 84.245 177.745 ;
        RECT 84.415 178.375 85.540 178.545 ;
        RECT 83.655 177.245 83.825 177.415 ;
        RECT 84.415 177.245 84.585 178.375 ;
        RECT 80.835 176.505 81.105 176.965 ;
        RECT 81.275 176.675 81.560 177.135 ;
        RECT 82.765 176.505 83.055 177.230 ;
        RECT 83.230 176.675 83.485 177.245 ;
        RECT 83.655 177.075 84.585 177.245 ;
        RECT 84.755 178.035 85.765 178.205 ;
        RECT 84.755 177.235 84.925 178.035 ;
        RECT 85.130 177.355 85.405 177.835 ;
        RECT 85.125 177.185 85.405 177.355 ;
        RECT 84.410 177.040 84.585 177.075 ;
        RECT 83.655 176.505 83.985 176.905 ;
        RECT 84.410 176.675 84.940 177.040 ;
        RECT 85.130 176.675 85.405 177.185 ;
        RECT 85.575 176.675 85.765 178.035 ;
        RECT 85.935 178.050 86.105 178.715 ;
        RECT 86.275 178.295 86.445 179.055 ;
        RECT 86.680 178.295 87.195 178.705 ;
        RECT 85.935 177.860 86.685 178.050 ;
        RECT 86.855 177.485 87.195 178.295 ;
        RECT 87.365 177.915 87.645 179.055 ;
        RECT 87.815 177.905 88.145 178.885 ;
        RECT 88.315 177.915 88.575 179.055 ;
        RECT 88.745 177.965 90.415 179.055 ;
        RECT 85.965 177.315 87.195 177.485 ;
        RECT 87.375 177.475 87.710 177.745 ;
        RECT 85.945 176.505 86.455 177.040 ;
        RECT 86.675 176.710 86.920 177.315 ;
        RECT 87.880 177.305 88.050 177.905 ;
        RECT 88.220 177.495 88.555 177.745 ;
        RECT 87.365 176.505 87.675 177.305 ;
        RECT 87.880 176.675 88.575 177.305 ;
        RECT 88.745 177.275 89.495 177.795 ;
        RECT 89.665 177.445 90.415 177.965 ;
        RECT 91.045 177.965 92.255 179.055 ;
        RECT 91.045 177.425 91.565 177.965 ;
        RECT 88.745 176.505 90.415 177.275 ;
        RECT 91.735 177.255 92.255 177.795 ;
        RECT 91.045 176.505 92.255 177.255 ;
        RECT 18.280 176.335 92.340 176.505 ;
        RECT 18.365 175.585 19.575 176.335 ;
        RECT 19.745 175.790 25.090 176.335 ;
        RECT 18.365 175.045 18.885 175.585 ;
        RECT 19.055 174.875 19.575 175.415 ;
        RECT 21.330 174.960 21.670 175.790 ;
        RECT 25.265 175.595 25.650 176.165 ;
        RECT 25.820 175.875 26.145 176.335 ;
        RECT 26.665 175.705 26.945 176.165 ;
        RECT 18.365 173.785 19.575 174.875 ;
        RECT 23.150 174.220 23.500 175.470 ;
        RECT 25.265 174.925 25.545 175.595 ;
        RECT 25.820 175.535 26.945 175.705 ;
        RECT 25.820 175.425 26.270 175.535 ;
        RECT 25.715 175.095 26.270 175.425 ;
        RECT 27.135 175.365 27.535 176.165 ;
        RECT 27.935 175.875 28.205 176.335 ;
        RECT 28.375 175.705 28.660 176.165 ;
        RECT 19.745 173.785 25.090 174.220 ;
        RECT 25.265 173.955 25.650 174.925 ;
        RECT 25.820 174.635 26.270 175.095 ;
        RECT 26.440 174.805 27.535 175.365 ;
        RECT 25.820 174.415 26.945 174.635 ;
        RECT 25.820 173.785 26.145 174.245 ;
        RECT 26.665 173.955 26.945 174.415 ;
        RECT 27.135 173.955 27.535 174.805 ;
        RECT 27.705 175.535 28.660 175.705 ;
        RECT 28.945 175.565 31.535 176.335 ;
        RECT 27.705 174.635 27.915 175.535 ;
        RECT 28.085 174.805 28.775 175.365 ;
        RECT 28.945 175.045 30.155 175.565 ;
        RECT 31.725 175.525 31.965 176.335 ;
        RECT 32.135 175.525 32.465 176.165 ;
        RECT 32.635 175.525 32.905 176.335 ;
        RECT 33.085 175.565 34.755 176.335 ;
        RECT 30.325 174.875 31.535 175.395 ;
        RECT 31.705 175.095 32.055 175.345 ;
        RECT 32.225 174.925 32.395 175.525 ;
        RECT 32.565 175.095 32.915 175.345 ;
        RECT 33.085 175.045 33.835 175.565 ;
        RECT 34.935 175.525 35.205 176.335 ;
        RECT 35.375 175.525 35.705 176.165 ;
        RECT 35.875 175.525 36.115 176.335 ;
        RECT 36.305 175.565 38.895 176.335 ;
        RECT 27.705 174.415 28.660 174.635 ;
        RECT 27.935 173.785 28.205 174.245 ;
        RECT 28.375 173.955 28.660 174.415 ;
        RECT 28.945 173.785 31.535 174.875 ;
        RECT 31.715 174.755 32.395 174.925 ;
        RECT 31.715 173.970 32.045 174.755 ;
        RECT 32.575 173.785 32.905 174.925 ;
        RECT 34.005 174.875 34.755 175.395 ;
        RECT 34.925 175.095 35.275 175.345 ;
        RECT 35.445 174.925 35.615 175.525 ;
        RECT 35.785 175.095 36.135 175.345 ;
        RECT 36.305 175.045 37.515 175.565 ;
        RECT 39.565 175.515 39.795 176.335 ;
        RECT 39.965 175.535 40.295 176.165 ;
        RECT 33.085 173.785 34.755 174.875 ;
        RECT 34.935 173.785 35.265 174.925 ;
        RECT 35.445 174.755 36.125 174.925 ;
        RECT 37.685 174.875 38.895 175.395 ;
        RECT 39.545 175.095 39.875 175.345 ;
        RECT 40.045 174.935 40.295 175.535 ;
        RECT 40.465 175.515 40.675 176.335 ;
        RECT 40.905 175.565 43.495 176.335 ;
        RECT 44.125 175.610 44.415 176.335 ;
        RECT 44.675 175.785 44.845 176.075 ;
        RECT 45.015 175.955 45.345 176.335 ;
        RECT 44.675 175.615 45.340 175.785 ;
        RECT 40.905 175.045 42.115 175.565 ;
        RECT 35.795 173.970 36.125 174.755 ;
        RECT 36.305 173.785 38.895 174.875 ;
        RECT 39.565 173.785 39.795 174.925 ;
        RECT 39.965 173.955 40.295 174.935 ;
        RECT 40.465 173.785 40.675 174.925 ;
        RECT 42.285 174.875 43.495 175.395 ;
        RECT 40.905 173.785 43.495 174.875 ;
        RECT 44.125 173.785 44.415 174.950 ;
        RECT 44.590 174.795 44.940 175.445 ;
        RECT 45.110 174.625 45.340 175.615 ;
        RECT 44.675 174.455 45.340 174.625 ;
        RECT 44.675 173.955 44.845 174.455 ;
        RECT 45.015 173.785 45.345 174.285 ;
        RECT 45.515 173.955 45.700 176.075 ;
        RECT 45.955 175.875 46.205 176.335 ;
        RECT 46.375 175.885 46.710 176.055 ;
        RECT 46.905 175.885 47.580 176.055 ;
        RECT 46.375 175.745 46.545 175.885 ;
        RECT 45.870 174.755 46.150 175.705 ;
        RECT 46.320 175.615 46.545 175.745 ;
        RECT 46.320 174.510 46.490 175.615 ;
        RECT 46.715 175.465 47.240 175.685 ;
        RECT 46.660 174.700 46.900 175.295 ;
        RECT 47.070 174.765 47.240 175.465 ;
        RECT 47.410 175.105 47.580 175.885 ;
        RECT 47.900 175.835 48.270 176.335 ;
        RECT 48.450 175.885 48.855 176.055 ;
        RECT 49.025 175.885 49.810 176.055 ;
        RECT 48.450 175.655 48.620 175.885 ;
        RECT 47.790 175.355 48.620 175.655 ;
        RECT 49.005 175.385 49.470 175.715 ;
        RECT 47.790 175.325 47.990 175.355 ;
        RECT 48.110 175.105 48.280 175.175 ;
        RECT 47.410 174.935 48.280 175.105 ;
        RECT 47.770 174.845 48.280 174.935 ;
        RECT 46.320 174.380 46.625 174.510 ;
        RECT 47.070 174.400 47.600 174.765 ;
        RECT 45.940 173.785 46.205 174.245 ;
        RECT 46.375 173.955 46.625 174.380 ;
        RECT 47.770 174.230 47.940 174.845 ;
        RECT 46.835 174.060 47.940 174.230 ;
        RECT 48.110 173.785 48.280 174.585 ;
        RECT 48.450 174.285 48.620 175.355 ;
        RECT 48.790 174.455 48.980 175.175 ;
        RECT 49.150 174.425 49.470 175.385 ;
        RECT 49.640 175.425 49.810 175.885 ;
        RECT 50.085 175.805 50.295 176.335 ;
        RECT 50.555 175.595 50.885 176.120 ;
        RECT 51.055 175.725 51.225 176.335 ;
        RECT 51.395 175.680 51.725 176.115 ;
        RECT 51.945 175.825 52.250 176.335 ;
        RECT 51.395 175.595 51.775 175.680 ;
        RECT 50.685 175.425 50.885 175.595 ;
        RECT 51.550 175.555 51.775 175.595 ;
        RECT 49.640 175.095 50.515 175.425 ;
        RECT 50.685 175.095 51.435 175.425 ;
        RECT 48.450 173.955 48.700 174.285 ;
        RECT 49.640 174.255 49.810 175.095 ;
        RECT 50.685 174.890 50.875 175.095 ;
        RECT 51.605 174.975 51.775 175.555 ;
        RECT 51.945 175.095 52.260 175.655 ;
        RECT 52.430 175.345 52.680 176.155 ;
        RECT 52.850 175.810 53.110 176.335 ;
        RECT 53.290 175.345 53.540 176.155 ;
        RECT 53.710 175.775 53.970 176.335 ;
        RECT 54.140 175.685 54.400 176.140 ;
        RECT 54.570 175.855 54.830 176.335 ;
        RECT 55.000 175.685 55.260 176.140 ;
        RECT 55.430 175.855 55.690 176.335 ;
        RECT 55.860 175.685 56.120 176.140 ;
        RECT 56.290 175.855 56.535 176.335 ;
        RECT 56.705 175.685 56.980 176.140 ;
        RECT 57.150 175.855 57.395 176.335 ;
        RECT 57.565 175.685 57.825 176.140 ;
        RECT 58.005 175.855 58.255 176.335 ;
        RECT 58.425 175.685 58.685 176.140 ;
        RECT 58.865 175.855 59.115 176.335 ;
        RECT 59.285 175.685 59.545 176.140 ;
        RECT 59.725 175.855 59.985 176.335 ;
        RECT 60.155 175.685 60.415 176.140 ;
        RECT 60.585 175.855 60.885 176.335 ;
        RECT 54.140 175.515 60.885 175.685 ;
        RECT 61.165 175.605 61.455 176.335 ;
        RECT 52.430 175.095 59.550 175.345 ;
        RECT 51.560 174.925 51.775 174.975 ;
        RECT 49.980 174.515 50.875 174.890 ;
        RECT 51.385 174.845 51.775 174.925 ;
        RECT 48.925 174.085 49.810 174.255 ;
        RECT 49.990 173.785 50.305 174.285 ;
        RECT 50.535 173.955 50.875 174.515 ;
        RECT 51.045 173.785 51.215 174.795 ;
        RECT 51.385 174.000 51.715 174.845 ;
        RECT 51.955 173.785 52.250 174.595 ;
        RECT 52.430 173.955 52.675 175.095 ;
        RECT 52.850 173.785 53.110 174.595 ;
        RECT 53.290 173.960 53.540 175.095 ;
        RECT 59.720 174.925 60.885 175.515 ;
        RECT 61.155 175.095 61.455 175.425 ;
        RECT 61.635 175.405 61.865 176.045 ;
        RECT 62.045 175.785 62.355 176.155 ;
        RECT 62.535 175.965 63.205 176.335 ;
        RECT 62.045 175.585 63.275 175.785 ;
        RECT 61.635 175.095 62.160 175.405 ;
        RECT 62.340 175.095 62.805 175.405 ;
        RECT 54.140 174.700 60.885 174.925 ;
        RECT 62.985 174.915 63.275 175.585 ;
        RECT 54.140 174.685 59.545 174.700 ;
        RECT 53.710 173.790 53.970 174.585 ;
        RECT 54.140 173.960 54.400 174.685 ;
        RECT 54.570 173.790 54.830 174.515 ;
        RECT 55.000 173.960 55.260 174.685 ;
        RECT 55.430 173.790 55.690 174.515 ;
        RECT 55.860 173.960 56.120 174.685 ;
        RECT 56.290 173.790 56.550 174.515 ;
        RECT 56.720 173.960 56.980 174.685 ;
        RECT 57.150 173.790 57.395 174.515 ;
        RECT 57.565 173.960 57.825 174.685 ;
        RECT 58.010 173.790 58.255 174.515 ;
        RECT 58.425 173.960 58.685 174.685 ;
        RECT 58.870 173.790 59.115 174.515 ;
        RECT 59.285 173.960 59.545 174.685 ;
        RECT 59.730 173.790 59.985 174.515 ;
        RECT 60.155 173.960 60.445 174.700 ;
        RECT 61.165 174.675 62.325 174.915 ;
        RECT 53.710 173.785 59.985 173.790 ;
        RECT 60.615 173.785 60.885 174.530 ;
        RECT 61.165 173.965 61.425 174.675 ;
        RECT 61.595 173.785 61.925 174.495 ;
        RECT 62.095 173.965 62.325 174.675 ;
        RECT 62.505 174.695 63.275 174.915 ;
        RECT 62.505 173.965 62.775 174.695 ;
        RECT 62.955 173.785 63.295 174.515 ;
        RECT 63.465 173.965 63.725 176.155 ;
        RECT 64.110 175.555 64.610 176.165 ;
        RECT 63.905 175.095 64.255 175.345 ;
        RECT 64.440 174.925 64.610 175.555 ;
        RECT 65.240 175.685 65.570 176.165 ;
        RECT 65.740 175.875 65.965 176.335 ;
        RECT 66.135 175.685 66.465 176.165 ;
        RECT 65.240 175.515 66.465 175.685 ;
        RECT 66.655 175.535 66.905 176.335 ;
        RECT 67.075 175.535 67.415 176.165 ;
        RECT 67.610 175.945 67.940 176.335 ;
        RECT 68.110 175.775 68.335 176.155 ;
        RECT 64.780 175.145 65.110 175.345 ;
        RECT 65.280 175.145 65.610 175.345 ;
        RECT 65.780 175.145 66.200 175.345 ;
        RECT 66.375 175.175 67.070 175.345 ;
        RECT 66.375 174.925 66.545 175.175 ;
        RECT 67.240 174.925 67.415 175.535 ;
        RECT 67.595 175.095 67.835 175.745 ;
        RECT 68.005 175.595 68.335 175.775 ;
        RECT 68.005 174.925 68.180 175.595 ;
        RECT 68.535 175.425 68.765 176.045 ;
        RECT 68.945 175.605 69.245 176.335 ;
        RECT 69.885 175.610 70.175 176.335 ;
        RECT 70.345 175.595 70.730 176.165 ;
        RECT 70.900 175.875 71.225 176.335 ;
        RECT 71.745 175.705 72.025 176.165 ;
        RECT 68.350 175.095 68.765 175.425 ;
        RECT 68.945 175.095 69.240 175.425 ;
        RECT 64.110 174.755 66.545 174.925 ;
        RECT 64.110 173.955 64.440 174.755 ;
        RECT 64.610 173.785 64.940 174.585 ;
        RECT 65.240 173.955 65.570 174.755 ;
        RECT 66.215 173.785 66.465 174.585 ;
        RECT 66.735 173.785 66.905 174.925 ;
        RECT 67.075 173.955 67.415 174.925 ;
        RECT 67.595 174.735 68.180 174.925 ;
        RECT 67.595 173.965 67.870 174.735 ;
        RECT 68.350 174.565 69.245 174.895 ;
        RECT 68.040 174.395 69.245 174.565 ;
        RECT 68.040 173.965 68.370 174.395 ;
        RECT 68.540 173.785 68.735 174.225 ;
        RECT 68.915 173.965 69.245 174.395 ;
        RECT 69.885 173.785 70.175 174.950 ;
        RECT 70.345 174.925 70.625 175.595 ;
        RECT 70.900 175.535 72.025 175.705 ;
        RECT 70.900 175.425 71.350 175.535 ;
        RECT 70.795 175.095 71.350 175.425 ;
        RECT 72.215 175.365 72.615 176.165 ;
        RECT 73.015 175.875 73.285 176.335 ;
        RECT 73.455 175.705 73.740 176.165 ;
        RECT 70.345 173.955 70.730 174.925 ;
        RECT 70.900 174.635 71.350 175.095 ;
        RECT 71.520 174.805 72.615 175.365 ;
        RECT 70.900 174.415 72.025 174.635 ;
        RECT 70.900 173.785 71.225 174.245 ;
        RECT 71.745 173.955 72.025 174.415 ;
        RECT 72.215 173.955 72.615 174.805 ;
        RECT 72.785 175.535 73.740 175.705 ;
        RECT 72.785 174.635 72.995 175.535 ;
        RECT 73.165 174.805 73.855 175.365 ;
        RECT 74.025 175.350 74.295 176.165 ;
        RECT 74.465 175.595 75.135 176.335 ;
        RECT 75.305 175.765 75.600 176.110 ;
        RECT 75.780 175.935 76.155 176.335 ;
        RECT 76.370 175.765 76.700 176.110 ;
        RECT 75.305 175.595 76.700 175.765 ;
        RECT 76.950 175.595 77.535 176.165 ;
        RECT 78.325 175.775 78.655 176.165 ;
        RECT 78.825 175.945 80.010 176.115 ;
        RECT 80.270 175.865 80.440 176.335 ;
        RECT 78.325 175.595 78.835 175.775 ;
        RECT 72.785 174.415 73.740 174.635 ;
        RECT 73.015 173.785 73.285 174.245 ;
        RECT 73.455 173.955 73.740 174.415 ;
        RECT 74.025 173.955 74.375 175.350 ;
        RECT 74.545 174.925 74.715 175.425 ;
        RECT 74.885 175.095 75.220 175.425 ;
        RECT 75.390 175.095 75.730 175.425 ;
        RECT 74.545 174.755 75.290 174.925 ;
        RECT 74.545 173.785 74.950 174.585 ;
        RECT 75.120 174.125 75.290 174.755 ;
        RECT 75.460 174.350 75.730 175.095 ;
        RECT 75.920 175.095 76.210 175.425 ;
        RECT 76.380 175.095 76.780 175.425 ;
        RECT 75.920 174.350 76.155 175.095 ;
        RECT 76.950 174.925 77.120 175.595 ;
        RECT 77.290 175.095 77.535 175.425 ;
        RECT 78.165 175.135 78.495 175.425 ;
        RECT 78.665 174.965 78.835 175.595 ;
        RECT 79.240 175.685 79.625 175.775 ;
        RECT 80.610 175.685 80.940 176.150 ;
        RECT 79.240 175.515 80.940 175.685 ;
        RECT 81.110 175.515 81.280 176.335 ;
        RECT 81.450 175.515 82.135 176.155 ;
        RECT 82.395 175.785 82.565 176.075 ;
        RECT 82.735 175.955 83.065 176.335 ;
        RECT 82.395 175.615 83.060 175.785 ;
        RECT 79.005 175.135 79.335 175.345 ;
        RECT 79.515 175.095 79.895 175.345 ;
        RECT 76.325 174.755 77.535 174.925 ;
        RECT 76.325 174.125 76.655 174.755 ;
        RECT 75.120 173.955 76.655 174.125 ;
        RECT 76.840 173.785 77.075 174.585 ;
        RECT 77.245 173.955 77.535 174.755 ;
        RECT 78.320 174.795 79.405 174.965 ;
        RECT 78.320 173.955 78.620 174.795 ;
        RECT 78.815 173.785 79.065 174.625 ;
        RECT 79.235 174.545 79.405 174.795 ;
        RECT 79.575 174.715 79.895 175.095 ;
        RECT 80.085 175.135 80.570 175.345 ;
        RECT 80.760 175.135 81.210 175.345 ;
        RECT 81.380 175.135 81.715 175.345 ;
        RECT 80.085 174.975 80.460 175.135 ;
        RECT 80.065 174.805 80.460 174.975 ;
        RECT 81.380 174.965 81.550 175.135 ;
        RECT 80.085 174.715 80.460 174.805 ;
        RECT 80.630 174.795 81.550 174.965 ;
        RECT 80.630 174.545 80.800 174.795 ;
        RECT 79.235 174.375 80.800 174.545 ;
        RECT 79.655 173.955 80.460 174.375 ;
        RECT 80.970 173.785 81.300 174.625 ;
        RECT 81.885 174.545 82.135 175.515 ;
        RECT 82.310 174.795 82.660 175.445 ;
        RECT 82.830 174.625 83.060 175.615 ;
        RECT 81.470 173.955 82.135 174.545 ;
        RECT 82.395 174.455 83.060 174.625 ;
        RECT 82.395 173.955 82.565 174.455 ;
        RECT 82.735 173.785 83.065 174.285 ;
        RECT 83.235 173.955 83.460 176.075 ;
        RECT 83.675 175.875 83.925 176.335 ;
        RECT 84.110 175.885 84.440 176.055 ;
        RECT 84.620 175.885 85.370 176.055 ;
        RECT 83.660 174.755 83.940 175.355 ;
        RECT 84.110 174.355 84.280 175.885 ;
        RECT 84.450 175.385 85.030 175.715 ;
        RECT 84.450 174.515 84.690 175.385 ;
        RECT 85.200 175.105 85.370 175.885 ;
        RECT 85.620 175.835 85.990 176.335 ;
        RECT 86.170 175.885 86.630 176.055 ;
        RECT 86.860 175.885 87.530 176.055 ;
        RECT 86.170 175.655 86.340 175.885 ;
        RECT 85.540 175.355 86.340 175.655 ;
        RECT 86.510 175.385 87.060 175.715 ;
        RECT 85.540 175.325 85.710 175.355 ;
        RECT 85.830 175.105 86.000 175.175 ;
        RECT 85.200 174.935 86.000 175.105 ;
        RECT 85.490 174.845 86.000 174.935 ;
        RECT 84.880 174.410 85.320 174.765 ;
        RECT 83.660 173.785 83.925 174.245 ;
        RECT 84.110 173.980 84.345 174.355 ;
        RECT 85.490 174.230 85.660 174.845 ;
        RECT 84.590 174.060 85.660 174.230 ;
        RECT 85.830 173.785 86.000 174.585 ;
        RECT 86.170 174.285 86.340 175.355 ;
        RECT 86.510 174.455 86.700 175.175 ;
        RECT 86.870 174.845 87.060 175.385 ;
        RECT 87.360 175.345 87.530 175.885 ;
        RECT 87.845 175.805 88.015 176.335 ;
        RECT 88.310 175.685 88.670 176.125 ;
        RECT 88.845 175.855 89.015 176.335 ;
        RECT 89.205 175.690 89.540 176.115 ;
        RECT 89.715 175.860 89.885 176.335 ;
        RECT 90.060 175.690 90.395 176.115 ;
        RECT 90.565 175.860 90.735 176.335 ;
        RECT 88.310 175.515 88.810 175.685 ;
        RECT 89.205 175.520 90.875 175.690 ;
        RECT 91.045 175.585 92.255 176.335 ;
        RECT 88.640 175.345 88.810 175.515 ;
        RECT 87.360 175.175 88.450 175.345 ;
        RECT 88.640 175.175 90.460 175.345 ;
        RECT 86.870 174.515 87.190 174.845 ;
        RECT 86.170 173.955 86.420 174.285 ;
        RECT 87.360 174.255 87.530 175.175 ;
        RECT 88.640 174.920 88.810 175.175 ;
        RECT 90.630 174.955 90.875 175.520 ;
        RECT 87.700 174.750 88.810 174.920 ;
        RECT 89.205 174.785 90.875 174.955 ;
        RECT 91.045 174.875 91.565 175.415 ;
        RECT 91.735 175.045 92.255 175.585 ;
        RECT 87.700 174.590 88.560 174.750 ;
        RECT 86.645 174.085 87.530 174.255 ;
        RECT 87.710 173.785 87.925 174.285 ;
        RECT 88.390 173.965 88.560 174.590 ;
        RECT 88.845 173.785 89.025 174.565 ;
        RECT 89.205 174.025 89.540 174.785 ;
        RECT 89.720 173.785 89.890 174.615 ;
        RECT 90.060 174.025 90.390 174.785 ;
        RECT 90.560 173.785 90.730 174.615 ;
        RECT 91.045 173.785 92.255 174.875 ;
        RECT 18.280 173.615 92.340 173.785 ;
        RECT 18.365 172.525 19.575 173.615 ;
        RECT 19.745 172.525 22.335 173.615 ;
        RECT 23.055 172.945 23.225 173.445 ;
        RECT 23.395 173.115 23.725 173.615 ;
        RECT 23.055 172.775 23.720 172.945 ;
        RECT 18.365 171.815 18.885 172.355 ;
        RECT 19.055 171.985 19.575 172.525 ;
        RECT 19.745 171.835 20.955 172.355 ;
        RECT 21.125 172.005 22.335 172.525 ;
        RECT 22.970 171.955 23.320 172.605 ;
        RECT 18.365 171.065 19.575 171.815 ;
        RECT 19.745 171.065 22.335 171.835 ;
        RECT 23.490 171.785 23.720 172.775 ;
        RECT 23.055 171.615 23.720 171.785 ;
        RECT 23.055 171.325 23.225 171.615 ;
        RECT 23.395 171.065 23.725 171.445 ;
        RECT 23.895 171.325 24.080 173.445 ;
        RECT 24.320 173.155 24.585 173.615 ;
        RECT 24.755 173.020 25.005 173.445 ;
        RECT 25.215 173.170 26.320 173.340 ;
        RECT 24.700 172.890 25.005 173.020 ;
        RECT 24.250 171.695 24.530 172.645 ;
        RECT 24.700 171.785 24.870 172.890 ;
        RECT 25.040 172.105 25.280 172.700 ;
        RECT 25.450 172.635 25.980 173.000 ;
        RECT 25.450 171.935 25.620 172.635 ;
        RECT 26.150 172.555 26.320 173.170 ;
        RECT 26.490 172.815 26.660 173.615 ;
        RECT 26.830 173.115 27.080 173.445 ;
        RECT 27.305 173.145 28.190 173.315 ;
        RECT 26.150 172.465 26.660 172.555 ;
        RECT 24.700 171.655 24.925 171.785 ;
        RECT 25.095 171.715 25.620 171.935 ;
        RECT 25.790 172.295 26.660 172.465 ;
        RECT 24.335 171.065 24.585 171.525 ;
        RECT 24.755 171.515 24.925 171.655 ;
        RECT 25.790 171.515 25.960 172.295 ;
        RECT 26.490 172.225 26.660 172.295 ;
        RECT 26.170 172.045 26.370 172.075 ;
        RECT 26.830 172.045 27.000 173.115 ;
        RECT 27.170 172.225 27.360 172.945 ;
        RECT 26.170 171.745 27.000 172.045 ;
        RECT 27.530 172.015 27.850 172.975 ;
        RECT 24.755 171.345 25.090 171.515 ;
        RECT 25.285 171.345 25.960 171.515 ;
        RECT 26.280 171.065 26.650 171.565 ;
        RECT 26.830 171.515 27.000 171.745 ;
        RECT 27.385 171.685 27.850 172.015 ;
        RECT 28.020 172.305 28.190 173.145 ;
        RECT 28.370 173.115 28.685 173.615 ;
        RECT 28.915 172.885 29.255 173.445 ;
        RECT 28.360 172.510 29.255 172.885 ;
        RECT 29.425 172.605 29.595 173.615 ;
        RECT 29.065 172.305 29.255 172.510 ;
        RECT 29.765 172.555 30.095 173.400 ;
        RECT 29.765 172.475 30.155 172.555 ;
        RECT 29.940 172.425 30.155 172.475 ;
        RECT 31.245 172.450 31.535 173.615 ;
        RECT 31.715 172.665 31.990 173.435 ;
        RECT 32.160 173.005 32.490 173.435 ;
        RECT 32.660 173.175 32.855 173.615 ;
        RECT 33.035 173.005 33.365 173.435 ;
        RECT 32.160 172.835 33.365 173.005 ;
        RECT 31.715 172.475 32.300 172.665 ;
        RECT 32.470 172.505 33.365 172.835 ;
        RECT 33.545 172.525 35.215 173.615 ;
        RECT 28.020 171.975 28.895 172.305 ;
        RECT 29.065 171.975 29.815 172.305 ;
        RECT 28.020 171.515 28.190 171.975 ;
        RECT 29.065 171.805 29.265 171.975 ;
        RECT 29.985 171.845 30.155 172.425 ;
        RECT 29.930 171.805 30.155 171.845 ;
        RECT 26.830 171.345 27.235 171.515 ;
        RECT 27.405 171.345 28.190 171.515 ;
        RECT 28.465 171.065 28.675 171.595 ;
        RECT 28.935 171.280 29.265 171.805 ;
        RECT 29.775 171.720 30.155 171.805 ;
        RECT 29.435 171.065 29.605 171.675 ;
        RECT 29.775 171.285 30.105 171.720 ;
        RECT 31.245 171.065 31.535 171.790 ;
        RECT 31.715 171.655 31.955 172.305 ;
        RECT 32.125 171.805 32.300 172.475 ;
        RECT 32.470 171.975 32.885 172.305 ;
        RECT 33.065 171.975 33.360 172.305 ;
        RECT 32.125 171.625 32.455 171.805 ;
        RECT 31.730 171.065 32.060 171.455 ;
        RECT 32.230 171.245 32.455 171.625 ;
        RECT 32.655 171.355 32.885 171.975 ;
        RECT 33.545 171.835 34.295 172.355 ;
        RECT 34.465 172.005 35.215 172.525 ;
        RECT 35.385 172.475 35.660 173.445 ;
        RECT 35.870 172.815 36.150 173.615 ;
        RECT 36.320 173.105 37.935 173.435 ;
        RECT 36.320 172.765 37.495 172.935 ;
        RECT 36.320 172.645 36.490 172.765 ;
        RECT 35.830 172.475 36.490 172.645 ;
        RECT 33.065 171.065 33.365 171.795 ;
        RECT 33.545 171.065 35.215 171.835 ;
        RECT 35.385 171.740 35.555 172.475 ;
        RECT 35.830 172.305 36.000 172.475 ;
        RECT 36.750 172.305 36.995 172.595 ;
        RECT 37.165 172.475 37.495 172.765 ;
        RECT 37.755 172.305 37.925 172.865 ;
        RECT 38.175 172.475 38.435 173.615 ;
        RECT 38.610 173.235 38.945 173.615 ;
        RECT 35.725 171.975 36.000 172.305 ;
        RECT 36.170 171.975 36.995 172.305 ;
        RECT 37.210 171.975 37.925 172.305 ;
        RECT 38.095 172.055 38.430 172.305 ;
        RECT 35.830 171.805 36.000 171.975 ;
        RECT 37.675 171.885 37.925 171.975 ;
        RECT 35.385 171.395 35.660 171.740 ;
        RECT 35.830 171.635 37.495 171.805 ;
        RECT 35.850 171.065 36.225 171.465 ;
        RECT 36.395 171.285 36.565 171.635 ;
        RECT 36.735 171.065 37.065 171.465 ;
        RECT 37.235 171.235 37.495 171.635 ;
        RECT 37.675 171.465 38.005 171.885 ;
        RECT 38.175 171.065 38.435 171.885 ;
        RECT 38.605 171.745 38.845 173.055 ;
        RECT 39.115 172.645 39.365 173.445 ;
        RECT 39.585 172.895 39.915 173.615 ;
        RECT 40.100 172.645 40.350 173.445 ;
        RECT 40.815 172.815 41.145 173.615 ;
        RECT 41.315 173.185 41.655 173.445 ;
        RECT 39.015 172.475 41.205 172.645 ;
        RECT 39.015 171.565 39.185 172.475 ;
        RECT 40.890 172.305 41.205 172.475 ;
        RECT 38.690 171.235 39.185 171.565 ;
        RECT 39.405 171.340 39.755 172.305 ;
        RECT 39.935 171.335 40.235 172.305 ;
        RECT 40.415 171.335 40.695 172.305 ;
        RECT 40.890 172.055 41.220 172.305 ;
        RECT 40.875 171.065 41.145 171.865 ;
        RECT 41.395 171.785 41.655 173.185 ;
        RECT 42.835 172.685 43.005 173.445 ;
        RECT 43.220 172.855 43.550 173.615 ;
        RECT 42.835 172.515 43.550 172.685 ;
        RECT 43.720 172.540 43.975 173.445 ;
        RECT 42.745 171.965 43.100 172.335 ;
        RECT 43.380 172.305 43.550 172.515 ;
        RECT 43.380 171.975 43.635 172.305 ;
        RECT 43.380 171.785 43.550 171.975 ;
        RECT 43.805 171.810 43.975 172.540 ;
        RECT 44.150 172.465 44.410 173.615 ;
        RECT 44.585 172.525 46.255 173.615 ;
        RECT 41.315 171.275 41.655 171.785 ;
        RECT 42.835 171.615 43.550 171.785 ;
        RECT 42.835 171.235 43.005 171.615 ;
        RECT 43.220 171.065 43.550 171.445 ;
        RECT 43.720 171.235 43.975 171.810 ;
        RECT 44.150 171.065 44.410 171.905 ;
        RECT 44.585 171.835 45.335 172.355 ;
        RECT 45.505 172.005 46.255 172.525 ;
        RECT 46.885 172.895 47.345 173.445 ;
        RECT 47.535 172.895 47.865 173.615 ;
        RECT 44.585 171.065 46.255 171.835 ;
        RECT 46.885 171.525 47.135 172.895 ;
        RECT 48.065 172.725 48.365 173.275 ;
        RECT 48.535 172.945 48.815 173.615 ;
        RECT 49.185 173.180 54.530 173.615 ;
        RECT 47.425 172.555 48.365 172.725 ;
        RECT 47.425 172.305 47.595 172.555 ;
        RECT 48.735 172.305 49.000 172.665 ;
        RECT 47.305 171.975 47.595 172.305 ;
        RECT 47.765 172.055 48.105 172.305 ;
        RECT 48.325 172.055 49.000 172.305 ;
        RECT 47.425 171.885 47.595 171.975 ;
        RECT 47.425 171.695 48.815 171.885 ;
        RECT 46.885 171.235 47.445 171.525 ;
        RECT 47.615 171.065 47.865 171.525 ;
        RECT 48.485 171.335 48.815 171.695 ;
        RECT 50.770 171.610 51.110 172.440 ;
        RECT 52.590 171.930 52.940 173.180 ;
        RECT 54.705 172.525 56.375 173.615 ;
        RECT 54.705 171.835 55.455 172.355 ;
        RECT 55.625 172.005 56.375 172.525 ;
        RECT 57.005 172.450 57.295 173.615 ;
        RECT 57.465 172.475 57.850 173.435 ;
        RECT 58.065 172.815 58.355 173.615 ;
        RECT 58.525 173.275 59.890 173.445 ;
        RECT 58.525 172.645 58.695 173.275 ;
        RECT 58.020 172.475 58.695 172.645 ;
        RECT 49.185 171.065 54.530 171.610 ;
        RECT 54.705 171.065 56.375 171.835 ;
        RECT 57.465 171.805 57.640 172.475 ;
        RECT 58.020 172.305 58.190 172.475 ;
        RECT 58.865 172.305 59.190 173.105 ;
        RECT 59.560 173.065 59.890 173.275 ;
        RECT 59.560 172.815 60.515 173.065 ;
        RECT 57.825 172.055 58.190 172.305 ;
        RECT 58.385 172.055 58.635 172.305 ;
        RECT 57.825 171.975 58.015 172.055 ;
        RECT 58.385 171.975 58.555 172.055 ;
        RECT 58.845 171.975 59.190 172.305 ;
        RECT 59.360 171.975 59.635 172.640 ;
        RECT 59.820 171.975 60.175 172.640 ;
        RECT 60.345 171.805 60.515 172.815 ;
        RECT 60.685 172.475 60.975 173.615 ;
        RECT 61.155 173.005 61.485 173.435 ;
        RECT 61.665 173.175 61.860 173.615 ;
        RECT 62.030 173.005 62.360 173.435 ;
        RECT 61.155 172.835 62.360 173.005 ;
        RECT 61.155 172.505 62.050 172.835 ;
        RECT 62.530 172.665 62.805 173.435 ;
        RECT 62.220 172.475 62.805 172.665 ;
        RECT 63.045 172.475 63.255 173.615 ;
        RECT 60.700 171.975 60.975 172.305 ;
        RECT 61.160 171.975 61.455 172.305 ;
        RECT 61.635 171.975 62.050 172.305 ;
        RECT 57.005 171.065 57.295 171.790 ;
        RECT 57.465 171.235 57.975 171.805 ;
        RECT 58.520 171.635 59.920 171.805 ;
        RECT 58.145 171.065 58.315 171.625 ;
        RECT 58.520 171.235 58.850 171.635 ;
        RECT 59.025 171.065 59.355 171.465 ;
        RECT 59.590 171.445 59.920 171.635 ;
        RECT 60.090 171.615 60.515 171.805 ;
        RECT 60.685 171.445 60.975 171.715 ;
        RECT 59.590 171.235 60.975 171.445 ;
        RECT 61.155 171.065 61.455 171.795 ;
        RECT 61.635 171.355 61.865 171.975 ;
        RECT 62.220 171.805 62.395 172.475 ;
        RECT 63.425 172.465 63.755 173.445 ;
        RECT 63.925 172.475 64.155 173.615 ;
        RECT 64.915 172.945 65.085 173.445 ;
        RECT 65.255 173.115 65.585 173.615 ;
        RECT 64.915 172.775 65.580 172.945 ;
        RECT 62.065 171.625 62.395 171.805 ;
        RECT 62.565 171.655 62.805 172.305 ;
        RECT 62.065 171.245 62.290 171.625 ;
        RECT 62.460 171.065 62.790 171.455 ;
        RECT 63.045 171.065 63.255 171.885 ;
        RECT 63.425 171.865 63.675 172.465 ;
        RECT 63.845 172.055 64.175 172.305 ;
        RECT 64.830 171.955 65.180 172.605 ;
        RECT 63.425 171.235 63.755 171.865 ;
        RECT 63.925 171.065 64.155 171.885 ;
        RECT 65.350 171.785 65.580 172.775 ;
        RECT 64.915 171.615 65.580 171.785 ;
        RECT 64.915 171.325 65.085 171.615 ;
        RECT 65.255 171.065 65.585 171.445 ;
        RECT 65.755 171.325 65.940 173.445 ;
        RECT 66.180 173.155 66.445 173.615 ;
        RECT 66.615 173.020 66.865 173.445 ;
        RECT 67.075 173.170 68.180 173.340 ;
        RECT 66.560 172.890 66.865 173.020 ;
        RECT 66.110 171.695 66.390 172.645 ;
        RECT 66.560 171.785 66.730 172.890 ;
        RECT 66.900 172.105 67.140 172.700 ;
        RECT 67.310 172.635 67.840 173.000 ;
        RECT 67.310 171.935 67.480 172.635 ;
        RECT 68.010 172.555 68.180 173.170 ;
        RECT 68.350 172.815 68.520 173.615 ;
        RECT 68.690 173.115 68.940 173.445 ;
        RECT 69.165 173.145 70.050 173.315 ;
        RECT 68.010 172.465 68.520 172.555 ;
        RECT 66.560 171.655 66.785 171.785 ;
        RECT 66.955 171.715 67.480 171.935 ;
        RECT 67.650 172.295 68.520 172.465 ;
        RECT 66.195 171.065 66.445 171.525 ;
        RECT 66.615 171.515 66.785 171.655 ;
        RECT 67.650 171.515 67.820 172.295 ;
        RECT 68.350 172.225 68.520 172.295 ;
        RECT 68.030 172.045 68.230 172.075 ;
        RECT 68.690 172.045 68.860 173.115 ;
        RECT 69.030 172.225 69.220 172.945 ;
        RECT 68.030 171.745 68.860 172.045 ;
        RECT 69.390 172.015 69.710 172.975 ;
        RECT 66.615 171.345 66.950 171.515 ;
        RECT 67.145 171.345 67.820 171.515 ;
        RECT 68.140 171.065 68.510 171.565 ;
        RECT 68.690 171.515 68.860 171.745 ;
        RECT 69.245 171.685 69.710 172.015 ;
        RECT 69.880 172.305 70.050 173.145 ;
        RECT 70.230 173.115 70.545 173.615 ;
        RECT 70.775 172.885 71.115 173.445 ;
        RECT 70.220 172.510 71.115 172.885 ;
        RECT 71.285 172.605 71.455 173.615 ;
        RECT 70.925 172.305 71.115 172.510 ;
        RECT 71.625 172.555 71.955 173.400 ;
        RECT 72.185 173.180 77.530 173.615 ;
        RECT 71.625 172.475 72.015 172.555 ;
        RECT 71.800 172.425 72.015 172.475 ;
        RECT 69.880 171.975 70.755 172.305 ;
        RECT 70.925 171.975 71.675 172.305 ;
        RECT 69.880 171.515 70.050 171.975 ;
        RECT 70.925 171.805 71.125 171.975 ;
        RECT 71.845 171.845 72.015 172.425 ;
        RECT 71.790 171.805 72.015 171.845 ;
        RECT 68.690 171.345 69.095 171.515 ;
        RECT 69.265 171.345 70.050 171.515 ;
        RECT 70.325 171.065 70.535 171.595 ;
        RECT 70.795 171.280 71.125 171.805 ;
        RECT 71.635 171.720 72.015 171.805 ;
        RECT 71.295 171.065 71.465 171.675 ;
        RECT 71.635 171.285 71.965 171.720 ;
        RECT 73.770 171.610 74.110 172.440 ;
        RECT 75.590 171.930 75.940 173.180 ;
        RECT 77.705 172.525 81.215 173.615 ;
        RECT 77.705 171.835 79.355 172.355 ;
        RECT 79.525 172.005 81.215 172.525 ;
        RECT 81.395 172.645 81.725 173.430 ;
        RECT 81.395 172.475 82.075 172.645 ;
        RECT 82.255 172.475 82.585 173.615 ;
        RECT 81.385 172.055 81.735 172.305 ;
        RECT 81.905 171.875 82.075 172.475 ;
        RECT 82.765 172.450 83.055 173.615 ;
        RECT 83.235 172.645 83.565 173.430 ;
        RECT 83.235 172.475 83.915 172.645 ;
        RECT 84.095 172.475 84.425 173.615 ;
        RECT 84.605 173.180 89.950 173.615 ;
        RECT 82.245 172.055 82.595 172.305 ;
        RECT 83.225 172.055 83.575 172.305 ;
        RECT 83.745 171.875 83.915 172.475 ;
        RECT 84.085 172.055 84.435 172.305 ;
        RECT 72.185 171.065 77.530 171.610 ;
        RECT 77.705 171.065 81.215 171.835 ;
        RECT 81.405 171.065 81.645 171.875 ;
        RECT 81.815 171.235 82.145 171.875 ;
        RECT 82.315 171.065 82.585 171.875 ;
        RECT 82.765 171.065 83.055 171.790 ;
        RECT 83.245 171.065 83.485 171.875 ;
        RECT 83.655 171.235 83.985 171.875 ;
        RECT 84.155 171.065 84.425 171.875 ;
        RECT 86.190 171.610 86.530 172.440 ;
        RECT 88.010 171.930 88.360 173.180 ;
        RECT 91.045 172.525 92.255 173.615 ;
        RECT 91.045 171.985 91.565 172.525 ;
        RECT 91.735 171.815 92.255 172.355 ;
        RECT 84.605 171.065 89.950 171.610 ;
        RECT 91.045 171.065 92.255 171.815 ;
        RECT 18.280 170.895 92.340 171.065 ;
        RECT 18.365 170.145 19.575 170.895 ;
        RECT 19.745 170.350 25.090 170.895 ;
        RECT 18.365 169.605 18.885 170.145 ;
        RECT 19.055 169.435 19.575 169.975 ;
        RECT 21.330 169.520 21.670 170.350 ;
        RECT 25.265 170.125 26.935 170.895 ;
        RECT 18.365 168.345 19.575 169.435 ;
        RECT 23.150 168.780 23.500 170.030 ;
        RECT 25.265 169.605 26.015 170.125 ;
        RECT 27.105 170.095 27.415 170.895 ;
        RECT 27.620 170.095 28.315 170.725 ;
        RECT 28.575 170.415 28.875 170.895 ;
        RECT 29.045 170.245 29.305 170.700 ;
        RECT 29.475 170.415 29.735 170.895 ;
        RECT 29.915 170.245 30.175 170.700 ;
        RECT 30.345 170.415 30.595 170.895 ;
        RECT 30.775 170.245 31.035 170.700 ;
        RECT 31.205 170.415 31.455 170.895 ;
        RECT 31.635 170.245 31.895 170.700 ;
        RECT 32.065 170.415 32.310 170.895 ;
        RECT 32.480 170.245 32.755 170.700 ;
        RECT 32.925 170.415 33.170 170.895 ;
        RECT 33.340 170.245 33.600 170.700 ;
        RECT 33.770 170.415 34.030 170.895 ;
        RECT 34.200 170.245 34.460 170.700 ;
        RECT 34.630 170.415 34.890 170.895 ;
        RECT 35.060 170.245 35.320 170.700 ;
        RECT 35.490 170.335 35.750 170.895 ;
        RECT 26.185 169.435 26.935 169.955 ;
        RECT 27.115 169.655 27.450 169.925 ;
        RECT 27.620 169.495 27.790 170.095 ;
        RECT 28.575 170.075 35.320 170.245 ;
        RECT 27.960 169.655 28.295 169.905 ;
        RECT 19.745 168.345 25.090 168.780 ;
        RECT 25.265 168.345 26.935 169.435 ;
        RECT 27.105 168.345 27.385 169.485 ;
        RECT 27.555 168.515 27.885 169.495 ;
        RECT 28.575 169.485 29.740 170.075 ;
        RECT 35.920 169.905 36.170 170.715 ;
        RECT 36.350 170.370 36.610 170.895 ;
        RECT 36.780 169.905 37.030 170.715 ;
        RECT 37.210 170.385 37.515 170.895 ;
        RECT 38.015 170.495 38.345 170.895 ;
        RECT 38.515 170.325 38.845 170.665 ;
        RECT 39.895 170.495 40.225 170.895 ;
        RECT 29.910 169.655 37.030 169.905 ;
        RECT 37.200 169.655 37.515 170.215 ;
        RECT 37.860 170.155 40.225 170.325 ;
        RECT 40.395 170.170 40.725 170.680 ;
        RECT 28.055 168.345 28.315 169.485 ;
        RECT 28.575 169.260 35.320 169.485 ;
        RECT 28.575 168.345 28.845 169.090 ;
        RECT 29.015 168.520 29.305 169.260 ;
        RECT 29.915 169.245 35.320 169.260 ;
        RECT 29.475 168.350 29.730 169.075 ;
        RECT 29.915 168.520 30.175 169.245 ;
        RECT 30.345 168.350 30.590 169.075 ;
        RECT 30.775 168.520 31.035 169.245 ;
        RECT 31.205 168.350 31.450 169.075 ;
        RECT 31.635 168.520 31.895 169.245 ;
        RECT 32.065 168.350 32.310 169.075 ;
        RECT 32.480 168.520 32.740 169.245 ;
        RECT 32.910 168.350 33.170 169.075 ;
        RECT 33.340 168.520 33.600 169.245 ;
        RECT 33.770 168.350 34.030 169.075 ;
        RECT 34.200 168.520 34.460 169.245 ;
        RECT 34.630 168.350 34.890 169.075 ;
        RECT 35.060 168.520 35.320 169.245 ;
        RECT 35.490 168.350 35.750 169.145 ;
        RECT 35.920 168.520 36.170 169.655 ;
        RECT 29.475 168.345 35.750 168.350 ;
        RECT 36.350 168.345 36.610 169.155 ;
        RECT 36.785 168.515 37.030 169.655 ;
        RECT 37.860 169.155 38.030 170.155 ;
        RECT 40.055 169.985 40.225 170.155 ;
        RECT 38.200 169.325 38.445 169.985 ;
        RECT 38.660 169.325 38.925 169.985 ;
        RECT 39.120 169.325 39.405 169.985 ;
        RECT 39.580 169.655 39.885 169.985 ;
        RECT 40.055 169.655 40.365 169.985 ;
        RECT 39.580 169.325 39.795 169.655 ;
        RECT 37.210 168.345 37.505 169.155 ;
        RECT 37.860 168.985 38.315 169.155 ;
        RECT 37.985 168.555 38.315 168.985 ;
        RECT 38.495 168.985 39.785 169.155 ;
        RECT 38.495 168.565 38.745 168.985 ;
        RECT 38.975 168.345 39.305 168.815 ;
        RECT 39.535 168.565 39.785 168.985 ;
        RECT 39.975 168.345 40.225 169.485 ;
        RECT 40.535 169.405 40.725 170.170 ;
        RECT 40.905 170.125 43.495 170.895 ;
        RECT 44.125 170.170 44.415 170.895 ;
        RECT 44.585 170.350 49.930 170.895 ;
        RECT 40.905 169.605 42.115 170.125 ;
        RECT 42.285 169.435 43.495 169.955 ;
        RECT 46.170 169.520 46.510 170.350 ;
        RECT 50.105 170.125 51.775 170.895 ;
        RECT 52.495 170.345 52.665 170.635 ;
        RECT 52.835 170.515 53.165 170.895 ;
        RECT 52.495 170.175 53.160 170.345 ;
        RECT 40.395 168.555 40.725 169.405 ;
        RECT 40.905 168.345 43.495 169.435 ;
        RECT 44.125 168.345 44.415 169.510 ;
        RECT 47.990 168.780 48.340 170.030 ;
        RECT 50.105 169.605 50.855 170.125 ;
        RECT 51.025 169.435 51.775 169.955 ;
        RECT 44.585 168.345 49.930 168.780 ;
        RECT 50.105 168.345 51.775 169.435 ;
        RECT 52.410 169.355 52.760 170.005 ;
        RECT 52.930 169.185 53.160 170.175 ;
        RECT 52.495 169.015 53.160 169.185 ;
        RECT 52.495 168.515 52.665 169.015 ;
        RECT 52.835 168.345 53.165 168.845 ;
        RECT 53.335 168.515 53.520 170.635 ;
        RECT 53.775 170.435 54.025 170.895 ;
        RECT 54.195 170.445 54.530 170.615 ;
        RECT 54.725 170.445 55.400 170.615 ;
        RECT 54.195 170.305 54.365 170.445 ;
        RECT 53.690 169.315 53.970 170.265 ;
        RECT 54.140 170.175 54.365 170.305 ;
        RECT 54.140 169.070 54.310 170.175 ;
        RECT 54.535 170.025 55.060 170.245 ;
        RECT 54.480 169.260 54.720 169.855 ;
        RECT 54.890 169.325 55.060 170.025 ;
        RECT 55.230 169.665 55.400 170.445 ;
        RECT 55.720 170.395 56.090 170.895 ;
        RECT 56.270 170.445 56.675 170.615 ;
        RECT 56.845 170.445 57.630 170.615 ;
        RECT 56.270 170.215 56.440 170.445 ;
        RECT 55.610 169.915 56.440 170.215 ;
        RECT 56.825 169.945 57.290 170.275 ;
        RECT 55.610 169.885 55.810 169.915 ;
        RECT 55.930 169.665 56.100 169.735 ;
        RECT 55.230 169.495 56.100 169.665 ;
        RECT 55.590 169.405 56.100 169.495 ;
        RECT 54.140 168.940 54.445 169.070 ;
        RECT 54.890 168.960 55.420 169.325 ;
        RECT 53.760 168.345 54.025 168.805 ;
        RECT 54.195 168.515 54.445 168.940 ;
        RECT 55.590 168.790 55.760 169.405 ;
        RECT 54.655 168.620 55.760 168.790 ;
        RECT 55.930 168.345 56.100 169.145 ;
        RECT 56.270 168.845 56.440 169.915 ;
        RECT 56.610 169.015 56.800 169.735 ;
        RECT 56.970 168.985 57.290 169.945 ;
        RECT 57.460 169.985 57.630 170.445 ;
        RECT 57.905 170.365 58.115 170.895 ;
        RECT 58.375 170.155 58.705 170.680 ;
        RECT 58.875 170.285 59.045 170.895 ;
        RECT 59.215 170.240 59.545 170.675 ;
        RECT 59.215 170.155 59.595 170.240 ;
        RECT 58.505 169.985 58.705 170.155 ;
        RECT 59.370 170.115 59.595 170.155 ;
        RECT 57.460 169.655 58.335 169.985 ;
        RECT 58.505 169.655 59.255 169.985 ;
        RECT 56.270 168.515 56.520 168.845 ;
        RECT 57.460 168.815 57.630 169.655 ;
        RECT 58.505 169.450 58.695 169.655 ;
        RECT 59.425 169.535 59.595 170.115 ;
        RECT 59.765 170.095 60.075 170.895 ;
        RECT 60.280 170.095 60.975 170.725 ;
        RECT 61.145 170.350 66.490 170.895 ;
        RECT 59.775 169.655 60.110 169.925 ;
        RECT 59.380 169.485 59.595 169.535 ;
        RECT 60.280 169.495 60.450 170.095 ;
        RECT 60.620 169.655 60.955 169.905 ;
        RECT 62.730 169.520 63.070 170.350 ;
        RECT 66.665 170.125 69.255 170.895 ;
        RECT 69.885 170.170 70.175 170.895 ;
        RECT 70.345 170.125 73.855 170.895 ;
        RECT 74.815 170.495 75.145 170.895 ;
        RECT 75.315 170.325 75.645 170.665 ;
        RECT 76.695 170.495 77.025 170.895 ;
        RECT 74.660 170.155 77.025 170.325 ;
        RECT 77.195 170.170 77.525 170.680 ;
        RECT 57.800 169.075 58.695 169.450 ;
        RECT 59.205 169.405 59.595 169.485 ;
        RECT 56.745 168.645 57.630 168.815 ;
        RECT 57.810 168.345 58.125 168.845 ;
        RECT 58.355 168.515 58.695 169.075 ;
        RECT 58.865 168.345 59.035 169.355 ;
        RECT 59.205 168.560 59.535 169.405 ;
        RECT 59.765 168.345 60.045 169.485 ;
        RECT 60.215 168.515 60.545 169.495 ;
        RECT 60.715 168.345 60.975 169.485 ;
        RECT 64.550 168.780 64.900 170.030 ;
        RECT 66.665 169.605 67.875 170.125 ;
        RECT 68.045 169.435 69.255 169.955 ;
        RECT 70.345 169.605 71.995 170.125 ;
        RECT 61.145 168.345 66.490 168.780 ;
        RECT 66.665 168.345 69.255 169.435 ;
        RECT 69.885 168.345 70.175 169.510 ;
        RECT 72.165 169.435 73.855 169.955 ;
        RECT 70.345 168.345 73.855 169.435 ;
        RECT 74.660 169.155 74.830 170.155 ;
        RECT 76.855 169.985 77.025 170.155 ;
        RECT 75.000 169.325 75.245 169.985 ;
        RECT 75.460 169.325 75.725 169.985 ;
        RECT 75.920 169.325 76.205 169.985 ;
        RECT 76.380 169.655 76.685 169.985 ;
        RECT 76.855 169.655 77.165 169.985 ;
        RECT 76.380 169.325 76.595 169.655 ;
        RECT 74.660 168.985 75.115 169.155 ;
        RECT 74.785 168.555 75.115 168.985 ;
        RECT 75.295 168.985 76.585 169.155 ;
        RECT 75.295 168.565 75.545 168.985 ;
        RECT 75.775 168.345 76.105 168.815 ;
        RECT 76.335 168.565 76.585 168.985 ;
        RECT 76.775 168.345 77.025 169.485 ;
        RECT 77.335 169.405 77.525 170.170 ;
        RECT 77.195 168.555 77.525 169.405 ;
        RECT 77.710 170.220 77.985 170.565 ;
        RECT 78.175 170.495 78.555 170.895 ;
        RECT 78.725 170.325 78.895 170.675 ;
        RECT 79.065 170.495 79.395 170.895 ;
        RECT 79.565 170.325 79.820 170.675 ;
        RECT 77.710 169.485 77.880 170.220 ;
        RECT 78.155 170.155 79.820 170.325 ;
        RECT 80.095 170.245 80.265 170.725 ;
        RECT 80.435 170.415 80.765 170.895 ;
        RECT 80.990 170.475 82.525 170.725 ;
        RECT 80.990 170.245 81.160 170.475 ;
        RECT 78.155 169.985 78.325 170.155 ;
        RECT 80.095 170.075 81.160 170.245 ;
        RECT 78.050 169.655 78.325 169.985 ;
        RECT 78.495 169.655 79.320 169.985 ;
        RECT 79.490 169.655 79.835 169.985 ;
        RECT 81.340 169.905 81.620 170.305 ;
        RECT 80.010 169.695 80.360 169.905 ;
        RECT 80.530 169.705 80.975 169.905 ;
        RECT 81.145 169.705 81.620 169.905 ;
        RECT 81.890 169.905 82.175 170.305 ;
        RECT 82.355 170.245 82.525 170.475 ;
        RECT 82.695 170.415 83.025 170.895 ;
        RECT 83.240 170.395 83.495 170.725 ;
        RECT 83.310 170.315 83.495 170.395 ;
        RECT 83.685 170.350 89.030 170.895 ;
        RECT 82.355 170.075 83.155 170.245 ;
        RECT 81.890 169.705 82.220 169.905 ;
        RECT 82.390 169.705 82.755 169.905 ;
        RECT 78.155 169.485 78.325 169.655 ;
        RECT 77.710 168.515 77.985 169.485 ;
        RECT 78.155 169.315 78.815 169.485 ;
        RECT 79.125 169.365 79.320 169.655 ;
        RECT 82.985 169.525 83.155 170.075 ;
        RECT 78.645 169.195 78.815 169.315 ;
        RECT 79.490 169.195 79.815 169.485 ;
        RECT 78.195 168.345 78.475 169.145 ;
        RECT 78.645 169.025 79.815 169.195 ;
        RECT 80.095 169.355 83.155 169.525 ;
        RECT 78.645 168.565 79.835 168.855 ;
        RECT 80.095 168.515 80.265 169.355 ;
        RECT 83.325 169.185 83.495 170.315 ;
        RECT 85.270 169.520 85.610 170.350 ;
        RECT 89.205 170.125 90.875 170.895 ;
        RECT 91.045 170.145 92.255 170.895 ;
        RECT 80.435 168.685 80.765 169.185 ;
        RECT 80.935 168.945 82.570 169.185 ;
        RECT 80.935 168.855 81.165 168.945 ;
        RECT 81.275 168.685 81.605 168.725 ;
        RECT 80.435 168.515 81.605 168.685 ;
        RECT 81.795 168.345 82.150 168.765 ;
        RECT 82.320 168.515 82.570 168.945 ;
        RECT 82.740 168.345 83.070 169.105 ;
        RECT 83.240 168.515 83.495 169.185 ;
        RECT 87.090 168.780 87.440 170.030 ;
        RECT 89.205 169.605 89.955 170.125 ;
        RECT 90.125 169.435 90.875 169.955 ;
        RECT 83.685 168.345 89.030 168.780 ;
        RECT 89.205 168.345 90.875 169.435 ;
        RECT 91.045 169.435 91.565 169.975 ;
        RECT 91.735 169.605 92.255 170.145 ;
        RECT 91.045 168.345 92.255 169.435 ;
        RECT 18.280 168.175 92.340 168.345 ;
        RECT 18.365 167.085 19.575 168.175 ;
        RECT 19.745 167.740 25.090 168.175 ;
        RECT 25.265 167.740 30.610 168.175 ;
        RECT 18.365 166.375 18.885 166.915 ;
        RECT 19.055 166.545 19.575 167.085 ;
        RECT 18.365 165.625 19.575 166.375 ;
        RECT 21.330 166.170 21.670 167.000 ;
        RECT 23.150 166.490 23.500 167.740 ;
        RECT 26.850 166.170 27.190 167.000 ;
        RECT 28.670 166.490 29.020 167.740 ;
        RECT 31.245 167.010 31.535 168.175 ;
        RECT 31.705 167.085 34.295 168.175 ;
        RECT 34.470 167.795 34.805 168.175 ;
        RECT 31.705 166.395 32.915 166.915 ;
        RECT 33.085 166.565 34.295 167.085 ;
        RECT 19.745 165.625 25.090 166.170 ;
        RECT 25.265 165.625 30.610 166.170 ;
        RECT 31.245 165.625 31.535 166.350 ;
        RECT 31.705 165.625 34.295 166.395 ;
        RECT 34.465 166.305 34.705 167.615 ;
        RECT 34.975 167.205 35.225 168.005 ;
        RECT 35.445 167.455 35.775 168.175 ;
        RECT 35.960 167.205 36.210 168.005 ;
        RECT 36.675 167.375 37.005 168.175 ;
        RECT 37.175 167.745 37.515 168.005 ;
        RECT 34.875 167.035 37.065 167.205 ;
        RECT 34.875 166.125 35.045 167.035 ;
        RECT 36.750 166.865 37.065 167.035 ;
        RECT 34.550 165.795 35.045 166.125 ;
        RECT 35.265 165.900 35.615 166.865 ;
        RECT 35.795 165.895 36.095 166.865 ;
        RECT 36.275 165.895 36.555 166.865 ;
        RECT 36.750 166.615 37.080 166.865 ;
        RECT 36.735 165.625 37.005 166.425 ;
        RECT 37.255 166.345 37.515 167.745 ;
        RECT 37.885 167.505 38.165 168.175 ;
        RECT 38.335 167.285 38.635 167.835 ;
        RECT 38.835 167.455 39.165 168.175 ;
        RECT 39.355 167.455 39.815 168.005 ;
        RECT 37.700 166.865 37.965 167.225 ;
        RECT 38.335 167.115 39.275 167.285 ;
        RECT 39.105 166.865 39.275 167.115 ;
        RECT 37.700 166.615 38.375 166.865 ;
        RECT 38.595 166.615 38.935 166.865 ;
        RECT 39.105 166.535 39.395 166.865 ;
        RECT 39.105 166.445 39.275 166.535 ;
        RECT 37.175 165.835 37.515 166.345 ;
        RECT 37.885 166.255 39.275 166.445 ;
        RECT 37.885 165.895 38.215 166.255 ;
        RECT 39.565 166.085 39.815 167.455 ;
        RECT 40.535 167.505 40.705 168.005 ;
        RECT 40.875 167.675 41.205 168.175 ;
        RECT 40.535 167.335 41.200 167.505 ;
        RECT 40.450 166.515 40.800 167.165 ;
        RECT 40.970 166.345 41.200 167.335 ;
        RECT 38.835 165.625 39.085 166.085 ;
        RECT 39.255 165.795 39.815 166.085 ;
        RECT 40.535 166.175 41.200 166.345 ;
        RECT 40.535 165.885 40.705 166.175 ;
        RECT 40.875 165.625 41.205 166.005 ;
        RECT 41.375 165.885 41.560 168.005 ;
        RECT 41.800 167.715 42.065 168.175 ;
        RECT 42.235 167.580 42.485 168.005 ;
        RECT 42.695 167.730 43.800 167.900 ;
        RECT 42.180 167.450 42.485 167.580 ;
        RECT 41.730 166.255 42.010 167.205 ;
        RECT 42.180 166.345 42.350 167.450 ;
        RECT 42.520 166.665 42.760 167.260 ;
        RECT 42.930 167.195 43.460 167.560 ;
        RECT 42.930 166.495 43.100 167.195 ;
        RECT 43.630 167.115 43.800 167.730 ;
        RECT 43.970 167.375 44.140 168.175 ;
        RECT 44.310 167.675 44.560 168.005 ;
        RECT 44.785 167.705 45.670 167.875 ;
        RECT 43.630 167.025 44.140 167.115 ;
        RECT 42.180 166.215 42.405 166.345 ;
        RECT 42.575 166.275 43.100 166.495 ;
        RECT 43.270 166.855 44.140 167.025 ;
        RECT 41.815 165.625 42.065 166.085 ;
        RECT 42.235 166.075 42.405 166.215 ;
        RECT 43.270 166.075 43.440 166.855 ;
        RECT 43.970 166.785 44.140 166.855 ;
        RECT 43.650 166.605 43.850 166.635 ;
        RECT 44.310 166.605 44.480 167.675 ;
        RECT 44.650 166.785 44.840 167.505 ;
        RECT 43.650 166.305 44.480 166.605 ;
        RECT 45.010 166.575 45.330 167.535 ;
        RECT 42.235 165.905 42.570 166.075 ;
        RECT 42.765 165.905 43.440 166.075 ;
        RECT 43.760 165.625 44.130 166.125 ;
        RECT 44.310 166.075 44.480 166.305 ;
        RECT 44.865 166.245 45.330 166.575 ;
        RECT 45.500 166.865 45.670 167.705 ;
        RECT 45.850 167.675 46.165 168.175 ;
        RECT 46.395 167.445 46.735 168.005 ;
        RECT 45.840 167.070 46.735 167.445 ;
        RECT 46.905 167.165 47.075 168.175 ;
        RECT 46.545 166.865 46.735 167.070 ;
        RECT 47.245 167.115 47.575 167.960 ;
        RECT 47.245 167.035 47.635 167.115 ;
        RECT 47.805 167.085 49.475 168.175 ;
        RECT 49.760 167.545 50.045 168.005 ;
        RECT 50.215 167.715 50.485 168.175 ;
        RECT 49.760 167.325 50.715 167.545 ;
        RECT 47.420 166.985 47.635 167.035 ;
        RECT 45.500 166.535 46.375 166.865 ;
        RECT 46.545 166.535 47.295 166.865 ;
        RECT 45.500 166.075 45.670 166.535 ;
        RECT 46.545 166.365 46.745 166.535 ;
        RECT 47.465 166.405 47.635 166.985 ;
        RECT 47.410 166.365 47.635 166.405 ;
        RECT 44.310 165.905 44.715 166.075 ;
        RECT 44.885 165.905 45.670 166.075 ;
        RECT 45.945 165.625 46.155 166.155 ;
        RECT 46.415 165.840 46.745 166.365 ;
        RECT 47.255 166.280 47.635 166.365 ;
        RECT 47.805 166.395 48.555 166.915 ;
        RECT 48.725 166.565 49.475 167.085 ;
        RECT 49.645 166.595 50.335 167.155 ;
        RECT 50.505 166.425 50.715 167.325 ;
        RECT 46.915 165.625 47.085 166.235 ;
        RECT 47.255 165.845 47.585 166.280 ;
        RECT 47.805 165.625 49.475 166.395 ;
        RECT 49.760 166.255 50.715 166.425 ;
        RECT 50.885 167.155 51.285 168.005 ;
        RECT 51.475 167.545 51.755 168.005 ;
        RECT 52.275 167.715 52.600 168.175 ;
        RECT 51.475 167.325 52.600 167.545 ;
        RECT 50.885 166.595 51.980 167.155 ;
        RECT 52.150 166.865 52.600 167.325 ;
        RECT 52.770 167.035 53.155 168.005 ;
        RECT 53.795 167.035 54.125 168.175 ;
        RECT 54.655 167.205 54.985 167.990 ;
        RECT 54.305 167.035 54.985 167.205 ;
        RECT 55.205 167.035 55.435 168.175 ;
        RECT 49.760 165.795 50.045 166.255 ;
        RECT 50.215 165.625 50.485 166.085 ;
        RECT 50.885 165.795 51.285 166.595 ;
        RECT 52.150 166.535 52.705 166.865 ;
        RECT 52.150 166.425 52.600 166.535 ;
        RECT 51.475 166.255 52.600 166.425 ;
        RECT 52.875 166.365 53.155 167.035 ;
        RECT 53.785 166.615 54.135 166.865 ;
        RECT 54.305 166.435 54.475 167.035 ;
        RECT 55.605 167.025 55.935 168.005 ;
        RECT 56.105 167.035 56.315 168.175 ;
        RECT 54.645 166.615 54.995 166.865 ;
        RECT 55.185 166.615 55.515 166.865 ;
        RECT 51.475 165.795 51.755 166.255 ;
        RECT 52.275 165.625 52.600 166.085 ;
        RECT 52.770 165.795 53.155 166.365 ;
        RECT 53.795 165.625 54.065 166.435 ;
        RECT 54.235 165.795 54.565 166.435 ;
        RECT 54.735 165.625 54.975 166.435 ;
        RECT 55.205 165.625 55.435 166.445 ;
        RECT 55.685 166.425 55.935 167.025 ;
        RECT 57.005 167.010 57.295 168.175 ;
        RECT 57.465 167.085 60.975 168.175 ;
        RECT 61.145 167.085 62.355 168.175 ;
        RECT 55.605 165.795 55.935 166.425 ;
        RECT 56.105 165.625 56.315 166.445 ;
        RECT 57.465 166.395 59.115 166.915 ;
        RECT 59.285 166.565 60.975 167.085 ;
        RECT 57.005 165.625 57.295 166.350 ;
        RECT 57.465 165.625 60.975 166.395 ;
        RECT 61.145 166.375 61.665 166.915 ;
        RECT 61.835 166.545 62.355 167.085 ;
        RECT 62.535 167.565 62.865 167.995 ;
        RECT 63.045 167.735 63.240 168.175 ;
        RECT 63.410 167.565 63.740 167.995 ;
        RECT 62.535 167.395 63.740 167.565 ;
        RECT 62.535 167.065 63.430 167.395 ;
        RECT 63.910 167.225 64.185 167.995 ;
        RECT 63.600 167.035 64.185 167.225 ;
        RECT 64.370 167.035 64.690 168.175 ;
        RECT 62.540 166.535 62.835 166.865 ;
        RECT 63.015 166.535 63.430 166.865 ;
        RECT 61.145 165.625 62.355 166.375 ;
        RECT 62.535 165.625 62.835 166.355 ;
        RECT 63.015 165.915 63.245 166.535 ;
        RECT 63.600 166.365 63.775 167.035 ;
        RECT 64.870 166.865 65.065 167.915 ;
        RECT 65.245 167.325 65.575 168.005 ;
        RECT 65.775 167.375 66.030 168.175 ;
        RECT 65.245 167.045 65.595 167.325 ;
        RECT 66.215 167.225 66.490 167.995 ;
        RECT 66.660 167.565 66.990 167.995 ;
        RECT 67.160 167.735 67.355 168.175 ;
        RECT 67.535 167.565 67.865 167.995 ;
        RECT 66.660 167.395 67.865 167.565 ;
        RECT 63.445 166.185 63.775 166.365 ;
        RECT 63.945 166.215 64.185 166.865 ;
        RECT 64.430 166.815 64.690 166.865 ;
        RECT 64.425 166.645 64.690 166.815 ;
        RECT 64.430 166.535 64.690 166.645 ;
        RECT 64.870 166.535 65.255 166.865 ;
        RECT 65.425 166.665 65.595 167.045 ;
        RECT 65.785 166.835 66.030 167.195 ;
        RECT 66.215 167.035 66.800 167.225 ;
        RECT 66.970 167.065 67.865 167.395 ;
        RECT 68.045 167.085 69.255 168.175 ;
        RECT 65.425 166.495 65.945 166.665 ;
        RECT 65.775 166.475 65.945 166.495 ;
        RECT 63.445 165.805 63.670 166.185 ;
        RECT 64.370 166.155 65.585 166.325 ;
        RECT 63.840 165.625 64.170 166.015 ;
        RECT 64.370 165.805 64.660 166.155 ;
        RECT 64.855 165.625 65.185 165.985 ;
        RECT 65.355 165.850 65.585 166.155 ;
        RECT 65.775 166.305 65.975 166.475 ;
        RECT 65.775 165.930 65.945 166.305 ;
        RECT 66.215 166.215 66.455 166.865 ;
        RECT 66.625 166.365 66.800 167.035 ;
        RECT 66.970 166.535 67.385 166.865 ;
        RECT 67.565 166.535 67.860 166.865 ;
        RECT 66.625 166.185 66.955 166.365 ;
        RECT 66.230 165.625 66.560 166.015 ;
        RECT 66.730 165.805 66.955 166.185 ;
        RECT 67.155 165.915 67.385 166.535 ;
        RECT 68.045 166.375 68.565 166.915 ;
        RECT 68.735 166.545 69.255 167.085 ;
        RECT 69.425 167.325 69.685 168.005 ;
        RECT 69.855 167.395 70.105 168.175 ;
        RECT 70.355 167.625 70.605 168.005 ;
        RECT 70.775 167.795 71.130 168.175 ;
        RECT 72.135 167.785 72.470 168.005 ;
        RECT 71.735 167.625 71.965 167.665 ;
        RECT 70.355 167.425 71.965 167.625 ;
        RECT 70.355 167.415 71.190 167.425 ;
        RECT 71.780 167.335 71.965 167.425 ;
        RECT 67.565 165.625 67.865 166.355 ;
        RECT 68.045 165.625 69.255 166.375 ;
        RECT 69.425 166.135 69.595 167.325 ;
        RECT 71.295 167.225 71.625 167.255 ;
        RECT 69.825 167.165 71.625 167.225 ;
        RECT 72.215 167.165 72.470 167.785 ;
        RECT 69.765 167.055 72.470 167.165 ;
        RECT 69.765 167.020 69.965 167.055 ;
        RECT 69.765 166.445 69.935 167.020 ;
        RECT 71.295 166.995 72.470 167.055 ;
        RECT 72.655 167.205 72.985 167.990 ;
        RECT 72.655 167.035 73.335 167.205 ;
        RECT 73.515 167.035 73.845 168.175 ;
        RECT 75.000 167.305 75.285 168.175 ;
        RECT 75.455 167.545 75.715 168.005 ;
        RECT 75.890 167.715 76.145 168.175 ;
        RECT 76.315 167.545 76.575 168.005 ;
        RECT 75.455 167.375 76.575 167.545 ;
        RECT 76.745 167.375 77.055 168.175 ;
        RECT 75.455 167.125 75.715 167.375 ;
        RECT 77.225 167.205 77.535 168.005 ;
        RECT 70.165 166.580 70.575 166.885 ;
        RECT 70.745 166.615 71.075 166.825 ;
        RECT 69.765 166.325 70.035 166.445 ;
        RECT 69.765 166.280 70.610 166.325 ;
        RECT 69.855 166.155 70.610 166.280 ;
        RECT 70.865 166.215 71.075 166.615 ;
        RECT 71.320 166.615 71.795 166.825 ;
        RECT 71.985 166.615 72.475 166.815 ;
        RECT 72.645 166.615 72.995 166.865 ;
        RECT 71.320 166.215 71.540 166.615 ;
        RECT 73.165 166.435 73.335 167.035 ;
        RECT 74.960 166.955 75.715 167.125 ;
        RECT 76.505 167.035 77.535 167.205 ;
        RECT 77.715 167.205 78.045 167.990 ;
        RECT 77.715 167.035 78.395 167.205 ;
        RECT 78.575 167.035 78.905 168.175 ;
        RECT 80.190 167.205 80.580 167.380 ;
        RECT 81.065 167.375 81.395 168.175 ;
        RECT 81.565 167.385 82.100 168.005 ;
        RECT 80.190 167.035 81.615 167.205 ;
        RECT 73.505 166.615 73.855 166.865 ;
        RECT 74.960 166.445 75.365 166.955 ;
        RECT 76.505 166.785 76.675 167.035 ;
        RECT 75.535 166.615 76.675 166.785 ;
        RECT 69.425 166.125 69.655 166.135 ;
        RECT 69.425 165.795 69.685 166.125 ;
        RECT 70.440 166.005 70.610 166.155 ;
        RECT 69.855 165.625 70.185 165.985 ;
        RECT 70.440 165.795 71.740 166.005 ;
        RECT 72.015 165.625 72.470 166.390 ;
        RECT 72.665 165.625 72.905 166.435 ;
        RECT 73.075 165.795 73.405 166.435 ;
        RECT 73.575 165.625 73.845 166.435 ;
        RECT 74.960 166.275 76.610 166.445 ;
        RECT 76.845 166.295 77.195 166.865 ;
        RECT 75.005 165.625 75.285 166.105 ;
        RECT 75.455 165.885 75.715 166.275 ;
        RECT 75.890 165.625 76.145 166.105 ;
        RECT 76.315 165.885 76.610 166.275 ;
        RECT 77.365 166.125 77.535 167.035 ;
        RECT 77.705 166.615 78.055 166.865 ;
        RECT 78.225 166.435 78.395 167.035 ;
        RECT 78.565 166.615 78.915 166.865 ;
        RECT 76.790 165.625 77.065 166.105 ;
        RECT 77.235 165.795 77.535 166.125 ;
        RECT 77.725 165.625 77.965 166.435 ;
        RECT 78.135 165.795 78.465 166.435 ;
        RECT 78.635 165.625 78.905 166.435 ;
        RECT 80.065 166.305 80.420 166.865 ;
        RECT 80.590 166.135 80.760 167.035 ;
        RECT 80.930 166.305 81.195 166.865 ;
        RECT 81.445 166.535 81.615 167.035 ;
        RECT 81.785 166.365 82.100 167.385 ;
        RECT 82.765 167.010 83.055 168.175 ;
        RECT 83.225 167.035 83.565 168.005 ;
        RECT 83.735 167.035 83.905 168.175 ;
        RECT 84.175 167.375 84.425 168.175 ;
        RECT 85.070 167.205 85.400 168.005 ;
        RECT 85.700 167.375 86.030 168.175 ;
        RECT 86.200 167.205 86.530 168.005 ;
        RECT 84.095 167.035 86.530 167.205 ;
        RECT 86.905 167.085 90.415 168.175 ;
        RECT 80.170 165.625 80.410 166.135 ;
        RECT 80.590 165.805 80.870 166.135 ;
        RECT 81.100 165.625 81.315 166.135 ;
        RECT 81.485 165.795 82.100 166.365 ;
        RECT 83.225 166.425 83.400 167.035 ;
        RECT 84.095 166.785 84.265 167.035 ;
        RECT 83.570 166.615 84.265 166.785 ;
        RECT 84.440 166.615 84.860 166.815 ;
        RECT 85.030 166.615 85.360 166.815 ;
        RECT 85.530 166.615 85.860 166.815 ;
        RECT 82.765 165.625 83.055 166.350 ;
        RECT 83.225 165.795 83.565 166.425 ;
        RECT 83.735 165.625 83.985 166.425 ;
        RECT 84.175 166.275 85.400 166.445 ;
        RECT 84.175 165.795 84.505 166.275 ;
        RECT 84.675 165.625 84.900 166.085 ;
        RECT 85.070 165.795 85.400 166.275 ;
        RECT 86.030 166.405 86.200 167.035 ;
        RECT 86.385 166.615 86.735 166.865 ;
        RECT 86.030 165.795 86.530 166.405 ;
        RECT 86.905 166.395 88.555 166.915 ;
        RECT 88.725 166.565 90.415 167.085 ;
        RECT 91.045 167.085 92.255 168.175 ;
        RECT 91.045 166.545 91.565 167.085 ;
        RECT 86.905 165.625 90.415 166.395 ;
        RECT 91.735 166.375 92.255 166.915 ;
        RECT 91.045 165.625 92.255 166.375 ;
        RECT 18.280 165.455 92.340 165.625 ;
        RECT 18.365 164.705 19.575 165.455 ;
        RECT 19.745 164.910 25.090 165.455 ;
        RECT 18.365 164.165 18.885 164.705 ;
        RECT 19.055 163.995 19.575 164.535 ;
        RECT 21.330 164.080 21.670 164.910 ;
        RECT 25.265 164.685 28.775 165.455 ;
        RECT 29.405 164.715 29.745 165.285 ;
        RECT 29.940 164.790 30.110 165.455 ;
        RECT 30.390 165.115 30.610 165.160 ;
        RECT 30.385 164.945 30.610 165.115 ;
        RECT 30.780 164.975 31.225 165.145 ;
        RECT 30.390 164.805 30.610 164.945 ;
        RECT 18.365 162.905 19.575 163.995 ;
        RECT 23.150 163.340 23.500 164.590 ;
        RECT 25.265 164.165 26.915 164.685 ;
        RECT 27.085 163.995 28.775 164.515 ;
        RECT 19.745 162.905 25.090 163.340 ;
        RECT 25.265 162.905 28.775 163.995 ;
        RECT 29.405 163.745 29.580 164.715 ;
        RECT 30.390 164.635 30.885 164.805 ;
        RECT 29.750 164.095 29.920 164.545 ;
        RECT 30.090 164.265 30.540 164.465 ;
        RECT 30.710 164.440 30.885 164.635 ;
        RECT 31.055 164.185 31.225 164.975 ;
        RECT 31.395 164.850 31.645 165.220 ;
        RECT 31.475 164.465 31.645 164.850 ;
        RECT 31.815 164.815 32.065 165.220 ;
        RECT 32.235 164.985 32.405 165.455 ;
        RECT 32.575 164.815 32.915 165.220 ;
        RECT 31.815 164.635 32.915 164.815 ;
        RECT 33.085 164.620 33.375 165.455 ;
        RECT 33.545 165.055 34.500 165.225 ;
        RECT 34.915 165.065 35.245 165.455 ;
        RECT 31.475 164.295 31.670 164.465 ;
        RECT 29.750 163.925 30.145 164.095 ;
        RECT 31.055 164.045 31.330 164.185 ;
        RECT 29.405 163.075 29.665 163.745 ;
        RECT 29.975 163.655 30.145 163.925 ;
        RECT 30.315 163.825 31.330 164.045 ;
        RECT 31.500 164.045 31.670 164.295 ;
        RECT 31.840 164.215 32.400 164.465 ;
        RECT 31.500 163.655 32.055 164.045 ;
        RECT 29.975 163.485 32.055 163.655 ;
        RECT 29.835 162.905 30.165 163.305 ;
        RECT 31.035 162.905 31.435 163.305 ;
        RECT 31.725 163.250 32.055 163.485 ;
        RECT 32.225 163.115 32.400 164.215 ;
        RECT 32.570 163.895 32.915 164.465 ;
        RECT 33.545 164.175 33.715 165.055 ;
        RECT 35.415 164.885 35.585 165.205 ;
        RECT 35.755 165.065 36.085 165.455 ;
        RECT 33.885 164.715 36.135 164.885 ;
        RECT 33.885 164.215 34.115 164.715 ;
        RECT 34.285 164.295 34.660 164.465 ;
        RECT 33.085 164.005 33.715 164.175 ;
        RECT 34.490 164.095 34.660 164.295 ;
        RECT 34.830 164.265 35.380 164.465 ;
        RECT 35.550 164.095 35.795 164.545 ;
        RECT 32.570 162.905 32.915 163.725 ;
        RECT 33.085 163.075 33.405 164.005 ;
        RECT 34.490 163.925 35.795 164.095 ;
        RECT 35.965 163.755 36.135 164.715 ;
        RECT 36.305 164.655 37.000 165.285 ;
        RECT 37.205 164.655 37.515 165.455 ;
        RECT 37.685 164.685 41.195 165.455 ;
        RECT 36.325 164.215 36.660 164.465 ;
        RECT 36.830 164.055 37.000 164.655 ;
        RECT 37.170 164.215 37.505 164.485 ;
        RECT 37.685 164.165 39.335 164.685 ;
        RECT 41.835 164.645 42.105 165.455 ;
        RECT 42.275 164.645 42.605 165.285 ;
        RECT 42.775 164.645 43.015 165.455 ;
        RECT 44.125 164.730 44.415 165.455 ;
        RECT 44.585 164.685 46.255 165.455 ;
        RECT 33.585 163.585 34.825 163.755 ;
        RECT 33.585 163.075 33.985 163.585 ;
        RECT 34.155 162.905 34.325 163.415 ;
        RECT 34.495 163.075 34.825 163.585 ;
        RECT 34.995 162.905 35.165 163.755 ;
        RECT 35.755 163.075 36.135 163.755 ;
        RECT 36.305 162.905 36.565 164.045 ;
        RECT 36.735 163.075 37.065 164.055 ;
        RECT 37.235 162.905 37.515 164.045 ;
        RECT 39.505 163.995 41.195 164.515 ;
        RECT 41.825 164.215 42.175 164.465 ;
        RECT 42.345 164.045 42.515 164.645 ;
        RECT 42.685 164.215 43.035 164.465 ;
        RECT 44.585 164.165 45.335 164.685 ;
        RECT 46.445 164.645 46.685 165.455 ;
        RECT 46.855 164.645 47.185 165.285 ;
        RECT 47.355 164.645 47.625 165.455 ;
        RECT 47.805 164.715 48.315 165.285 ;
        RECT 48.485 164.895 48.655 165.455 ;
        RECT 48.860 164.885 49.190 165.285 ;
        RECT 49.365 165.055 49.695 165.455 ;
        RECT 49.930 165.075 51.315 165.285 ;
        RECT 49.930 164.885 50.260 165.075 ;
        RECT 48.860 164.715 50.260 164.885 ;
        RECT 50.430 164.715 50.855 164.905 ;
        RECT 51.025 164.805 51.315 165.075 ;
        RECT 51.485 164.910 56.830 165.455 ;
        RECT 57.005 164.910 62.350 165.455 ;
        RECT 62.525 164.910 67.870 165.455 ;
        RECT 37.685 162.905 41.195 163.995 ;
        RECT 41.835 162.905 42.165 164.045 ;
        RECT 42.345 163.875 43.025 164.045 ;
        RECT 42.695 163.090 43.025 163.875 ;
        RECT 44.125 162.905 44.415 164.070 ;
        RECT 45.505 163.995 46.255 164.515 ;
        RECT 46.425 164.215 46.775 164.465 ;
        RECT 46.945 164.045 47.115 164.645 ;
        RECT 47.285 164.215 47.635 164.465 ;
        RECT 47.805 164.045 47.980 164.715 ;
        RECT 48.165 164.465 48.355 164.545 ;
        RECT 48.725 164.465 48.895 164.545 ;
        RECT 48.165 164.215 48.530 164.465 ;
        RECT 48.725 164.215 48.975 164.465 ;
        RECT 49.185 164.215 49.530 164.545 ;
        RECT 48.360 164.045 48.530 164.215 ;
        RECT 44.585 162.905 46.255 163.995 ;
        RECT 46.435 163.875 47.115 164.045 ;
        RECT 46.435 163.090 46.765 163.875 ;
        RECT 47.295 162.905 47.625 164.045 ;
        RECT 47.805 163.085 48.190 164.045 ;
        RECT 48.360 163.875 49.035 164.045 ;
        RECT 48.405 162.905 48.695 163.705 ;
        RECT 48.865 163.245 49.035 163.875 ;
        RECT 49.205 163.415 49.530 164.215 ;
        RECT 49.700 163.880 49.975 164.545 ;
        RECT 50.160 163.880 50.515 164.545 ;
        RECT 50.685 163.705 50.855 164.715 ;
        RECT 51.040 164.215 51.315 164.545 ;
        RECT 53.070 164.080 53.410 164.910 ;
        RECT 49.900 163.455 50.855 163.705 ;
        RECT 49.900 163.245 50.230 163.455 ;
        RECT 48.865 163.075 50.230 163.245 ;
        RECT 51.025 162.905 51.315 164.045 ;
        RECT 54.890 163.340 55.240 164.590 ;
        RECT 58.590 164.080 58.930 164.910 ;
        RECT 60.410 163.340 60.760 164.590 ;
        RECT 64.110 164.080 64.450 164.910 ;
        RECT 68.045 164.685 69.715 165.455 ;
        RECT 69.885 164.730 70.175 165.455 ;
        RECT 70.345 164.685 73.855 165.455 ;
        RECT 74.025 164.705 75.235 165.455 ;
        RECT 75.415 164.725 75.715 165.455 ;
        RECT 65.930 163.340 66.280 164.590 ;
        RECT 68.045 164.165 68.795 164.685 ;
        RECT 68.965 163.995 69.715 164.515 ;
        RECT 70.345 164.165 71.995 164.685 ;
        RECT 51.485 162.905 56.830 163.340 ;
        RECT 57.005 162.905 62.350 163.340 ;
        RECT 62.525 162.905 67.870 163.340 ;
        RECT 68.045 162.905 69.715 163.995 ;
        RECT 69.885 162.905 70.175 164.070 ;
        RECT 72.165 163.995 73.855 164.515 ;
        RECT 74.025 164.165 74.545 164.705 ;
        RECT 75.895 164.545 76.125 165.165 ;
        RECT 76.325 164.895 76.550 165.275 ;
        RECT 76.720 165.065 77.050 165.455 ;
        RECT 76.325 164.715 76.655 164.895 ;
        RECT 74.715 163.995 75.235 164.535 ;
        RECT 75.420 164.215 75.715 164.545 ;
        RECT 75.895 164.215 76.310 164.545 ;
        RECT 76.480 164.045 76.655 164.715 ;
        RECT 76.825 164.215 77.065 164.865 ;
        RECT 78.165 164.805 78.425 165.285 ;
        RECT 78.595 164.915 78.845 165.455 ;
        RECT 70.345 162.905 73.855 163.995 ;
        RECT 74.025 162.905 75.235 163.995 ;
        RECT 75.415 163.685 76.310 164.015 ;
        RECT 76.480 163.855 77.065 164.045 ;
        RECT 75.415 163.515 76.620 163.685 ;
        RECT 75.415 163.085 75.745 163.515 ;
        RECT 75.925 162.905 76.120 163.345 ;
        RECT 76.290 163.085 76.620 163.515 ;
        RECT 76.790 163.085 77.065 163.855 ;
        RECT 78.165 163.775 78.335 164.805 ;
        RECT 79.015 164.775 79.235 165.235 ;
        RECT 78.985 164.750 79.235 164.775 ;
        RECT 78.505 164.155 78.735 164.550 ;
        RECT 78.905 164.325 79.235 164.750 ;
        RECT 79.405 165.075 80.295 165.245 ;
        RECT 79.405 164.350 79.575 165.075 ;
        RECT 79.745 164.520 80.295 164.905 ;
        RECT 80.465 164.685 82.135 165.455 ;
        RECT 82.395 164.905 82.565 165.195 ;
        RECT 82.735 165.075 83.065 165.455 ;
        RECT 82.395 164.735 83.060 164.905 ;
        RECT 79.405 164.280 80.295 164.350 ;
        RECT 79.400 164.255 80.295 164.280 ;
        RECT 79.390 164.240 80.295 164.255 ;
        RECT 79.385 164.225 80.295 164.240 ;
        RECT 79.375 164.220 80.295 164.225 ;
        RECT 79.370 164.210 80.295 164.220 ;
        RECT 79.365 164.200 80.295 164.210 ;
        RECT 79.355 164.195 80.295 164.200 ;
        RECT 79.345 164.185 80.295 164.195 ;
        RECT 79.335 164.180 80.295 164.185 ;
        RECT 79.335 164.175 79.670 164.180 ;
        RECT 79.320 164.170 79.670 164.175 ;
        RECT 79.305 164.160 79.670 164.170 ;
        RECT 79.280 164.155 79.670 164.160 ;
        RECT 78.505 164.150 79.670 164.155 ;
        RECT 78.505 164.115 79.640 164.150 ;
        RECT 78.505 164.090 79.605 164.115 ;
        RECT 78.505 164.060 79.575 164.090 ;
        RECT 78.505 164.030 79.555 164.060 ;
        RECT 78.505 164.000 79.535 164.030 ;
        RECT 78.505 163.990 79.465 164.000 ;
        RECT 78.505 163.980 79.440 163.990 ;
        RECT 78.505 163.965 79.420 163.980 ;
        RECT 78.505 163.950 79.400 163.965 ;
        RECT 78.610 163.940 79.395 163.950 ;
        RECT 78.610 163.905 79.380 163.940 ;
        RECT 78.165 163.075 78.440 163.775 ;
        RECT 78.610 163.655 79.365 163.905 ;
        RECT 79.535 163.585 79.865 163.830 ;
        RECT 80.035 163.730 80.295 164.180 ;
        RECT 80.465 164.165 81.215 164.685 ;
        RECT 81.385 163.995 82.135 164.515 ;
        RECT 79.680 163.560 79.865 163.585 ;
        RECT 79.680 163.460 80.295 163.560 ;
        RECT 78.610 162.905 78.865 163.450 ;
        RECT 79.035 163.075 79.515 163.415 ;
        RECT 79.690 162.905 80.295 163.460 ;
        RECT 80.465 162.905 82.135 163.995 ;
        RECT 82.310 163.915 82.660 164.565 ;
        RECT 82.830 163.745 83.060 164.735 ;
        RECT 82.395 163.575 83.060 163.745 ;
        RECT 82.395 163.075 82.565 163.575 ;
        RECT 82.735 162.905 83.065 163.405 ;
        RECT 83.235 163.075 83.460 165.195 ;
        RECT 83.675 164.995 83.925 165.455 ;
        RECT 84.110 165.005 84.440 165.175 ;
        RECT 84.620 165.005 85.370 165.175 ;
        RECT 83.660 163.875 83.940 164.475 ;
        RECT 84.110 163.475 84.280 165.005 ;
        RECT 84.450 164.505 85.030 164.835 ;
        RECT 84.450 163.635 84.690 164.505 ;
        RECT 85.200 164.225 85.370 165.005 ;
        RECT 85.620 164.955 85.990 165.455 ;
        RECT 86.170 165.005 86.630 165.175 ;
        RECT 86.860 165.005 87.530 165.175 ;
        RECT 86.170 164.775 86.340 165.005 ;
        RECT 85.540 164.475 86.340 164.775 ;
        RECT 86.510 164.505 87.060 164.835 ;
        RECT 85.540 164.445 85.710 164.475 ;
        RECT 85.830 164.225 86.000 164.295 ;
        RECT 85.200 164.055 86.000 164.225 ;
        RECT 85.490 163.965 86.000 164.055 ;
        RECT 84.880 163.530 85.320 163.885 ;
        RECT 83.660 162.905 83.925 163.365 ;
        RECT 84.110 163.100 84.345 163.475 ;
        RECT 85.490 163.350 85.660 163.965 ;
        RECT 84.590 163.180 85.660 163.350 ;
        RECT 85.830 162.905 86.000 163.705 ;
        RECT 86.170 163.405 86.340 164.475 ;
        RECT 86.510 163.575 86.700 164.295 ;
        RECT 86.870 163.965 87.060 164.505 ;
        RECT 87.360 164.465 87.530 165.005 ;
        RECT 87.845 164.925 88.015 165.455 ;
        RECT 88.310 164.805 88.670 165.245 ;
        RECT 88.845 164.975 89.015 165.455 ;
        RECT 89.205 164.810 89.540 165.235 ;
        RECT 89.715 164.980 89.885 165.455 ;
        RECT 90.060 164.810 90.395 165.235 ;
        RECT 90.565 164.980 90.735 165.455 ;
        RECT 88.310 164.635 88.810 164.805 ;
        RECT 89.205 164.640 90.875 164.810 ;
        RECT 91.045 164.705 92.255 165.455 ;
        RECT 88.640 164.465 88.810 164.635 ;
        RECT 87.360 164.295 88.450 164.465 ;
        RECT 88.640 164.295 90.460 164.465 ;
        RECT 86.870 163.635 87.190 163.965 ;
        RECT 86.170 163.075 86.420 163.405 ;
        RECT 87.360 163.375 87.530 164.295 ;
        RECT 88.640 164.040 88.810 164.295 ;
        RECT 90.630 164.075 90.875 164.640 ;
        RECT 87.700 163.870 88.810 164.040 ;
        RECT 89.205 163.905 90.875 164.075 ;
        RECT 91.045 163.995 91.565 164.535 ;
        RECT 91.735 164.165 92.255 164.705 ;
        RECT 87.700 163.710 88.560 163.870 ;
        RECT 86.645 163.205 87.530 163.375 ;
        RECT 87.710 162.905 87.925 163.405 ;
        RECT 88.390 163.085 88.560 163.710 ;
        RECT 88.845 162.905 89.025 163.685 ;
        RECT 89.205 163.145 89.540 163.905 ;
        RECT 89.720 162.905 89.890 163.735 ;
        RECT 90.060 163.145 90.390 163.905 ;
        RECT 90.560 162.905 90.730 163.735 ;
        RECT 91.045 162.905 92.255 163.995 ;
        RECT 18.280 162.735 92.340 162.905 ;
        RECT 18.365 161.645 19.575 162.735 ;
        RECT 19.745 161.645 22.335 162.735 ;
        RECT 22.595 162.065 22.765 162.565 ;
        RECT 22.935 162.235 23.265 162.735 ;
        RECT 22.595 161.895 23.260 162.065 ;
        RECT 18.365 160.935 18.885 161.475 ;
        RECT 19.055 161.105 19.575 161.645 ;
        RECT 19.745 160.955 20.955 161.475 ;
        RECT 21.125 161.125 22.335 161.645 ;
        RECT 22.510 161.075 22.860 161.725 ;
        RECT 18.365 160.185 19.575 160.935 ;
        RECT 19.745 160.185 22.335 160.955 ;
        RECT 23.030 160.905 23.260 161.895 ;
        RECT 22.595 160.735 23.260 160.905 ;
        RECT 22.595 160.445 22.765 160.735 ;
        RECT 22.935 160.185 23.265 160.565 ;
        RECT 23.435 160.445 23.620 162.565 ;
        RECT 23.860 162.275 24.125 162.735 ;
        RECT 24.295 162.140 24.545 162.565 ;
        RECT 24.755 162.290 25.860 162.460 ;
        RECT 24.240 162.010 24.545 162.140 ;
        RECT 23.790 160.815 24.070 161.765 ;
        RECT 24.240 160.905 24.410 162.010 ;
        RECT 24.580 161.225 24.820 161.820 ;
        RECT 24.990 161.755 25.520 162.120 ;
        RECT 24.990 161.055 25.160 161.755 ;
        RECT 25.690 161.675 25.860 162.290 ;
        RECT 26.030 161.935 26.200 162.735 ;
        RECT 26.370 162.235 26.620 162.565 ;
        RECT 26.845 162.265 27.730 162.435 ;
        RECT 25.690 161.585 26.200 161.675 ;
        RECT 24.240 160.775 24.465 160.905 ;
        RECT 24.635 160.835 25.160 161.055 ;
        RECT 25.330 161.415 26.200 161.585 ;
        RECT 23.875 160.185 24.125 160.645 ;
        RECT 24.295 160.635 24.465 160.775 ;
        RECT 25.330 160.635 25.500 161.415 ;
        RECT 26.030 161.345 26.200 161.415 ;
        RECT 25.710 161.165 25.910 161.195 ;
        RECT 26.370 161.165 26.540 162.235 ;
        RECT 26.710 161.345 26.900 162.065 ;
        RECT 25.710 160.865 26.540 161.165 ;
        RECT 27.070 161.135 27.390 162.095 ;
        RECT 24.295 160.465 24.630 160.635 ;
        RECT 24.825 160.465 25.500 160.635 ;
        RECT 25.820 160.185 26.190 160.685 ;
        RECT 26.370 160.635 26.540 160.865 ;
        RECT 26.925 160.805 27.390 161.135 ;
        RECT 27.560 161.425 27.730 162.265 ;
        RECT 27.910 162.235 28.225 162.735 ;
        RECT 28.455 162.005 28.795 162.565 ;
        RECT 27.900 161.630 28.795 162.005 ;
        RECT 28.965 161.725 29.135 162.735 ;
        RECT 28.605 161.425 28.795 161.630 ;
        RECT 29.305 161.675 29.635 162.520 ;
        RECT 29.875 161.765 30.205 162.550 ;
        RECT 29.305 161.595 29.695 161.675 ;
        RECT 29.875 161.595 30.555 161.765 ;
        RECT 30.735 161.595 31.065 162.735 ;
        RECT 29.480 161.545 29.695 161.595 ;
        RECT 27.560 161.095 28.435 161.425 ;
        RECT 28.605 161.095 29.355 161.425 ;
        RECT 27.560 160.635 27.730 161.095 ;
        RECT 28.605 160.925 28.805 161.095 ;
        RECT 29.525 160.965 29.695 161.545 ;
        RECT 29.865 161.175 30.215 161.425 ;
        RECT 30.385 160.995 30.555 161.595 ;
        RECT 31.245 161.570 31.535 162.735 ;
        RECT 31.705 161.645 34.295 162.735 ;
        RECT 30.725 161.175 31.075 161.425 ;
        RECT 29.470 160.925 29.695 160.965 ;
        RECT 26.370 160.465 26.775 160.635 ;
        RECT 26.945 160.465 27.730 160.635 ;
        RECT 28.005 160.185 28.215 160.715 ;
        RECT 28.475 160.400 28.805 160.925 ;
        RECT 29.315 160.840 29.695 160.925 ;
        RECT 28.975 160.185 29.145 160.795 ;
        RECT 29.315 160.405 29.645 160.840 ;
        RECT 29.885 160.185 30.125 160.995 ;
        RECT 30.295 160.355 30.625 160.995 ;
        RECT 30.795 160.185 31.065 160.995 ;
        RECT 31.705 160.955 32.915 161.475 ;
        RECT 33.085 161.125 34.295 161.645 ;
        RECT 34.925 161.595 35.200 162.565 ;
        RECT 35.410 161.935 35.690 162.735 ;
        RECT 35.860 162.225 37.475 162.555 ;
        RECT 35.860 161.885 37.035 162.055 ;
        RECT 35.860 161.765 36.030 161.885 ;
        RECT 35.370 161.595 36.030 161.765 ;
        RECT 31.245 160.185 31.535 160.910 ;
        RECT 31.705 160.185 34.295 160.955 ;
        RECT 34.925 160.860 35.095 161.595 ;
        RECT 35.370 161.425 35.540 161.595 ;
        RECT 36.290 161.425 36.535 161.715 ;
        RECT 36.705 161.595 37.035 161.885 ;
        RECT 37.295 161.425 37.465 161.985 ;
        RECT 37.715 161.595 37.975 162.735 ;
        RECT 38.155 161.765 38.485 162.550 ;
        RECT 38.155 161.595 38.835 161.765 ;
        RECT 39.015 161.595 39.345 162.735 ;
        RECT 39.525 161.645 43.035 162.735 ;
        RECT 35.265 161.095 35.540 161.425 ;
        RECT 35.710 161.095 36.535 161.425 ;
        RECT 36.750 161.095 37.465 161.425 ;
        RECT 37.635 161.175 37.970 161.425 ;
        RECT 38.145 161.175 38.495 161.425 ;
        RECT 35.370 160.925 35.540 161.095 ;
        RECT 37.215 161.005 37.465 161.095 ;
        RECT 34.925 160.515 35.200 160.860 ;
        RECT 35.370 160.755 37.035 160.925 ;
        RECT 35.390 160.185 35.765 160.585 ;
        RECT 35.935 160.405 36.105 160.755 ;
        RECT 36.275 160.185 36.605 160.585 ;
        RECT 36.775 160.355 37.035 160.755 ;
        RECT 37.215 160.585 37.545 161.005 ;
        RECT 37.715 160.185 37.975 161.005 ;
        RECT 38.665 160.995 38.835 161.595 ;
        RECT 39.005 161.175 39.355 161.425 ;
        RECT 38.165 160.185 38.405 160.995 ;
        RECT 38.575 160.355 38.905 160.995 ;
        RECT 39.075 160.185 39.345 160.995 ;
        RECT 39.525 160.955 41.175 161.475 ;
        RECT 41.345 161.125 43.035 161.645 ;
        RECT 44.125 161.595 44.510 162.555 ;
        RECT 44.725 161.935 45.015 162.735 ;
        RECT 45.185 162.395 46.550 162.565 ;
        RECT 45.185 161.765 45.355 162.395 ;
        RECT 44.680 161.595 45.355 161.765 ;
        RECT 39.525 160.185 43.035 160.955 ;
        RECT 44.125 160.925 44.300 161.595 ;
        RECT 44.680 161.425 44.850 161.595 ;
        RECT 45.525 161.425 45.850 162.225 ;
        RECT 46.220 162.185 46.550 162.395 ;
        RECT 46.220 161.935 47.175 162.185 ;
        RECT 44.485 161.175 44.850 161.425 ;
        RECT 45.045 161.175 45.295 161.425 ;
        RECT 44.485 161.095 44.675 161.175 ;
        RECT 45.045 161.095 45.215 161.175 ;
        RECT 45.505 161.095 45.850 161.425 ;
        RECT 46.020 161.095 46.295 161.760 ;
        RECT 46.480 161.095 46.835 161.760 ;
        RECT 47.005 160.925 47.175 161.935 ;
        RECT 47.345 161.595 47.635 162.735 ;
        RECT 47.815 162.355 48.145 162.735 ;
        RECT 47.360 161.095 47.635 161.425 ;
        RECT 44.125 160.355 44.635 160.925 ;
        RECT 45.180 160.755 46.580 160.925 ;
        RECT 44.805 160.185 44.975 160.745 ;
        RECT 45.180 160.355 45.510 160.755 ;
        RECT 45.685 160.185 46.015 160.585 ;
        RECT 46.250 160.565 46.580 160.755 ;
        RECT 46.750 160.735 47.175 160.925 ;
        RECT 47.845 160.855 48.050 162.175 ;
        RECT 48.320 161.765 48.570 162.565 ;
        RECT 48.790 162.015 49.120 162.735 ;
        RECT 49.305 161.765 49.555 162.565 ;
        RECT 49.955 161.935 50.285 162.735 ;
        RECT 50.455 162.395 50.790 162.565 ;
        RECT 50.455 162.225 50.795 162.395 ;
        RECT 48.220 161.595 50.275 161.765 ;
        RECT 50.455 161.595 50.790 162.225 ;
        RECT 50.965 161.935 51.295 162.735 ;
        RECT 51.545 161.595 51.755 162.735 ;
        RECT 47.345 160.565 47.635 160.835 ;
        RECT 48.220 160.685 48.390 161.595 ;
        RECT 46.250 160.355 47.635 160.565 ;
        RECT 47.895 160.355 48.390 160.685 ;
        RECT 48.610 160.520 48.965 161.425 ;
        RECT 49.140 161.405 49.310 161.425 ;
        RECT 49.140 160.515 49.440 161.405 ;
        RECT 49.620 160.515 49.880 161.425 ;
        RECT 50.050 161.415 50.275 161.595 ;
        RECT 50.050 161.175 50.445 161.415 ;
        RECT 50.050 160.185 50.285 160.990 ;
        RECT 50.615 160.905 50.790 161.595 ;
        RECT 51.925 161.585 52.255 162.565 ;
        RECT 52.425 161.595 52.655 162.735 ;
        RECT 53.325 162.225 53.625 162.735 ;
        RECT 53.795 162.055 54.125 162.565 ;
        RECT 54.295 162.225 54.925 162.735 ;
        RECT 55.505 162.225 55.885 162.395 ;
        RECT 56.055 162.225 56.355 162.735 ;
        RECT 55.715 162.055 55.885 162.225 ;
        RECT 53.325 161.885 55.545 162.055 ;
        RECT 50.455 160.440 50.790 160.905 ;
        RECT 50.455 160.395 50.785 160.440 ;
        RECT 50.975 160.185 51.305 160.910 ;
        RECT 51.545 160.185 51.755 161.005 ;
        RECT 51.925 160.985 52.175 161.585 ;
        RECT 52.345 161.175 52.675 161.425 ;
        RECT 51.925 160.355 52.255 160.985 ;
        RECT 52.425 160.185 52.655 161.005 ;
        RECT 53.325 160.925 53.495 161.885 ;
        RECT 53.665 161.545 55.205 161.715 ;
        RECT 53.665 161.095 53.910 161.545 ;
        RECT 54.170 161.175 54.865 161.375 ;
        RECT 55.035 161.345 55.205 161.545 ;
        RECT 55.375 161.685 55.545 161.885 ;
        RECT 55.715 161.855 56.375 162.055 ;
        RECT 55.375 161.515 56.035 161.685 ;
        RECT 55.035 161.175 55.635 161.345 ;
        RECT 55.865 161.095 56.035 161.515 ;
        RECT 53.325 160.380 53.790 160.925 ;
        RECT 54.295 160.185 54.465 161.005 ;
        RECT 54.635 160.925 55.545 161.005 ;
        RECT 56.205 160.925 56.375 161.855 ;
        RECT 57.005 161.570 57.295 162.735 ;
        RECT 57.465 161.915 57.810 162.735 ;
        RECT 57.465 161.175 57.810 161.745 ;
        RECT 57.980 161.425 58.155 162.525 ;
        RECT 58.325 162.155 58.655 162.390 ;
        RECT 58.945 162.335 59.345 162.735 ;
        RECT 60.215 162.335 60.545 162.735 ;
        RECT 58.325 161.985 60.405 162.155 ;
        RECT 58.325 161.595 58.880 161.985 ;
        RECT 57.980 161.175 58.540 161.425 ;
        RECT 58.710 161.345 58.880 161.595 ;
        RECT 59.050 161.595 60.065 161.815 ;
        RECT 60.235 161.715 60.405 161.985 ;
        RECT 60.715 161.895 60.975 162.565 ;
        RECT 59.050 161.455 59.325 161.595 ;
        RECT 60.235 161.545 60.630 161.715 ;
        RECT 58.710 161.175 58.905 161.345 ;
        RECT 54.635 160.835 55.885 160.925 ;
        RECT 54.635 160.355 54.965 160.835 ;
        RECT 55.375 160.755 55.885 160.835 ;
        RECT 55.135 160.185 55.485 160.575 ;
        RECT 55.655 160.355 55.885 160.755 ;
        RECT 56.055 160.445 56.375 160.925 ;
        RECT 57.005 160.185 57.295 160.910 ;
        RECT 57.465 160.825 58.565 161.005 ;
        RECT 57.465 160.420 57.805 160.825 ;
        RECT 57.975 160.185 58.145 160.655 ;
        RECT 58.315 160.420 58.565 160.825 ;
        RECT 58.735 160.790 58.905 161.175 ;
        RECT 58.735 160.420 58.985 160.790 ;
        RECT 59.155 160.665 59.325 161.455 ;
        RECT 59.495 161.005 59.670 161.200 ;
        RECT 59.840 161.175 60.290 161.375 ;
        RECT 60.460 161.095 60.630 161.545 ;
        RECT 59.495 160.835 59.990 161.005 ;
        RECT 60.800 160.925 60.975 161.895 ;
        RECT 59.770 160.695 59.990 160.835 ;
        RECT 59.155 160.495 59.600 160.665 ;
        RECT 59.770 160.525 59.995 160.695 ;
        RECT 59.770 160.480 59.990 160.525 ;
        RECT 60.270 160.185 60.440 160.850 ;
        RECT 60.635 160.355 60.975 160.925 ;
        RECT 62.065 161.130 62.345 162.565 ;
        RECT 62.515 161.960 63.225 162.735 ;
        RECT 63.395 161.790 63.725 162.565 ;
        RECT 62.575 161.575 63.725 161.790 ;
        RECT 62.065 160.355 62.405 161.130 ;
        RECT 62.575 161.005 62.860 161.575 ;
        RECT 63.045 161.175 63.515 161.405 ;
        RECT 63.920 161.375 64.135 162.490 ;
        RECT 64.315 162.015 64.645 162.735 ;
        RECT 64.835 161.785 65.110 162.555 ;
        RECT 65.280 162.125 65.610 162.555 ;
        RECT 65.780 162.295 65.975 162.735 ;
        RECT 66.155 162.125 66.485 162.555 ;
        RECT 65.280 161.955 66.485 162.125 ;
        RECT 64.425 161.375 64.655 161.715 ;
        RECT 64.835 161.595 65.420 161.785 ;
        RECT 65.590 161.625 66.485 161.955 ;
        RECT 66.665 161.645 69.255 162.735 ;
        RECT 63.685 161.195 64.135 161.375 ;
        RECT 63.685 161.175 64.015 161.195 ;
        RECT 64.325 161.175 64.655 161.375 ;
        RECT 62.575 160.815 63.285 161.005 ;
        RECT 62.985 160.675 63.285 160.815 ;
        RECT 63.475 160.815 64.655 161.005 ;
        RECT 63.475 160.735 63.805 160.815 ;
        RECT 62.985 160.665 63.300 160.675 ;
        RECT 62.985 160.655 63.310 160.665 ;
        RECT 62.985 160.650 63.320 160.655 ;
        RECT 62.575 160.185 62.745 160.645 ;
        RECT 62.985 160.640 63.325 160.650 ;
        RECT 62.985 160.635 63.330 160.640 ;
        RECT 62.985 160.625 63.335 160.635 ;
        RECT 62.985 160.620 63.340 160.625 ;
        RECT 62.985 160.355 63.345 160.620 ;
        RECT 63.975 160.185 64.145 160.645 ;
        RECT 64.315 160.355 64.655 160.815 ;
        RECT 64.835 160.775 65.075 161.425 ;
        RECT 65.245 160.925 65.420 161.595 ;
        RECT 65.590 161.095 66.005 161.425 ;
        RECT 66.185 161.095 66.480 161.425 ;
        RECT 65.245 160.745 65.575 160.925 ;
        RECT 64.850 160.185 65.180 160.575 ;
        RECT 65.350 160.365 65.575 160.745 ;
        RECT 65.775 160.475 66.005 161.095 ;
        RECT 66.665 160.955 67.875 161.475 ;
        RECT 68.045 161.125 69.255 161.645 ;
        RECT 69.890 161.595 70.210 162.735 ;
        RECT 70.390 161.425 70.585 162.475 ;
        RECT 70.765 161.885 71.095 162.565 ;
        RECT 71.295 161.935 71.550 162.735 ;
        RECT 70.765 161.605 71.115 161.885 ;
        RECT 69.950 161.375 70.210 161.425 ;
        RECT 69.945 161.205 70.210 161.375 ;
        RECT 69.950 161.095 70.210 161.205 ;
        RECT 70.390 161.095 70.775 161.425 ;
        RECT 70.945 161.225 71.115 161.605 ;
        RECT 71.305 161.395 71.550 161.755 ;
        RECT 71.725 161.595 72.005 162.735 ;
        RECT 72.175 161.585 72.505 162.565 ;
        RECT 72.675 161.595 72.935 162.735 ;
        RECT 73.105 161.645 76.615 162.735 ;
        RECT 76.785 161.645 77.995 162.735 ;
        RECT 70.945 161.055 71.465 161.225 ;
        RECT 71.735 161.155 72.070 161.425 ;
        RECT 66.185 160.185 66.485 160.915 ;
        RECT 66.665 160.185 69.255 160.955 ;
        RECT 69.890 160.715 71.105 160.885 ;
        RECT 69.890 160.365 70.180 160.715 ;
        RECT 70.375 160.185 70.705 160.545 ;
        RECT 70.875 160.410 71.105 160.715 ;
        RECT 71.295 160.695 71.465 161.055 ;
        RECT 72.240 160.985 72.410 161.585 ;
        RECT 72.580 161.175 72.915 161.425 ;
        RECT 71.295 160.525 71.495 160.695 ;
        RECT 71.295 160.490 71.465 160.525 ;
        RECT 71.725 160.185 72.035 160.985 ;
        RECT 72.240 160.355 72.935 160.985 ;
        RECT 73.105 160.955 74.755 161.475 ;
        RECT 74.925 161.125 76.615 161.645 ;
        RECT 73.105 160.185 76.615 160.955 ;
        RECT 76.785 160.935 77.305 161.475 ;
        RECT 77.475 161.105 77.995 161.645 ;
        RECT 78.165 161.580 78.505 162.565 ;
        RECT 78.675 162.305 79.085 162.735 ;
        RECT 79.830 162.315 80.160 162.735 ;
        RECT 80.330 162.135 80.655 162.565 ;
        RECT 78.675 161.965 80.655 162.135 ;
        RECT 76.785 160.185 77.995 160.935 ;
        RECT 78.165 160.925 78.420 161.580 ;
        RECT 78.675 161.425 78.940 161.965 ;
        RECT 79.155 161.625 79.780 161.795 ;
        RECT 78.590 161.095 78.940 161.425 ;
        RECT 79.110 161.095 79.440 161.425 ;
        RECT 79.610 160.925 79.780 161.625 ;
        RECT 78.165 160.550 78.525 160.925 ;
        RECT 78.225 160.525 78.395 160.550 ;
        RECT 78.790 160.185 78.960 160.925 ;
        RECT 79.240 160.755 79.780 160.925 ;
        RECT 79.950 161.555 80.655 161.965 ;
        RECT 81.130 161.635 81.460 162.735 ;
        RECT 82.765 161.570 83.055 162.735 ;
        RECT 83.225 161.595 83.610 162.565 ;
        RECT 83.780 162.275 84.105 162.735 ;
        RECT 84.625 162.105 84.905 162.565 ;
        RECT 83.780 161.885 84.905 162.105 ;
        RECT 79.240 160.550 79.410 160.755 ;
        RECT 79.950 160.355 80.120 161.555 ;
        RECT 80.290 161.175 80.860 161.385 ;
        RECT 81.030 161.175 81.675 161.385 ;
        RECT 80.350 160.835 81.520 161.005 ;
        RECT 83.225 160.925 83.505 161.595 ;
        RECT 83.780 161.425 84.230 161.885 ;
        RECT 85.095 161.715 85.495 162.565 ;
        RECT 85.895 162.275 86.165 162.735 ;
        RECT 86.335 162.105 86.620 162.565 ;
        RECT 83.675 161.095 84.230 161.425 ;
        RECT 84.400 161.155 85.495 161.715 ;
        RECT 83.780 160.985 84.230 161.095 ;
        RECT 80.350 160.355 80.680 160.835 ;
        RECT 80.850 160.185 81.020 160.655 ;
        RECT 81.190 160.370 81.520 160.835 ;
        RECT 82.765 160.185 83.055 160.910 ;
        RECT 83.225 160.355 83.610 160.925 ;
        RECT 83.780 160.815 84.905 160.985 ;
        RECT 83.780 160.185 84.105 160.645 ;
        RECT 84.625 160.355 84.905 160.815 ;
        RECT 85.095 160.355 85.495 161.155 ;
        RECT 85.665 161.885 86.620 162.105 ;
        RECT 86.905 162.305 87.245 162.565 ;
        RECT 85.665 160.985 85.875 161.885 ;
        RECT 86.045 161.155 86.735 161.715 ;
        RECT 85.665 160.815 86.620 160.985 ;
        RECT 85.895 160.185 86.165 160.645 ;
        RECT 86.335 160.355 86.620 160.815 ;
        RECT 86.905 160.905 87.165 162.305 ;
        RECT 87.415 161.935 87.745 162.735 ;
        RECT 88.210 161.765 88.460 162.565 ;
        RECT 88.645 162.015 88.975 162.735 ;
        RECT 89.195 161.765 89.445 162.565 ;
        RECT 89.615 162.355 89.950 162.735 ;
        RECT 87.355 161.595 89.545 161.765 ;
        RECT 87.355 161.425 87.670 161.595 ;
        RECT 87.340 161.175 87.670 161.425 ;
        RECT 86.905 160.395 87.245 160.905 ;
        RECT 87.415 160.185 87.685 160.985 ;
        RECT 87.865 160.455 88.145 161.425 ;
        RECT 88.325 160.455 88.625 161.425 ;
        RECT 88.805 160.460 89.155 161.425 ;
        RECT 89.375 160.685 89.545 161.595 ;
        RECT 89.715 160.865 89.955 162.175 ;
        RECT 91.045 161.645 92.255 162.735 ;
        RECT 91.045 161.105 91.565 161.645 ;
        RECT 91.735 160.935 92.255 161.475 ;
        RECT 89.375 160.355 89.870 160.685 ;
        RECT 91.045 160.185 92.255 160.935 ;
        RECT 18.280 160.015 92.340 160.185 ;
        RECT 18.365 159.265 19.575 160.015 ;
        RECT 19.745 159.470 25.090 160.015 ;
        RECT 25.265 159.470 30.610 160.015 ;
        RECT 18.365 158.725 18.885 159.265 ;
        RECT 19.055 158.555 19.575 159.095 ;
        RECT 21.330 158.640 21.670 159.470 ;
        RECT 18.365 157.465 19.575 158.555 ;
        RECT 23.150 157.900 23.500 159.150 ;
        RECT 26.850 158.640 27.190 159.470 ;
        RECT 30.785 159.245 33.375 160.015 ;
        RECT 34.030 159.625 34.360 160.015 ;
        RECT 34.530 159.455 34.755 159.835 ;
        RECT 28.670 157.900 29.020 159.150 ;
        RECT 30.785 158.725 31.995 159.245 ;
        RECT 32.165 158.555 33.375 159.075 ;
        RECT 34.015 158.775 34.255 159.425 ;
        RECT 34.425 159.275 34.755 159.455 ;
        RECT 34.425 158.605 34.600 159.275 ;
        RECT 34.955 159.105 35.185 159.725 ;
        RECT 35.365 159.285 35.665 160.015 ;
        RECT 35.845 159.215 36.540 159.845 ;
        RECT 36.745 159.215 37.055 160.015 ;
        RECT 38.145 159.275 38.530 159.845 ;
        RECT 38.700 159.555 39.025 160.015 ;
        RECT 39.545 159.385 39.825 159.845 ;
        RECT 34.770 158.775 35.185 159.105 ;
        RECT 35.365 158.775 35.660 159.105 ;
        RECT 35.865 158.775 36.200 159.025 ;
        RECT 36.370 158.655 36.540 159.215 ;
        RECT 36.710 158.775 37.045 159.045 ;
        RECT 36.365 158.615 36.540 158.655 ;
        RECT 19.745 157.465 25.090 157.900 ;
        RECT 25.265 157.465 30.610 157.900 ;
        RECT 30.785 157.465 33.375 158.555 ;
        RECT 34.015 158.415 34.600 158.605 ;
        RECT 34.015 157.645 34.290 158.415 ;
        RECT 34.770 158.245 35.665 158.575 ;
        RECT 34.460 158.075 35.665 158.245 ;
        RECT 34.460 157.645 34.790 158.075 ;
        RECT 34.960 157.465 35.155 157.905 ;
        RECT 35.335 157.645 35.665 158.075 ;
        RECT 35.845 157.465 36.105 158.605 ;
        RECT 36.275 157.635 36.605 158.615 ;
        RECT 38.145 158.605 38.425 159.275 ;
        RECT 38.700 159.215 39.825 159.385 ;
        RECT 38.700 159.105 39.150 159.215 ;
        RECT 38.595 158.775 39.150 159.105 ;
        RECT 40.015 159.045 40.415 159.845 ;
        RECT 40.815 159.555 41.085 160.015 ;
        RECT 41.255 159.385 41.540 159.845 ;
        RECT 36.775 157.465 37.055 158.605 ;
        RECT 38.145 157.635 38.530 158.605 ;
        RECT 38.700 158.315 39.150 158.775 ;
        RECT 39.320 158.485 40.415 159.045 ;
        RECT 38.700 158.095 39.825 158.315 ;
        RECT 38.700 157.465 39.025 157.925 ;
        RECT 39.545 157.635 39.825 158.095 ;
        RECT 40.015 157.635 40.415 158.485 ;
        RECT 40.585 159.215 41.540 159.385 ;
        RECT 40.585 158.315 40.795 159.215 ;
        RECT 41.835 159.205 42.105 160.015 ;
        RECT 42.275 159.205 42.605 159.845 ;
        RECT 42.775 159.205 43.015 160.015 ;
        RECT 44.125 159.290 44.415 160.015 ;
        RECT 45.530 159.625 45.860 160.015 ;
        RECT 46.030 159.455 46.255 159.835 ;
        RECT 40.965 158.485 41.655 159.045 ;
        RECT 41.825 158.775 42.175 159.025 ;
        RECT 42.345 158.605 42.515 159.205 ;
        RECT 42.685 158.775 43.035 159.025 ;
        RECT 45.515 158.775 45.755 159.425 ;
        RECT 45.925 159.275 46.255 159.455 ;
        RECT 40.585 158.095 41.540 158.315 ;
        RECT 40.815 157.465 41.085 157.925 ;
        RECT 41.255 157.635 41.540 158.095 ;
        RECT 41.835 157.465 42.165 158.605 ;
        RECT 42.345 158.435 43.025 158.605 ;
        RECT 42.695 157.650 43.025 158.435 ;
        RECT 44.125 157.465 44.415 158.630 ;
        RECT 45.925 158.605 46.100 159.275 ;
        RECT 46.455 159.105 46.685 159.725 ;
        RECT 46.865 159.285 47.165 160.015 ;
        RECT 47.345 159.365 47.605 159.845 ;
        RECT 47.775 159.475 48.025 160.015 ;
        RECT 46.270 158.775 46.685 159.105 ;
        RECT 46.865 158.775 47.160 159.105 ;
        RECT 45.515 158.415 46.100 158.605 ;
        RECT 45.515 157.645 45.790 158.415 ;
        RECT 46.270 158.245 47.165 158.575 ;
        RECT 45.960 158.075 47.165 158.245 ;
        RECT 45.960 157.645 46.290 158.075 ;
        RECT 46.460 157.465 46.655 157.905 ;
        RECT 46.835 157.645 47.165 158.075 ;
        RECT 47.345 158.335 47.515 159.365 ;
        RECT 48.195 159.310 48.415 159.795 ;
        RECT 47.685 158.715 47.915 159.110 ;
        RECT 48.085 158.885 48.415 159.310 ;
        RECT 48.585 159.635 49.475 159.805 ;
        RECT 48.585 158.910 48.755 159.635 ;
        RECT 48.925 159.080 49.475 159.465 ;
        RECT 49.760 159.385 50.045 159.845 ;
        RECT 50.215 159.555 50.485 160.015 ;
        RECT 49.760 159.215 50.715 159.385 ;
        RECT 48.585 158.840 49.475 158.910 ;
        RECT 48.580 158.815 49.475 158.840 ;
        RECT 48.570 158.800 49.475 158.815 ;
        RECT 48.565 158.785 49.475 158.800 ;
        RECT 48.555 158.780 49.475 158.785 ;
        RECT 48.550 158.770 49.475 158.780 ;
        RECT 48.545 158.760 49.475 158.770 ;
        RECT 48.535 158.755 49.475 158.760 ;
        RECT 48.525 158.745 49.475 158.755 ;
        RECT 48.515 158.740 49.475 158.745 ;
        RECT 48.515 158.735 48.850 158.740 ;
        RECT 48.500 158.730 48.850 158.735 ;
        RECT 48.485 158.720 48.850 158.730 ;
        RECT 48.460 158.715 48.850 158.720 ;
        RECT 47.685 158.710 48.850 158.715 ;
        RECT 47.685 158.675 48.820 158.710 ;
        RECT 47.685 158.650 48.785 158.675 ;
        RECT 47.685 158.620 48.755 158.650 ;
        RECT 47.685 158.590 48.735 158.620 ;
        RECT 47.685 158.560 48.715 158.590 ;
        RECT 47.685 158.550 48.645 158.560 ;
        RECT 47.685 158.540 48.620 158.550 ;
        RECT 47.685 158.525 48.600 158.540 ;
        RECT 47.685 158.510 48.580 158.525 ;
        RECT 47.790 158.500 48.575 158.510 ;
        RECT 47.790 158.465 48.560 158.500 ;
        RECT 47.345 157.635 47.620 158.335 ;
        RECT 47.790 158.215 48.545 158.465 ;
        RECT 48.715 158.145 49.045 158.390 ;
        RECT 49.215 158.290 49.475 158.740 ;
        RECT 49.645 158.485 50.335 159.045 ;
        RECT 50.505 158.315 50.715 159.215 ;
        RECT 48.860 158.120 49.045 158.145 ;
        RECT 48.860 158.020 49.475 158.120 ;
        RECT 47.790 157.465 48.045 158.010 ;
        RECT 48.215 157.635 48.695 157.975 ;
        RECT 48.870 157.465 49.475 158.020 ;
        RECT 49.760 158.095 50.715 158.315 ;
        RECT 50.885 159.045 51.285 159.845 ;
        RECT 51.475 159.385 51.755 159.845 ;
        RECT 52.275 159.555 52.600 160.015 ;
        RECT 51.475 159.215 52.600 159.385 ;
        RECT 52.770 159.275 53.155 159.845 ;
        RECT 52.150 159.105 52.600 159.215 ;
        RECT 50.885 158.485 51.980 159.045 ;
        RECT 52.150 158.775 52.705 159.105 ;
        RECT 49.760 157.635 50.045 158.095 ;
        RECT 50.215 157.465 50.485 157.925 ;
        RECT 50.885 157.635 51.285 158.485 ;
        RECT 52.150 158.315 52.600 158.775 ;
        RECT 52.875 158.605 53.155 159.275 ;
        RECT 53.335 159.205 53.605 160.015 ;
        RECT 53.775 159.205 54.105 159.845 ;
        RECT 54.275 159.205 54.515 160.015 ;
        RECT 54.705 159.505 55.010 160.015 ;
        RECT 53.325 158.775 53.675 159.025 ;
        RECT 53.845 158.605 54.015 159.205 ;
        RECT 54.185 158.775 54.535 159.025 ;
        RECT 54.705 158.775 55.020 159.335 ;
        RECT 55.190 159.025 55.440 159.835 ;
        RECT 55.610 159.490 55.870 160.015 ;
        RECT 56.050 159.025 56.300 159.835 ;
        RECT 56.470 159.455 56.730 160.015 ;
        RECT 56.900 159.365 57.160 159.820 ;
        RECT 57.330 159.535 57.590 160.015 ;
        RECT 57.760 159.365 58.020 159.820 ;
        RECT 58.190 159.535 58.450 160.015 ;
        RECT 58.620 159.365 58.880 159.820 ;
        RECT 59.050 159.535 59.295 160.015 ;
        RECT 59.465 159.365 59.740 159.820 ;
        RECT 59.910 159.535 60.155 160.015 ;
        RECT 60.325 159.365 60.585 159.820 ;
        RECT 60.765 159.535 61.015 160.015 ;
        RECT 61.185 159.365 61.445 159.820 ;
        RECT 61.625 159.535 61.875 160.015 ;
        RECT 62.045 159.365 62.305 159.820 ;
        RECT 62.485 159.535 62.745 160.015 ;
        RECT 62.915 159.365 63.175 159.820 ;
        RECT 63.345 159.535 63.645 160.015 ;
        RECT 56.900 159.195 63.645 159.365 ;
        RECT 55.190 158.775 62.310 159.025 ;
        RECT 51.475 158.095 52.600 158.315 ;
        RECT 51.475 157.635 51.755 158.095 ;
        RECT 52.275 157.465 52.600 157.925 ;
        RECT 52.770 157.635 53.155 158.605 ;
        RECT 53.335 157.465 53.665 158.605 ;
        RECT 53.845 158.435 54.525 158.605 ;
        RECT 54.195 157.650 54.525 158.435 ;
        RECT 54.715 157.465 55.010 158.275 ;
        RECT 55.190 157.635 55.435 158.775 ;
        RECT 55.610 157.465 55.870 158.275 ;
        RECT 56.050 157.640 56.300 158.775 ;
        RECT 62.480 158.605 63.645 159.195 ;
        RECT 63.905 159.245 65.575 160.015 ;
        RECT 65.745 159.275 66.130 159.845 ;
        RECT 66.300 159.555 66.625 160.015 ;
        RECT 67.145 159.385 67.425 159.845 ;
        RECT 63.905 158.725 64.655 159.245 ;
        RECT 56.900 158.380 63.645 158.605 ;
        RECT 64.825 158.555 65.575 159.075 ;
        RECT 56.900 158.365 62.305 158.380 ;
        RECT 56.470 157.470 56.730 158.265 ;
        RECT 56.900 157.640 57.160 158.365 ;
        RECT 57.330 157.470 57.590 158.195 ;
        RECT 57.760 157.640 58.020 158.365 ;
        RECT 58.190 157.470 58.450 158.195 ;
        RECT 58.620 157.640 58.880 158.365 ;
        RECT 59.050 157.470 59.310 158.195 ;
        RECT 59.480 157.640 59.740 158.365 ;
        RECT 59.910 157.470 60.155 158.195 ;
        RECT 60.325 157.640 60.585 158.365 ;
        RECT 60.770 157.470 61.015 158.195 ;
        RECT 61.185 157.640 61.445 158.365 ;
        RECT 61.630 157.470 61.875 158.195 ;
        RECT 62.045 157.640 62.305 158.365 ;
        RECT 62.490 157.470 62.745 158.195 ;
        RECT 62.915 157.640 63.205 158.380 ;
        RECT 56.470 157.465 62.745 157.470 ;
        RECT 63.375 157.465 63.645 158.210 ;
        RECT 63.905 157.465 65.575 158.555 ;
        RECT 65.745 158.605 66.025 159.275 ;
        RECT 66.300 159.215 67.425 159.385 ;
        RECT 66.300 159.105 66.750 159.215 ;
        RECT 66.195 158.775 66.750 159.105 ;
        RECT 67.615 159.045 68.015 159.845 ;
        RECT 68.415 159.555 68.685 160.015 ;
        RECT 68.855 159.385 69.140 159.845 ;
        RECT 65.745 157.635 66.130 158.605 ;
        RECT 66.300 158.315 66.750 158.775 ;
        RECT 66.920 158.485 68.015 159.045 ;
        RECT 66.300 158.095 67.425 158.315 ;
        RECT 66.300 157.465 66.625 157.925 ;
        RECT 67.145 157.635 67.425 158.095 ;
        RECT 67.615 157.635 68.015 158.485 ;
        RECT 68.185 159.215 69.140 159.385 ;
        RECT 69.885 159.290 70.175 160.015 ;
        RECT 70.345 159.265 71.555 160.015 ;
        RECT 71.735 159.285 72.035 160.015 ;
        RECT 68.185 158.315 68.395 159.215 ;
        RECT 68.565 158.485 69.255 159.045 ;
        RECT 70.345 158.725 70.865 159.265 ;
        RECT 72.215 159.105 72.445 159.725 ;
        RECT 72.645 159.455 72.870 159.835 ;
        RECT 73.040 159.625 73.370 160.015 ;
        RECT 72.645 159.275 72.975 159.455 ;
        RECT 68.185 158.095 69.140 158.315 ;
        RECT 68.415 157.465 68.685 157.925 ;
        RECT 68.855 157.635 69.140 158.095 ;
        RECT 69.885 157.465 70.175 158.630 ;
        RECT 71.035 158.555 71.555 159.095 ;
        RECT 71.740 158.775 72.035 159.105 ;
        RECT 72.215 158.775 72.630 159.105 ;
        RECT 72.800 158.605 72.975 159.275 ;
        RECT 73.145 158.775 73.385 159.425 ;
        RECT 73.565 159.245 75.235 160.015 ;
        RECT 75.405 159.515 75.705 159.845 ;
        RECT 75.875 159.535 76.150 160.015 ;
        RECT 73.565 158.725 74.315 159.245 ;
        RECT 70.345 157.465 71.555 158.555 ;
        RECT 71.735 158.245 72.630 158.575 ;
        RECT 72.800 158.415 73.385 158.605 ;
        RECT 74.485 158.555 75.235 159.075 ;
        RECT 71.735 158.075 72.940 158.245 ;
        RECT 71.735 157.645 72.065 158.075 ;
        RECT 72.245 157.465 72.440 157.905 ;
        RECT 72.610 157.645 72.940 158.075 ;
        RECT 73.110 157.645 73.385 158.415 ;
        RECT 73.565 157.465 75.235 158.555 ;
        RECT 75.405 158.605 75.575 159.515 ;
        RECT 76.330 159.365 76.625 159.755 ;
        RECT 76.795 159.535 77.050 160.015 ;
        RECT 77.225 159.365 77.485 159.755 ;
        RECT 77.655 159.535 77.935 160.015 ;
        RECT 75.745 158.775 76.095 159.345 ;
        RECT 76.330 159.195 77.980 159.365 ;
        RECT 76.265 158.855 77.405 159.025 ;
        RECT 76.265 158.605 76.435 158.855 ;
        RECT 77.575 158.685 77.980 159.195 ;
        RECT 78.165 159.265 79.375 160.015 ;
        RECT 79.635 159.465 79.805 159.755 ;
        RECT 79.975 159.635 80.305 160.015 ;
        RECT 79.635 159.295 80.300 159.465 ;
        RECT 78.165 158.725 78.685 159.265 ;
        RECT 75.405 158.435 76.435 158.605 ;
        RECT 77.225 158.515 77.980 158.685 ;
        RECT 78.855 158.555 79.375 159.095 ;
        RECT 75.405 157.635 75.715 158.435 ;
        RECT 77.225 158.265 77.485 158.515 ;
        RECT 75.885 157.465 76.195 158.265 ;
        RECT 76.365 158.095 77.485 158.265 ;
        RECT 76.365 157.635 76.625 158.095 ;
        RECT 76.795 157.465 77.050 157.925 ;
        RECT 77.225 157.635 77.485 158.095 ;
        RECT 77.655 157.465 77.940 158.335 ;
        RECT 78.165 157.465 79.375 158.555 ;
        RECT 79.550 158.475 79.900 159.125 ;
        RECT 80.070 158.305 80.300 159.295 ;
        RECT 79.635 158.135 80.300 158.305 ;
        RECT 79.635 157.635 79.805 158.135 ;
        RECT 79.975 157.465 80.305 157.965 ;
        RECT 80.475 157.635 80.700 159.755 ;
        RECT 80.915 159.555 81.165 160.015 ;
        RECT 81.350 159.565 81.680 159.735 ;
        RECT 81.860 159.565 82.610 159.735 ;
        RECT 80.900 158.435 81.180 159.035 ;
        RECT 81.350 158.035 81.520 159.565 ;
        RECT 81.690 159.065 82.270 159.395 ;
        RECT 81.690 158.195 81.930 159.065 ;
        RECT 82.440 158.785 82.610 159.565 ;
        RECT 82.860 159.515 83.230 160.015 ;
        RECT 83.410 159.565 83.870 159.735 ;
        RECT 84.100 159.565 84.770 159.735 ;
        RECT 83.410 159.335 83.580 159.565 ;
        RECT 82.780 159.035 83.580 159.335 ;
        RECT 83.750 159.065 84.300 159.395 ;
        RECT 82.780 159.005 82.950 159.035 ;
        RECT 83.070 158.785 83.240 158.855 ;
        RECT 82.440 158.615 83.240 158.785 ;
        RECT 82.730 158.525 83.240 158.615 ;
        RECT 82.120 158.090 82.560 158.445 ;
        RECT 80.900 157.465 81.165 157.925 ;
        RECT 81.350 157.660 81.585 158.035 ;
        RECT 82.730 157.910 82.900 158.525 ;
        RECT 81.830 157.740 82.900 157.910 ;
        RECT 83.070 157.465 83.240 158.265 ;
        RECT 83.410 157.965 83.580 159.035 ;
        RECT 83.750 158.135 83.940 158.855 ;
        RECT 84.110 158.525 84.300 159.065 ;
        RECT 84.600 159.025 84.770 159.565 ;
        RECT 85.085 159.485 85.255 160.015 ;
        RECT 85.550 159.365 85.910 159.805 ;
        RECT 86.085 159.535 86.255 160.015 ;
        RECT 86.445 159.370 86.780 159.795 ;
        RECT 86.955 159.540 87.125 160.015 ;
        RECT 87.300 159.370 87.635 159.795 ;
        RECT 87.805 159.540 87.975 160.015 ;
        RECT 85.550 159.195 86.050 159.365 ;
        RECT 86.445 159.200 88.115 159.370 ;
        RECT 85.880 159.025 86.050 159.195 ;
        RECT 84.600 158.855 85.690 159.025 ;
        RECT 85.880 158.855 87.700 159.025 ;
        RECT 84.110 158.195 84.430 158.525 ;
        RECT 83.410 157.635 83.660 157.965 ;
        RECT 84.600 157.935 84.770 158.855 ;
        RECT 85.880 158.600 86.050 158.855 ;
        RECT 87.870 158.635 88.115 159.200 ;
        RECT 88.285 159.245 90.875 160.015 ;
        RECT 91.045 159.265 92.255 160.015 ;
        RECT 88.285 158.725 89.495 159.245 ;
        RECT 84.940 158.430 86.050 158.600 ;
        RECT 86.445 158.465 88.115 158.635 ;
        RECT 89.665 158.555 90.875 159.075 ;
        RECT 84.940 158.270 85.800 158.430 ;
        RECT 83.885 157.765 84.770 157.935 ;
        RECT 84.950 157.465 85.165 157.965 ;
        RECT 85.630 157.645 85.800 158.270 ;
        RECT 86.085 157.465 86.265 158.245 ;
        RECT 86.445 157.705 86.780 158.465 ;
        RECT 86.960 157.465 87.130 158.295 ;
        RECT 87.300 157.705 87.630 158.465 ;
        RECT 87.800 157.465 87.970 158.295 ;
        RECT 88.285 157.465 90.875 158.555 ;
        RECT 91.045 158.555 91.565 159.095 ;
        RECT 91.735 158.725 92.255 159.265 ;
        RECT 91.045 157.465 92.255 158.555 ;
        RECT 18.280 157.295 92.340 157.465 ;
        RECT 18.365 156.205 19.575 157.295 ;
        RECT 19.745 156.860 25.090 157.295 ;
        RECT 25.265 156.860 30.610 157.295 ;
        RECT 18.365 155.495 18.885 156.035 ;
        RECT 19.055 155.665 19.575 156.205 ;
        RECT 18.365 154.745 19.575 155.495 ;
        RECT 21.330 155.290 21.670 156.120 ;
        RECT 23.150 155.610 23.500 156.860 ;
        RECT 26.850 155.290 27.190 156.120 ;
        RECT 28.670 155.610 29.020 156.860 ;
        RECT 31.245 156.130 31.535 157.295 ;
        RECT 32.255 156.625 32.425 157.125 ;
        RECT 32.595 156.795 32.925 157.295 ;
        RECT 32.255 156.455 32.920 156.625 ;
        RECT 32.170 155.635 32.520 156.285 ;
        RECT 19.745 154.745 25.090 155.290 ;
        RECT 25.265 154.745 30.610 155.290 ;
        RECT 31.245 154.745 31.535 155.470 ;
        RECT 32.690 155.465 32.920 156.455 ;
        RECT 32.255 155.295 32.920 155.465 ;
        RECT 32.255 155.005 32.425 155.295 ;
        RECT 32.595 154.745 32.925 155.125 ;
        RECT 33.095 155.005 33.280 157.125 ;
        RECT 33.520 156.835 33.785 157.295 ;
        RECT 33.955 156.700 34.205 157.125 ;
        RECT 34.415 156.850 35.520 157.020 ;
        RECT 33.900 156.570 34.205 156.700 ;
        RECT 33.450 155.375 33.730 156.325 ;
        RECT 33.900 155.465 34.070 156.570 ;
        RECT 34.240 155.785 34.480 156.380 ;
        RECT 34.650 156.315 35.180 156.680 ;
        RECT 34.650 155.615 34.820 156.315 ;
        RECT 35.350 156.235 35.520 156.850 ;
        RECT 35.690 156.495 35.860 157.295 ;
        RECT 36.030 156.795 36.280 157.125 ;
        RECT 36.505 156.825 37.390 156.995 ;
        RECT 35.350 156.145 35.860 156.235 ;
        RECT 33.900 155.335 34.125 155.465 ;
        RECT 34.295 155.395 34.820 155.615 ;
        RECT 34.990 155.975 35.860 156.145 ;
        RECT 33.535 154.745 33.785 155.205 ;
        RECT 33.955 155.195 34.125 155.335 ;
        RECT 34.990 155.195 35.160 155.975 ;
        RECT 35.690 155.905 35.860 155.975 ;
        RECT 35.370 155.725 35.570 155.755 ;
        RECT 36.030 155.725 36.200 156.795 ;
        RECT 36.370 155.905 36.560 156.625 ;
        RECT 35.370 155.425 36.200 155.725 ;
        RECT 36.730 155.695 37.050 156.655 ;
        RECT 33.955 155.025 34.290 155.195 ;
        RECT 34.485 155.025 35.160 155.195 ;
        RECT 35.480 154.745 35.850 155.245 ;
        RECT 36.030 155.195 36.200 155.425 ;
        RECT 36.585 155.365 37.050 155.695 ;
        RECT 37.220 155.985 37.390 156.825 ;
        RECT 37.570 156.795 37.885 157.295 ;
        RECT 38.115 156.565 38.455 157.125 ;
        RECT 37.560 156.190 38.455 156.565 ;
        RECT 38.625 156.285 38.795 157.295 ;
        RECT 38.265 155.985 38.455 156.190 ;
        RECT 38.965 156.235 39.295 157.080 ;
        RECT 40.535 156.625 40.705 157.125 ;
        RECT 40.875 156.795 41.205 157.295 ;
        RECT 40.535 156.455 41.200 156.625 ;
        RECT 38.965 156.155 39.355 156.235 ;
        RECT 39.140 156.105 39.355 156.155 ;
        RECT 37.220 155.655 38.095 155.985 ;
        RECT 38.265 155.655 39.015 155.985 ;
        RECT 37.220 155.195 37.390 155.655 ;
        RECT 38.265 155.485 38.465 155.655 ;
        RECT 39.185 155.525 39.355 156.105 ;
        RECT 40.450 155.635 40.800 156.285 ;
        RECT 39.130 155.485 39.355 155.525 ;
        RECT 36.030 155.025 36.435 155.195 ;
        RECT 36.605 155.025 37.390 155.195 ;
        RECT 37.665 154.745 37.875 155.275 ;
        RECT 38.135 154.960 38.465 155.485 ;
        RECT 38.975 155.400 39.355 155.485 ;
        RECT 40.970 155.465 41.200 156.455 ;
        RECT 38.635 154.745 38.805 155.355 ;
        RECT 38.975 154.965 39.305 155.400 ;
        RECT 40.535 155.295 41.200 155.465 ;
        RECT 40.535 155.005 40.705 155.295 ;
        RECT 40.875 154.745 41.205 155.125 ;
        RECT 41.375 155.005 41.560 157.125 ;
        RECT 41.800 156.835 42.065 157.295 ;
        RECT 42.235 156.700 42.485 157.125 ;
        RECT 42.695 156.850 43.800 157.020 ;
        RECT 42.180 156.570 42.485 156.700 ;
        RECT 41.730 155.375 42.010 156.325 ;
        RECT 42.180 155.465 42.350 156.570 ;
        RECT 42.520 155.785 42.760 156.380 ;
        RECT 42.930 156.315 43.460 156.680 ;
        RECT 42.930 155.615 43.100 156.315 ;
        RECT 43.630 156.235 43.800 156.850 ;
        RECT 43.970 156.495 44.140 157.295 ;
        RECT 44.310 156.795 44.560 157.125 ;
        RECT 44.785 156.825 45.670 156.995 ;
        RECT 43.630 156.145 44.140 156.235 ;
        RECT 42.180 155.335 42.405 155.465 ;
        RECT 42.575 155.395 43.100 155.615 ;
        RECT 43.270 155.975 44.140 156.145 ;
        RECT 41.815 154.745 42.065 155.205 ;
        RECT 42.235 155.195 42.405 155.335 ;
        RECT 43.270 155.195 43.440 155.975 ;
        RECT 43.970 155.905 44.140 155.975 ;
        RECT 43.650 155.725 43.850 155.755 ;
        RECT 44.310 155.725 44.480 156.795 ;
        RECT 44.650 155.905 44.840 156.625 ;
        RECT 43.650 155.425 44.480 155.725 ;
        RECT 45.010 155.695 45.330 156.655 ;
        RECT 42.235 155.025 42.570 155.195 ;
        RECT 42.765 155.025 43.440 155.195 ;
        RECT 43.760 154.745 44.130 155.245 ;
        RECT 44.310 155.195 44.480 155.425 ;
        RECT 44.865 155.365 45.330 155.695 ;
        RECT 45.500 155.985 45.670 156.825 ;
        RECT 45.850 156.795 46.165 157.295 ;
        RECT 46.395 156.565 46.735 157.125 ;
        RECT 45.840 156.190 46.735 156.565 ;
        RECT 46.905 156.285 47.075 157.295 ;
        RECT 46.545 155.985 46.735 156.190 ;
        RECT 47.245 156.235 47.575 157.080 ;
        RECT 47.245 156.155 47.635 156.235 ;
        RECT 47.805 156.205 49.475 157.295 ;
        RECT 49.705 156.235 50.035 157.080 ;
        RECT 50.205 156.285 50.375 157.295 ;
        RECT 50.545 156.565 50.885 157.125 ;
        RECT 51.115 156.795 51.430 157.295 ;
        RECT 51.610 156.825 52.495 156.995 ;
        RECT 47.420 156.105 47.635 156.155 ;
        RECT 45.500 155.655 46.375 155.985 ;
        RECT 46.545 155.655 47.295 155.985 ;
        RECT 45.500 155.195 45.670 155.655 ;
        RECT 46.545 155.485 46.745 155.655 ;
        RECT 47.465 155.525 47.635 156.105 ;
        RECT 47.410 155.485 47.635 155.525 ;
        RECT 44.310 155.025 44.715 155.195 ;
        RECT 44.885 155.025 45.670 155.195 ;
        RECT 45.945 154.745 46.155 155.275 ;
        RECT 46.415 154.960 46.745 155.485 ;
        RECT 47.255 155.400 47.635 155.485 ;
        RECT 47.805 155.515 48.555 156.035 ;
        RECT 48.725 155.685 49.475 156.205 ;
        RECT 49.645 156.155 50.035 156.235 ;
        RECT 50.545 156.190 51.440 156.565 ;
        RECT 49.645 156.105 49.860 156.155 ;
        RECT 49.645 155.525 49.815 156.105 ;
        RECT 50.545 155.985 50.735 156.190 ;
        RECT 51.610 155.985 51.780 156.825 ;
        RECT 52.720 156.795 52.970 157.125 ;
        RECT 49.985 155.655 50.735 155.985 ;
        RECT 50.905 155.655 51.780 155.985 ;
        RECT 46.915 154.745 47.085 155.355 ;
        RECT 47.255 154.965 47.585 155.400 ;
        RECT 47.805 154.745 49.475 155.515 ;
        RECT 49.645 155.485 49.870 155.525 ;
        RECT 50.535 155.485 50.735 155.655 ;
        RECT 49.645 155.400 50.025 155.485 ;
        RECT 49.695 154.965 50.025 155.400 ;
        RECT 50.195 154.745 50.365 155.355 ;
        RECT 50.535 154.960 50.865 155.485 ;
        RECT 51.125 154.745 51.335 155.275 ;
        RECT 51.610 155.195 51.780 155.655 ;
        RECT 51.950 155.695 52.270 156.655 ;
        RECT 52.440 155.905 52.630 156.625 ;
        RECT 52.800 155.725 52.970 156.795 ;
        RECT 53.140 156.495 53.310 157.295 ;
        RECT 53.480 156.850 54.585 157.020 ;
        RECT 53.480 156.235 53.650 156.850 ;
        RECT 54.795 156.700 55.045 157.125 ;
        RECT 55.215 156.835 55.480 157.295 ;
        RECT 53.820 156.315 54.350 156.680 ;
        RECT 54.795 156.570 55.100 156.700 ;
        RECT 53.140 156.145 53.650 156.235 ;
        RECT 53.140 155.975 54.010 156.145 ;
        RECT 53.140 155.905 53.310 155.975 ;
        RECT 53.430 155.725 53.630 155.755 ;
        RECT 51.950 155.365 52.415 155.695 ;
        RECT 52.800 155.425 53.630 155.725 ;
        RECT 52.800 155.195 52.970 155.425 ;
        RECT 51.610 155.025 52.395 155.195 ;
        RECT 52.565 155.025 52.970 155.195 ;
        RECT 53.150 154.745 53.520 155.245 ;
        RECT 53.840 155.195 54.010 155.975 ;
        RECT 54.180 155.615 54.350 156.315 ;
        RECT 54.520 155.785 54.760 156.380 ;
        RECT 54.180 155.395 54.705 155.615 ;
        RECT 54.930 155.465 55.100 156.570 ;
        RECT 54.875 155.335 55.100 155.465 ;
        RECT 55.270 155.375 55.550 156.325 ;
        RECT 54.875 155.195 55.045 155.335 ;
        RECT 53.840 155.025 54.515 155.195 ;
        RECT 54.710 155.025 55.045 155.195 ;
        RECT 55.215 154.745 55.465 155.205 ;
        RECT 55.720 155.005 55.905 157.125 ;
        RECT 56.075 156.795 56.405 157.295 ;
        RECT 56.575 156.625 56.745 157.125 ;
        RECT 56.080 156.455 56.745 156.625 ;
        RECT 56.080 155.465 56.310 156.455 ;
        RECT 56.480 155.635 56.830 156.285 ;
        RECT 57.005 156.130 57.295 157.295 ;
        RECT 57.465 156.205 60.055 157.295 ;
        RECT 60.315 156.625 60.485 157.125 ;
        RECT 60.655 156.795 60.985 157.295 ;
        RECT 60.315 156.455 60.980 156.625 ;
        RECT 57.465 155.515 58.675 156.035 ;
        RECT 58.845 155.685 60.055 156.205 ;
        RECT 60.230 155.635 60.580 156.285 ;
        RECT 56.080 155.295 56.745 155.465 ;
        RECT 56.075 154.745 56.405 155.125 ;
        RECT 56.575 155.005 56.745 155.295 ;
        RECT 57.005 154.745 57.295 155.470 ;
        RECT 57.465 154.745 60.055 155.515 ;
        RECT 60.750 155.465 60.980 156.455 ;
        RECT 60.315 155.295 60.980 155.465 ;
        RECT 60.315 155.005 60.485 155.295 ;
        RECT 60.655 154.745 60.985 155.125 ;
        RECT 61.155 155.005 61.340 157.125 ;
        RECT 61.580 156.835 61.845 157.295 ;
        RECT 62.015 156.700 62.265 157.125 ;
        RECT 62.475 156.850 63.580 157.020 ;
        RECT 61.960 156.570 62.265 156.700 ;
        RECT 61.510 155.375 61.790 156.325 ;
        RECT 61.960 155.465 62.130 156.570 ;
        RECT 62.300 155.785 62.540 156.380 ;
        RECT 62.710 156.315 63.240 156.680 ;
        RECT 62.710 155.615 62.880 156.315 ;
        RECT 63.410 156.235 63.580 156.850 ;
        RECT 63.750 156.495 63.920 157.295 ;
        RECT 64.090 156.795 64.340 157.125 ;
        RECT 64.565 156.825 65.450 156.995 ;
        RECT 63.410 156.145 63.920 156.235 ;
        RECT 61.960 155.335 62.185 155.465 ;
        RECT 62.355 155.395 62.880 155.615 ;
        RECT 63.050 155.975 63.920 156.145 ;
        RECT 61.595 154.745 61.845 155.205 ;
        RECT 62.015 155.195 62.185 155.335 ;
        RECT 63.050 155.195 63.220 155.975 ;
        RECT 63.750 155.905 63.920 155.975 ;
        RECT 63.430 155.725 63.630 155.755 ;
        RECT 64.090 155.725 64.260 156.795 ;
        RECT 64.430 155.905 64.620 156.625 ;
        RECT 63.430 155.425 64.260 155.725 ;
        RECT 64.790 155.695 65.110 156.655 ;
        RECT 62.015 155.025 62.350 155.195 ;
        RECT 62.545 155.025 63.220 155.195 ;
        RECT 63.540 154.745 63.910 155.245 ;
        RECT 64.090 155.195 64.260 155.425 ;
        RECT 64.645 155.365 65.110 155.695 ;
        RECT 65.280 155.985 65.450 156.825 ;
        RECT 65.630 156.795 65.945 157.295 ;
        RECT 66.175 156.565 66.515 157.125 ;
        RECT 65.620 156.190 66.515 156.565 ;
        RECT 66.685 156.285 66.855 157.295 ;
        RECT 66.325 155.985 66.515 156.190 ;
        RECT 67.025 156.235 67.355 157.080 ;
        RECT 67.025 156.155 67.415 156.235 ;
        RECT 67.585 156.205 71.095 157.295 ;
        RECT 72.275 156.625 72.445 157.125 ;
        RECT 72.615 156.795 72.945 157.295 ;
        RECT 72.275 156.455 72.940 156.625 ;
        RECT 67.200 156.105 67.415 156.155 ;
        RECT 65.280 155.655 66.155 155.985 ;
        RECT 66.325 155.655 67.075 155.985 ;
        RECT 65.280 155.195 65.450 155.655 ;
        RECT 66.325 155.485 66.525 155.655 ;
        RECT 67.245 155.525 67.415 156.105 ;
        RECT 67.190 155.485 67.415 155.525 ;
        RECT 64.090 155.025 64.495 155.195 ;
        RECT 64.665 155.025 65.450 155.195 ;
        RECT 65.725 154.745 65.935 155.275 ;
        RECT 66.195 154.960 66.525 155.485 ;
        RECT 67.035 155.400 67.415 155.485 ;
        RECT 67.585 155.515 69.235 156.035 ;
        RECT 69.405 155.685 71.095 156.205 ;
        RECT 72.190 155.635 72.540 156.285 ;
        RECT 66.695 154.745 66.865 155.355 ;
        RECT 67.035 154.965 67.365 155.400 ;
        RECT 67.585 154.745 71.095 155.515 ;
        RECT 72.710 155.465 72.940 156.455 ;
        RECT 72.275 155.295 72.940 155.465 ;
        RECT 72.275 155.005 72.445 155.295 ;
        RECT 72.615 154.745 72.945 155.125 ;
        RECT 73.115 155.005 73.340 157.125 ;
        RECT 73.540 156.835 73.805 157.295 ;
        RECT 73.990 156.725 74.225 157.100 ;
        RECT 74.470 156.850 75.540 157.020 ;
        RECT 73.540 155.725 73.820 156.325 ;
        RECT 73.555 154.745 73.805 155.205 ;
        RECT 73.990 155.195 74.160 156.725 ;
        RECT 74.330 155.695 74.570 156.565 ;
        RECT 74.760 156.315 75.200 156.670 ;
        RECT 75.370 156.235 75.540 156.850 ;
        RECT 75.710 156.495 75.880 157.295 ;
        RECT 76.050 156.795 76.300 157.125 ;
        RECT 76.525 156.825 77.410 156.995 ;
        RECT 75.370 156.145 75.880 156.235 ;
        RECT 75.080 155.975 75.880 156.145 ;
        RECT 74.330 155.365 74.910 155.695 ;
        RECT 75.080 155.195 75.250 155.975 ;
        RECT 75.710 155.905 75.880 155.975 ;
        RECT 75.420 155.725 75.590 155.755 ;
        RECT 76.050 155.725 76.220 156.795 ;
        RECT 76.390 155.905 76.580 156.625 ;
        RECT 76.750 156.235 77.070 156.565 ;
        RECT 75.420 155.425 76.220 155.725 ;
        RECT 76.750 155.695 76.940 156.235 ;
        RECT 73.990 155.025 74.320 155.195 ;
        RECT 74.500 155.025 75.250 155.195 ;
        RECT 75.500 154.745 75.870 155.245 ;
        RECT 76.050 155.195 76.220 155.425 ;
        RECT 76.390 155.365 76.940 155.695 ;
        RECT 77.240 155.905 77.410 156.825 ;
        RECT 77.590 156.795 77.805 157.295 ;
        RECT 78.270 156.490 78.440 157.115 ;
        RECT 78.725 156.515 78.905 157.295 ;
        RECT 77.580 156.330 78.440 156.490 ;
        RECT 77.580 156.160 78.690 156.330 ;
        RECT 78.520 155.905 78.690 156.160 ;
        RECT 79.085 156.295 79.420 157.055 ;
        RECT 79.600 156.465 79.770 157.295 ;
        RECT 79.940 156.295 80.270 157.055 ;
        RECT 80.440 156.465 80.610 157.295 ;
        RECT 79.085 156.125 80.755 156.295 ;
        RECT 80.925 156.205 82.595 157.295 ;
        RECT 77.240 155.735 78.330 155.905 ;
        RECT 78.520 155.735 80.340 155.905 ;
        RECT 77.240 155.195 77.410 155.735 ;
        RECT 78.520 155.565 78.690 155.735 ;
        RECT 78.190 155.395 78.690 155.565 ;
        RECT 80.510 155.560 80.755 156.125 ;
        RECT 76.050 155.025 76.510 155.195 ;
        RECT 76.740 155.025 77.410 155.195 ;
        RECT 77.725 154.745 77.895 155.275 ;
        RECT 78.190 154.955 78.550 155.395 ;
        RECT 79.085 155.390 80.755 155.560 ;
        RECT 80.925 155.515 81.675 156.035 ;
        RECT 81.845 155.685 82.595 156.205 ;
        RECT 82.765 156.130 83.055 157.295 ;
        RECT 83.225 156.860 88.570 157.295 ;
        RECT 78.725 154.745 78.895 155.225 ;
        RECT 79.085 154.965 79.420 155.390 ;
        RECT 79.595 154.745 79.765 155.220 ;
        RECT 79.940 154.965 80.275 155.390 ;
        RECT 80.445 154.745 80.615 155.220 ;
        RECT 80.925 154.745 82.595 155.515 ;
        RECT 82.765 154.745 83.055 155.470 ;
        RECT 84.810 155.290 85.150 156.120 ;
        RECT 86.630 155.610 86.980 156.860 ;
        RECT 88.745 156.205 90.415 157.295 ;
        RECT 88.745 155.515 89.495 156.035 ;
        RECT 89.665 155.685 90.415 156.205 ;
        RECT 91.045 156.205 92.255 157.295 ;
        RECT 91.045 155.665 91.565 156.205 ;
        RECT 83.225 154.745 88.570 155.290 ;
        RECT 88.745 154.745 90.415 155.515 ;
        RECT 91.735 155.495 92.255 156.035 ;
        RECT 91.045 154.745 92.255 155.495 ;
        RECT 18.280 154.575 92.340 154.745 ;
        RECT 18.365 153.825 19.575 154.575 ;
        RECT 19.745 154.030 25.090 154.575 ;
        RECT 25.265 154.030 30.610 154.575 ;
        RECT 30.785 154.030 36.130 154.575 ;
        RECT 36.305 154.030 41.650 154.575 ;
        RECT 18.365 153.285 18.885 153.825 ;
        RECT 19.055 153.115 19.575 153.655 ;
        RECT 21.330 153.200 21.670 154.030 ;
        RECT 18.365 152.025 19.575 153.115 ;
        RECT 23.150 152.460 23.500 153.710 ;
        RECT 26.850 153.200 27.190 154.030 ;
        RECT 28.670 152.460 29.020 153.710 ;
        RECT 32.370 153.200 32.710 154.030 ;
        RECT 34.190 152.460 34.540 153.710 ;
        RECT 37.890 153.200 38.230 154.030 ;
        RECT 41.825 153.805 43.495 154.575 ;
        RECT 44.125 153.850 44.415 154.575 ;
        RECT 44.585 154.030 49.930 154.575 ;
        RECT 50.105 154.030 55.450 154.575 ;
        RECT 55.625 154.030 60.970 154.575 ;
        RECT 61.145 154.030 66.490 154.575 ;
        RECT 39.710 152.460 40.060 153.710 ;
        RECT 41.825 153.285 42.575 153.805 ;
        RECT 42.745 153.115 43.495 153.635 ;
        RECT 46.170 153.200 46.510 154.030 ;
        RECT 19.745 152.025 25.090 152.460 ;
        RECT 25.265 152.025 30.610 152.460 ;
        RECT 30.785 152.025 36.130 152.460 ;
        RECT 36.305 152.025 41.650 152.460 ;
        RECT 41.825 152.025 43.495 153.115 ;
        RECT 44.125 152.025 44.415 153.190 ;
        RECT 47.990 152.460 48.340 153.710 ;
        RECT 51.690 153.200 52.030 154.030 ;
        RECT 53.510 152.460 53.860 153.710 ;
        RECT 57.210 153.200 57.550 154.030 ;
        RECT 59.030 152.460 59.380 153.710 ;
        RECT 62.730 153.200 63.070 154.030 ;
        RECT 66.665 153.805 69.255 154.575 ;
        RECT 69.885 153.850 70.175 154.575 ;
        RECT 70.345 154.030 75.690 154.575 ;
        RECT 75.865 154.030 81.210 154.575 ;
        RECT 81.385 154.030 86.730 154.575 ;
        RECT 64.550 152.460 64.900 153.710 ;
        RECT 66.665 153.285 67.875 153.805 ;
        RECT 68.045 153.115 69.255 153.635 ;
        RECT 71.930 153.200 72.270 154.030 ;
        RECT 44.585 152.025 49.930 152.460 ;
        RECT 50.105 152.025 55.450 152.460 ;
        RECT 55.625 152.025 60.970 152.460 ;
        RECT 61.145 152.025 66.490 152.460 ;
        RECT 66.665 152.025 69.255 153.115 ;
        RECT 69.885 152.025 70.175 153.190 ;
        RECT 73.750 152.460 74.100 153.710 ;
        RECT 77.450 153.200 77.790 154.030 ;
        RECT 79.270 152.460 79.620 153.710 ;
        RECT 82.970 153.200 83.310 154.030 ;
        RECT 86.905 153.805 90.415 154.575 ;
        RECT 91.045 153.825 92.255 154.575 ;
        RECT 84.790 152.460 85.140 153.710 ;
        RECT 86.905 153.285 88.555 153.805 ;
        RECT 88.725 153.115 90.415 153.635 ;
        RECT 70.345 152.025 75.690 152.460 ;
        RECT 75.865 152.025 81.210 152.460 ;
        RECT 81.385 152.025 86.730 152.460 ;
        RECT 86.905 152.025 90.415 153.115 ;
        RECT 91.045 153.115 91.565 153.655 ;
        RECT 91.735 153.285 92.255 153.825 ;
        RECT 91.045 152.025 92.255 153.115 ;
        RECT 18.280 151.855 92.340 152.025 ;
        RECT 18.365 150.765 19.575 151.855 ;
        RECT 19.745 151.420 25.090 151.855 ;
        RECT 25.265 151.420 30.610 151.855 ;
        RECT 18.365 150.055 18.885 150.595 ;
        RECT 19.055 150.225 19.575 150.765 ;
        RECT 18.365 149.305 19.575 150.055 ;
        RECT 21.330 149.850 21.670 150.680 ;
        RECT 23.150 150.170 23.500 151.420 ;
        RECT 26.850 149.850 27.190 150.680 ;
        RECT 28.670 150.170 29.020 151.420 ;
        RECT 31.245 150.690 31.535 151.855 ;
        RECT 31.705 151.420 37.050 151.855 ;
        RECT 37.225 151.420 42.570 151.855 ;
        RECT 42.745 151.420 48.090 151.855 ;
        RECT 48.265 151.420 53.610 151.855 ;
        RECT 19.745 149.305 25.090 149.850 ;
        RECT 25.265 149.305 30.610 149.850 ;
        RECT 31.245 149.305 31.535 150.030 ;
        RECT 33.290 149.850 33.630 150.680 ;
        RECT 35.110 150.170 35.460 151.420 ;
        RECT 38.810 149.850 39.150 150.680 ;
        RECT 40.630 150.170 40.980 151.420 ;
        RECT 44.330 149.850 44.670 150.680 ;
        RECT 46.150 150.170 46.500 151.420 ;
        RECT 49.850 149.850 50.190 150.680 ;
        RECT 51.670 150.170 52.020 151.420 ;
        RECT 53.785 150.765 56.375 151.855 ;
        RECT 53.785 150.075 54.995 150.595 ;
        RECT 55.165 150.245 56.375 150.765 ;
        RECT 57.005 150.690 57.295 151.855 ;
        RECT 57.465 151.420 62.810 151.855 ;
        RECT 31.705 149.305 37.050 149.850 ;
        RECT 37.225 149.305 42.570 149.850 ;
        RECT 42.745 149.305 48.090 149.850 ;
        RECT 48.265 149.305 53.610 149.850 ;
        RECT 53.785 149.305 56.375 150.075 ;
        RECT 57.005 149.305 57.295 150.030 ;
        RECT 59.050 149.850 59.390 150.680 ;
        RECT 60.870 150.170 61.220 151.420 ;
        RECT 63.995 151.185 64.165 151.685 ;
        RECT 64.335 151.355 64.665 151.855 ;
        RECT 63.995 151.015 64.660 151.185 ;
        RECT 63.910 150.195 64.260 150.845 ;
        RECT 64.430 150.025 64.660 151.015 ;
        RECT 63.995 149.855 64.660 150.025 ;
        RECT 57.465 149.305 62.810 149.850 ;
        RECT 63.995 149.565 64.165 149.855 ;
        RECT 64.335 149.305 64.665 149.685 ;
        RECT 64.835 149.565 65.060 151.685 ;
        RECT 65.260 151.395 65.525 151.855 ;
        RECT 65.710 151.285 65.945 151.660 ;
        RECT 66.190 151.410 67.260 151.580 ;
        RECT 65.260 150.285 65.540 150.885 ;
        RECT 65.275 149.305 65.525 149.765 ;
        RECT 65.710 149.755 65.880 151.285 ;
        RECT 66.050 150.255 66.290 151.125 ;
        RECT 66.480 150.875 66.920 151.230 ;
        RECT 67.090 150.795 67.260 151.410 ;
        RECT 67.430 151.055 67.600 151.855 ;
        RECT 67.770 151.355 68.020 151.685 ;
        RECT 68.245 151.385 69.130 151.555 ;
        RECT 67.090 150.705 67.600 150.795 ;
        RECT 66.800 150.535 67.600 150.705 ;
        RECT 66.050 149.925 66.630 150.255 ;
        RECT 66.800 149.755 66.970 150.535 ;
        RECT 67.430 150.465 67.600 150.535 ;
        RECT 67.140 150.285 67.310 150.315 ;
        RECT 67.770 150.285 67.940 151.355 ;
        RECT 68.110 150.465 68.300 151.185 ;
        RECT 68.470 150.795 68.790 151.125 ;
        RECT 67.140 149.985 67.940 150.285 ;
        RECT 68.470 150.255 68.660 150.795 ;
        RECT 65.710 149.585 66.040 149.755 ;
        RECT 66.220 149.585 66.970 149.755 ;
        RECT 67.220 149.305 67.590 149.805 ;
        RECT 67.770 149.755 67.940 149.985 ;
        RECT 68.110 149.925 68.660 150.255 ;
        RECT 68.960 150.465 69.130 151.385 ;
        RECT 69.310 151.355 69.525 151.855 ;
        RECT 69.990 151.050 70.160 151.675 ;
        RECT 70.445 151.075 70.625 151.855 ;
        RECT 69.300 150.890 70.160 151.050 ;
        RECT 69.300 150.720 70.410 150.890 ;
        RECT 70.240 150.465 70.410 150.720 ;
        RECT 70.805 150.855 71.140 151.615 ;
        RECT 71.320 151.025 71.490 151.855 ;
        RECT 71.660 150.855 71.990 151.615 ;
        RECT 72.160 151.025 72.330 151.855 ;
        RECT 72.645 151.420 77.990 151.855 ;
        RECT 70.805 150.685 72.475 150.855 ;
        RECT 68.960 150.295 70.050 150.465 ;
        RECT 70.240 150.295 72.060 150.465 ;
        RECT 68.960 149.755 69.130 150.295 ;
        RECT 70.240 150.125 70.410 150.295 ;
        RECT 69.910 149.955 70.410 150.125 ;
        RECT 72.230 150.120 72.475 150.685 ;
        RECT 67.770 149.585 68.230 149.755 ;
        RECT 68.460 149.585 69.130 149.755 ;
        RECT 69.445 149.305 69.615 149.835 ;
        RECT 69.910 149.515 70.270 149.955 ;
        RECT 70.805 149.950 72.475 150.120 ;
        RECT 70.445 149.305 70.615 149.785 ;
        RECT 70.805 149.525 71.140 149.950 ;
        RECT 71.315 149.305 71.485 149.780 ;
        RECT 71.660 149.525 71.995 149.950 ;
        RECT 74.230 149.850 74.570 150.680 ;
        RECT 76.050 150.170 76.400 151.420 ;
        RECT 78.165 150.765 81.675 151.855 ;
        RECT 78.165 150.075 79.815 150.595 ;
        RECT 79.985 150.245 81.675 150.765 ;
        RECT 82.765 150.690 83.055 151.855 ;
        RECT 83.225 151.420 88.570 151.855 ;
        RECT 72.165 149.305 72.335 149.780 ;
        RECT 72.645 149.305 77.990 149.850 ;
        RECT 78.165 149.305 81.675 150.075 ;
        RECT 82.765 149.305 83.055 150.030 ;
        RECT 84.810 149.850 85.150 150.680 ;
        RECT 86.630 150.170 86.980 151.420 ;
        RECT 88.745 150.765 90.415 151.855 ;
        RECT 88.745 150.075 89.495 150.595 ;
        RECT 89.665 150.245 90.415 150.765 ;
        RECT 91.045 150.765 92.255 151.855 ;
        RECT 91.045 150.225 91.565 150.765 ;
        RECT 83.225 149.305 88.570 149.850 ;
        RECT 88.745 149.305 90.415 150.075 ;
        RECT 91.735 150.055 92.255 150.595 ;
        RECT 91.045 149.305 92.255 150.055 ;
        RECT 18.280 149.135 92.340 149.305 ;
        RECT 18.365 148.385 19.575 149.135 ;
        RECT 19.745 148.590 25.090 149.135 ;
        RECT 25.265 148.590 30.610 149.135 ;
        RECT 30.785 148.590 36.130 149.135 ;
        RECT 36.305 148.590 41.650 149.135 ;
        RECT 18.365 147.845 18.885 148.385 ;
        RECT 19.055 147.675 19.575 148.215 ;
        RECT 21.330 147.760 21.670 148.590 ;
        RECT 18.365 146.585 19.575 147.675 ;
        RECT 23.150 147.020 23.500 148.270 ;
        RECT 26.850 147.760 27.190 148.590 ;
        RECT 28.670 147.020 29.020 148.270 ;
        RECT 32.370 147.760 32.710 148.590 ;
        RECT 34.190 147.020 34.540 148.270 ;
        RECT 37.890 147.760 38.230 148.590 ;
        RECT 41.825 148.365 43.495 149.135 ;
        RECT 44.125 148.410 44.415 149.135 ;
        RECT 44.585 148.590 49.930 149.135 ;
        RECT 50.105 148.590 55.450 149.135 ;
        RECT 55.625 148.590 60.970 149.135 ;
        RECT 61.145 148.590 66.490 149.135 ;
        RECT 39.710 147.020 40.060 148.270 ;
        RECT 41.825 147.845 42.575 148.365 ;
        RECT 42.745 147.675 43.495 148.195 ;
        RECT 46.170 147.760 46.510 148.590 ;
        RECT 19.745 146.585 25.090 147.020 ;
        RECT 25.265 146.585 30.610 147.020 ;
        RECT 30.785 146.585 36.130 147.020 ;
        RECT 36.305 146.585 41.650 147.020 ;
        RECT 41.825 146.585 43.495 147.675 ;
        RECT 44.125 146.585 44.415 147.750 ;
        RECT 47.990 147.020 48.340 148.270 ;
        RECT 51.690 147.760 52.030 148.590 ;
        RECT 53.510 147.020 53.860 148.270 ;
        RECT 57.210 147.760 57.550 148.590 ;
        RECT 59.030 147.020 59.380 148.270 ;
        RECT 62.730 147.760 63.070 148.590 ;
        RECT 66.665 148.365 69.255 149.135 ;
        RECT 69.885 148.410 70.175 149.135 ;
        RECT 70.345 148.590 75.690 149.135 ;
        RECT 75.865 148.590 81.210 149.135 ;
        RECT 81.385 148.590 86.730 149.135 ;
        RECT 64.550 147.020 64.900 148.270 ;
        RECT 66.665 147.845 67.875 148.365 ;
        RECT 68.045 147.675 69.255 148.195 ;
        RECT 71.930 147.760 72.270 148.590 ;
        RECT 44.585 146.585 49.930 147.020 ;
        RECT 50.105 146.585 55.450 147.020 ;
        RECT 55.625 146.585 60.970 147.020 ;
        RECT 61.145 146.585 66.490 147.020 ;
        RECT 66.665 146.585 69.255 147.675 ;
        RECT 69.885 146.585 70.175 147.750 ;
        RECT 73.750 147.020 74.100 148.270 ;
        RECT 77.450 147.760 77.790 148.590 ;
        RECT 79.270 147.020 79.620 148.270 ;
        RECT 82.970 147.760 83.310 148.590 ;
        RECT 86.905 148.365 90.415 149.135 ;
        RECT 91.045 148.385 92.255 149.135 ;
        RECT 84.790 147.020 85.140 148.270 ;
        RECT 86.905 147.845 88.555 148.365 ;
        RECT 88.725 147.675 90.415 148.195 ;
        RECT 70.345 146.585 75.690 147.020 ;
        RECT 75.865 146.585 81.210 147.020 ;
        RECT 81.385 146.585 86.730 147.020 ;
        RECT 86.905 146.585 90.415 147.675 ;
        RECT 91.045 147.675 91.565 148.215 ;
        RECT 91.735 147.845 92.255 148.385 ;
        RECT 91.045 146.585 92.255 147.675 ;
        RECT 18.280 146.415 92.340 146.585 ;
        RECT 18.365 145.325 19.575 146.415 ;
        RECT 19.745 145.980 25.090 146.415 ;
        RECT 25.265 145.980 30.610 146.415 ;
        RECT 18.365 144.615 18.885 145.155 ;
        RECT 19.055 144.785 19.575 145.325 ;
        RECT 18.365 143.865 19.575 144.615 ;
        RECT 21.330 144.410 21.670 145.240 ;
        RECT 23.150 144.730 23.500 145.980 ;
        RECT 26.850 144.410 27.190 145.240 ;
        RECT 28.670 144.730 29.020 145.980 ;
        RECT 31.245 145.250 31.535 146.415 ;
        RECT 31.705 145.980 37.050 146.415 ;
        RECT 37.225 145.980 42.570 146.415 ;
        RECT 42.745 145.980 48.090 146.415 ;
        RECT 48.265 145.980 53.610 146.415 ;
        RECT 19.745 143.865 25.090 144.410 ;
        RECT 25.265 143.865 30.610 144.410 ;
        RECT 31.245 143.865 31.535 144.590 ;
        RECT 33.290 144.410 33.630 145.240 ;
        RECT 35.110 144.730 35.460 145.980 ;
        RECT 38.810 144.410 39.150 145.240 ;
        RECT 40.630 144.730 40.980 145.980 ;
        RECT 44.330 144.410 44.670 145.240 ;
        RECT 46.150 144.730 46.500 145.980 ;
        RECT 49.850 144.410 50.190 145.240 ;
        RECT 51.670 144.730 52.020 145.980 ;
        RECT 53.785 145.325 56.375 146.415 ;
        RECT 53.785 144.635 54.995 145.155 ;
        RECT 55.165 144.805 56.375 145.325 ;
        RECT 57.005 145.250 57.295 146.415 ;
        RECT 57.465 145.980 62.810 146.415 ;
        RECT 62.985 145.980 68.330 146.415 ;
        RECT 68.505 145.980 73.850 146.415 ;
        RECT 74.025 145.980 79.370 146.415 ;
        RECT 31.705 143.865 37.050 144.410 ;
        RECT 37.225 143.865 42.570 144.410 ;
        RECT 42.745 143.865 48.090 144.410 ;
        RECT 48.265 143.865 53.610 144.410 ;
        RECT 53.785 143.865 56.375 144.635 ;
        RECT 57.005 143.865 57.295 144.590 ;
        RECT 59.050 144.410 59.390 145.240 ;
        RECT 60.870 144.730 61.220 145.980 ;
        RECT 64.570 144.410 64.910 145.240 ;
        RECT 66.390 144.730 66.740 145.980 ;
        RECT 70.090 144.410 70.430 145.240 ;
        RECT 71.910 144.730 72.260 145.980 ;
        RECT 75.610 144.410 75.950 145.240 ;
        RECT 77.430 144.730 77.780 145.980 ;
        RECT 79.545 145.325 82.135 146.415 ;
        RECT 79.545 144.635 80.755 145.155 ;
        RECT 80.925 144.805 82.135 145.325 ;
        RECT 82.765 145.250 83.055 146.415 ;
        RECT 83.225 145.980 88.570 146.415 ;
        RECT 57.465 143.865 62.810 144.410 ;
        RECT 62.985 143.865 68.330 144.410 ;
        RECT 68.505 143.865 73.850 144.410 ;
        RECT 74.025 143.865 79.370 144.410 ;
        RECT 79.545 143.865 82.135 144.635 ;
        RECT 82.765 143.865 83.055 144.590 ;
        RECT 84.810 144.410 85.150 145.240 ;
        RECT 86.630 144.730 86.980 145.980 ;
        RECT 88.745 145.325 90.415 146.415 ;
        RECT 88.745 144.635 89.495 145.155 ;
        RECT 89.665 144.805 90.415 145.325 ;
        RECT 91.045 145.325 92.255 146.415 ;
        RECT 91.045 144.785 91.565 145.325 ;
        RECT 83.225 143.865 88.570 144.410 ;
        RECT 88.745 143.865 90.415 144.635 ;
        RECT 91.735 144.615 92.255 145.155 ;
        RECT 91.045 143.865 92.255 144.615 ;
        RECT 18.280 143.695 92.340 143.865 ;
        RECT 18.365 142.945 19.575 143.695 ;
        RECT 19.745 143.150 25.090 143.695 ;
        RECT 25.265 143.150 30.610 143.695 ;
        RECT 30.785 143.150 36.130 143.695 ;
        RECT 36.305 143.150 41.650 143.695 ;
        RECT 18.365 142.405 18.885 142.945 ;
        RECT 19.055 142.235 19.575 142.775 ;
        RECT 21.330 142.320 21.670 143.150 ;
        RECT 18.365 141.145 19.575 142.235 ;
        RECT 23.150 141.580 23.500 142.830 ;
        RECT 26.850 142.320 27.190 143.150 ;
        RECT 28.670 141.580 29.020 142.830 ;
        RECT 32.370 142.320 32.710 143.150 ;
        RECT 34.190 141.580 34.540 142.830 ;
        RECT 37.890 142.320 38.230 143.150 ;
        RECT 41.825 142.925 43.495 143.695 ;
        RECT 44.125 142.970 44.415 143.695 ;
        RECT 44.585 143.150 49.930 143.695 ;
        RECT 50.105 143.150 55.450 143.695 ;
        RECT 55.625 143.150 60.970 143.695 ;
        RECT 61.145 143.150 66.490 143.695 ;
        RECT 39.710 141.580 40.060 142.830 ;
        RECT 41.825 142.405 42.575 142.925 ;
        RECT 42.745 142.235 43.495 142.755 ;
        RECT 46.170 142.320 46.510 143.150 ;
        RECT 19.745 141.145 25.090 141.580 ;
        RECT 25.265 141.145 30.610 141.580 ;
        RECT 30.785 141.145 36.130 141.580 ;
        RECT 36.305 141.145 41.650 141.580 ;
        RECT 41.825 141.145 43.495 142.235 ;
        RECT 44.125 141.145 44.415 142.310 ;
        RECT 47.990 141.580 48.340 142.830 ;
        RECT 51.690 142.320 52.030 143.150 ;
        RECT 53.510 141.580 53.860 142.830 ;
        RECT 57.210 142.320 57.550 143.150 ;
        RECT 59.030 141.580 59.380 142.830 ;
        RECT 62.730 142.320 63.070 143.150 ;
        RECT 66.665 142.925 69.255 143.695 ;
        RECT 69.885 142.970 70.175 143.695 ;
        RECT 70.345 143.150 75.690 143.695 ;
        RECT 75.865 143.150 81.210 143.695 ;
        RECT 81.385 143.150 86.730 143.695 ;
        RECT 64.550 141.580 64.900 142.830 ;
        RECT 66.665 142.405 67.875 142.925 ;
        RECT 68.045 142.235 69.255 142.755 ;
        RECT 71.930 142.320 72.270 143.150 ;
        RECT 44.585 141.145 49.930 141.580 ;
        RECT 50.105 141.145 55.450 141.580 ;
        RECT 55.625 141.145 60.970 141.580 ;
        RECT 61.145 141.145 66.490 141.580 ;
        RECT 66.665 141.145 69.255 142.235 ;
        RECT 69.885 141.145 70.175 142.310 ;
        RECT 73.750 141.580 74.100 142.830 ;
        RECT 77.450 142.320 77.790 143.150 ;
        RECT 79.270 141.580 79.620 142.830 ;
        RECT 82.970 142.320 83.310 143.150 ;
        RECT 86.905 142.925 90.415 143.695 ;
        RECT 91.045 142.945 92.255 143.695 ;
        RECT 84.790 141.580 85.140 142.830 ;
        RECT 86.905 142.405 88.555 142.925 ;
        RECT 88.725 142.235 90.415 142.755 ;
        RECT 70.345 141.145 75.690 141.580 ;
        RECT 75.865 141.145 81.210 141.580 ;
        RECT 81.385 141.145 86.730 141.580 ;
        RECT 86.905 141.145 90.415 142.235 ;
        RECT 91.045 142.235 91.565 142.775 ;
        RECT 91.735 142.405 92.255 142.945 ;
        RECT 112.990 142.690 113.340 144.850 ;
        RECT 113.990 142.690 114.340 144.850 ;
        RECT 114.990 142.690 115.340 144.850 ;
        RECT 115.990 142.690 116.340 144.850 ;
        RECT 116.990 142.690 117.340 144.850 ;
        RECT 117.990 142.690 118.340 144.850 ;
        RECT 118.990 142.690 119.340 144.850 ;
        RECT 119.990 142.690 120.340 144.850 ;
        RECT 91.045 141.145 92.255 142.235 ;
        RECT 18.280 140.975 92.340 141.145 ;
        RECT 18.365 139.885 19.575 140.975 ;
        RECT 19.745 140.540 25.090 140.975 ;
        RECT 25.265 140.540 30.610 140.975 ;
        RECT 18.365 139.175 18.885 139.715 ;
        RECT 19.055 139.345 19.575 139.885 ;
        RECT 18.365 138.425 19.575 139.175 ;
        RECT 21.330 138.970 21.670 139.800 ;
        RECT 23.150 139.290 23.500 140.540 ;
        RECT 26.850 138.970 27.190 139.800 ;
        RECT 28.670 139.290 29.020 140.540 ;
        RECT 31.245 139.810 31.535 140.975 ;
        RECT 31.705 140.540 37.050 140.975 ;
        RECT 37.225 140.540 42.570 140.975 ;
        RECT 42.745 140.540 48.090 140.975 ;
        RECT 48.265 140.540 53.610 140.975 ;
        RECT 19.745 138.425 25.090 138.970 ;
        RECT 25.265 138.425 30.610 138.970 ;
        RECT 31.245 138.425 31.535 139.150 ;
        RECT 33.290 138.970 33.630 139.800 ;
        RECT 35.110 139.290 35.460 140.540 ;
        RECT 38.810 138.970 39.150 139.800 ;
        RECT 40.630 139.290 40.980 140.540 ;
        RECT 44.330 138.970 44.670 139.800 ;
        RECT 46.150 139.290 46.500 140.540 ;
        RECT 49.850 138.970 50.190 139.800 ;
        RECT 51.670 139.290 52.020 140.540 ;
        RECT 53.785 139.885 56.375 140.975 ;
        RECT 53.785 139.195 54.995 139.715 ;
        RECT 55.165 139.365 56.375 139.885 ;
        RECT 57.005 139.810 57.295 140.975 ;
        RECT 57.465 140.540 62.810 140.975 ;
        RECT 62.985 140.540 68.330 140.975 ;
        RECT 68.505 140.540 73.850 140.975 ;
        RECT 74.025 140.540 79.370 140.975 ;
        RECT 31.705 138.425 37.050 138.970 ;
        RECT 37.225 138.425 42.570 138.970 ;
        RECT 42.745 138.425 48.090 138.970 ;
        RECT 48.265 138.425 53.610 138.970 ;
        RECT 53.785 138.425 56.375 139.195 ;
        RECT 57.005 138.425 57.295 139.150 ;
        RECT 59.050 138.970 59.390 139.800 ;
        RECT 60.870 139.290 61.220 140.540 ;
        RECT 64.570 138.970 64.910 139.800 ;
        RECT 66.390 139.290 66.740 140.540 ;
        RECT 70.090 138.970 70.430 139.800 ;
        RECT 71.910 139.290 72.260 140.540 ;
        RECT 75.610 138.970 75.950 139.800 ;
        RECT 77.430 139.290 77.780 140.540 ;
        RECT 79.545 139.885 82.135 140.975 ;
        RECT 79.545 139.195 80.755 139.715 ;
        RECT 80.925 139.365 82.135 139.885 ;
        RECT 82.765 139.810 83.055 140.975 ;
        RECT 83.225 140.540 88.570 140.975 ;
        RECT 57.465 138.425 62.810 138.970 ;
        RECT 62.985 138.425 68.330 138.970 ;
        RECT 68.505 138.425 73.850 138.970 ;
        RECT 74.025 138.425 79.370 138.970 ;
        RECT 79.545 138.425 82.135 139.195 ;
        RECT 82.765 138.425 83.055 139.150 ;
        RECT 84.810 138.970 85.150 139.800 ;
        RECT 86.630 139.290 86.980 140.540 ;
        RECT 88.745 139.885 90.415 140.975 ;
        RECT 88.745 139.195 89.495 139.715 ;
        RECT 89.665 139.365 90.415 139.885 ;
        RECT 91.045 139.885 92.255 140.975 ;
        RECT 91.045 139.345 91.565 139.885 ;
        RECT 83.225 138.425 88.570 138.970 ;
        RECT 88.745 138.425 90.415 139.195 ;
        RECT 91.735 139.175 92.255 139.715 ;
        RECT 112.990 139.530 113.340 141.690 ;
        RECT 113.990 139.530 114.340 141.690 ;
        RECT 114.990 139.530 115.340 141.690 ;
        RECT 115.990 139.530 116.340 141.690 ;
        RECT 116.990 139.530 117.340 141.690 ;
        RECT 117.990 139.530 118.340 141.690 ;
        RECT 118.990 139.530 119.340 141.690 ;
        RECT 119.990 139.530 120.340 141.690 ;
        RECT 91.045 138.425 92.255 139.175 ;
        RECT 18.280 138.255 92.340 138.425 ;
        RECT 18.365 137.505 19.575 138.255 ;
        RECT 19.745 137.710 25.090 138.255 ;
        RECT 25.265 137.710 30.610 138.255 ;
        RECT 30.785 137.710 36.130 138.255 ;
        RECT 36.305 137.710 41.650 138.255 ;
        RECT 18.365 136.965 18.885 137.505 ;
        RECT 19.055 136.795 19.575 137.335 ;
        RECT 21.330 136.880 21.670 137.710 ;
        RECT 18.365 135.705 19.575 136.795 ;
        RECT 23.150 136.140 23.500 137.390 ;
        RECT 26.850 136.880 27.190 137.710 ;
        RECT 28.670 136.140 29.020 137.390 ;
        RECT 32.370 136.880 32.710 137.710 ;
        RECT 34.190 136.140 34.540 137.390 ;
        RECT 37.890 136.880 38.230 137.710 ;
        RECT 41.825 137.485 43.495 138.255 ;
        RECT 44.125 137.530 44.415 138.255 ;
        RECT 44.585 137.710 49.930 138.255 ;
        RECT 50.105 137.710 55.450 138.255 ;
        RECT 55.625 137.710 60.970 138.255 ;
        RECT 61.145 137.710 66.490 138.255 ;
        RECT 39.710 136.140 40.060 137.390 ;
        RECT 41.825 136.965 42.575 137.485 ;
        RECT 42.745 136.795 43.495 137.315 ;
        RECT 46.170 136.880 46.510 137.710 ;
        RECT 19.745 135.705 25.090 136.140 ;
        RECT 25.265 135.705 30.610 136.140 ;
        RECT 30.785 135.705 36.130 136.140 ;
        RECT 36.305 135.705 41.650 136.140 ;
        RECT 41.825 135.705 43.495 136.795 ;
        RECT 44.125 135.705 44.415 136.870 ;
        RECT 47.990 136.140 48.340 137.390 ;
        RECT 51.690 136.880 52.030 137.710 ;
        RECT 53.510 136.140 53.860 137.390 ;
        RECT 57.210 136.880 57.550 137.710 ;
        RECT 59.030 136.140 59.380 137.390 ;
        RECT 62.730 136.880 63.070 137.710 ;
        RECT 66.665 137.485 69.255 138.255 ;
        RECT 69.885 137.530 70.175 138.255 ;
        RECT 70.345 137.710 75.690 138.255 ;
        RECT 75.865 137.710 81.210 138.255 ;
        RECT 81.385 137.710 86.730 138.255 ;
        RECT 64.550 136.140 64.900 137.390 ;
        RECT 66.665 136.965 67.875 137.485 ;
        RECT 68.045 136.795 69.255 137.315 ;
        RECT 71.930 136.880 72.270 137.710 ;
        RECT 44.585 135.705 49.930 136.140 ;
        RECT 50.105 135.705 55.450 136.140 ;
        RECT 55.625 135.705 60.970 136.140 ;
        RECT 61.145 135.705 66.490 136.140 ;
        RECT 66.665 135.705 69.255 136.795 ;
        RECT 69.885 135.705 70.175 136.870 ;
        RECT 73.750 136.140 74.100 137.390 ;
        RECT 77.450 136.880 77.790 137.710 ;
        RECT 79.270 136.140 79.620 137.390 ;
        RECT 82.970 136.880 83.310 137.710 ;
        RECT 86.905 137.485 90.415 138.255 ;
        RECT 91.045 137.505 92.255 138.255 ;
        RECT 84.790 136.140 85.140 137.390 ;
        RECT 86.905 136.965 88.555 137.485 ;
        RECT 88.725 136.795 90.415 137.315 ;
        RECT 70.345 135.705 75.690 136.140 ;
        RECT 75.865 135.705 81.210 136.140 ;
        RECT 81.385 135.705 86.730 136.140 ;
        RECT 86.905 135.705 90.415 136.795 ;
        RECT 91.045 136.795 91.565 137.335 ;
        RECT 91.735 136.965 92.255 137.505 ;
        RECT 91.045 135.705 92.255 136.795 ;
        RECT 112.990 136.690 113.340 138.850 ;
        RECT 113.990 136.190 114.340 138.350 ;
        RECT 114.990 136.190 115.340 138.350 ;
        RECT 115.990 136.190 116.340 138.350 ;
        RECT 116.990 136.190 117.340 138.350 ;
        RECT 117.990 136.190 118.340 138.350 ;
        RECT 118.990 136.190 119.340 138.350 ;
        RECT 119.990 136.190 120.340 138.350 ;
        RECT 18.280 135.535 92.340 135.705 ;
        RECT 18.365 134.445 19.575 135.535 ;
        RECT 19.745 135.100 25.090 135.535 ;
        RECT 25.265 135.100 30.610 135.535 ;
        RECT 18.365 133.735 18.885 134.275 ;
        RECT 19.055 133.905 19.575 134.445 ;
        RECT 18.365 132.985 19.575 133.735 ;
        RECT 21.330 133.530 21.670 134.360 ;
        RECT 23.150 133.850 23.500 135.100 ;
        RECT 26.850 133.530 27.190 134.360 ;
        RECT 28.670 133.850 29.020 135.100 ;
        RECT 31.245 134.370 31.535 135.535 ;
        RECT 31.705 135.100 37.050 135.535 ;
        RECT 37.225 135.100 42.570 135.535 ;
        RECT 19.745 132.985 25.090 133.530 ;
        RECT 25.265 132.985 30.610 133.530 ;
        RECT 31.245 132.985 31.535 133.710 ;
        RECT 33.290 133.530 33.630 134.360 ;
        RECT 35.110 133.850 35.460 135.100 ;
        RECT 38.810 133.530 39.150 134.360 ;
        RECT 40.630 133.850 40.980 135.100 ;
        RECT 42.745 134.445 43.955 135.535 ;
        RECT 42.745 133.735 43.265 134.275 ;
        RECT 43.435 133.905 43.955 134.445 ;
        RECT 44.125 134.370 44.415 135.535 ;
        RECT 44.585 135.100 49.930 135.535 ;
        RECT 50.105 135.100 55.450 135.535 ;
        RECT 31.705 132.985 37.050 133.530 ;
        RECT 37.225 132.985 42.570 133.530 ;
        RECT 42.745 132.985 43.955 133.735 ;
        RECT 44.125 132.985 44.415 133.710 ;
        RECT 46.170 133.530 46.510 134.360 ;
        RECT 47.990 133.850 48.340 135.100 ;
        RECT 51.690 133.530 52.030 134.360 ;
        RECT 53.510 133.850 53.860 135.100 ;
        RECT 55.625 134.445 56.835 135.535 ;
        RECT 55.625 133.735 56.145 134.275 ;
        RECT 56.315 133.905 56.835 134.445 ;
        RECT 57.005 134.370 57.295 135.535 ;
        RECT 57.465 135.100 62.810 135.535 ;
        RECT 62.985 135.100 68.330 135.535 ;
        RECT 44.585 132.985 49.930 133.530 ;
        RECT 50.105 132.985 55.450 133.530 ;
        RECT 55.625 132.985 56.835 133.735 ;
        RECT 57.005 132.985 57.295 133.710 ;
        RECT 59.050 133.530 59.390 134.360 ;
        RECT 60.870 133.850 61.220 135.100 ;
        RECT 64.570 133.530 64.910 134.360 ;
        RECT 66.390 133.850 66.740 135.100 ;
        RECT 68.505 134.445 69.715 135.535 ;
        RECT 68.505 133.735 69.025 134.275 ;
        RECT 69.195 133.905 69.715 134.445 ;
        RECT 69.885 134.370 70.175 135.535 ;
        RECT 70.345 135.100 75.690 135.535 ;
        RECT 75.865 135.100 81.210 135.535 ;
        RECT 57.465 132.985 62.810 133.530 ;
        RECT 62.985 132.985 68.330 133.530 ;
        RECT 68.505 132.985 69.715 133.735 ;
        RECT 69.885 132.985 70.175 133.710 ;
        RECT 71.930 133.530 72.270 134.360 ;
        RECT 73.750 133.850 74.100 135.100 ;
        RECT 77.450 133.530 77.790 134.360 ;
        RECT 79.270 133.850 79.620 135.100 ;
        RECT 81.385 134.445 82.595 135.535 ;
        RECT 81.385 133.735 81.905 134.275 ;
        RECT 82.075 133.905 82.595 134.445 ;
        RECT 82.765 134.370 83.055 135.535 ;
        RECT 83.225 135.100 88.570 135.535 ;
        RECT 70.345 132.985 75.690 133.530 ;
        RECT 75.865 132.985 81.210 133.530 ;
        RECT 81.385 132.985 82.595 133.735 ;
        RECT 82.765 132.985 83.055 133.710 ;
        RECT 84.810 133.530 85.150 134.360 ;
        RECT 86.630 133.850 86.980 135.100 ;
        RECT 88.745 134.445 90.415 135.535 ;
        RECT 88.745 133.755 89.495 134.275 ;
        RECT 89.665 133.925 90.415 134.445 ;
        RECT 91.045 134.445 92.255 135.535 ;
        RECT 91.045 133.905 91.565 134.445 ;
        RECT 83.225 132.985 88.570 133.530 ;
        RECT 88.745 132.985 90.415 133.755 ;
        RECT 91.735 133.735 92.255 134.275 ;
        RECT 91.045 132.985 92.255 133.735 ;
        RECT 112.990 133.530 113.340 135.690 ;
        RECT 113.990 133.530 114.340 135.690 ;
        RECT 114.990 133.530 115.340 135.690 ;
        RECT 115.990 133.530 116.340 135.690 ;
        RECT 116.990 133.530 117.340 135.690 ;
        RECT 117.990 133.530 118.340 135.690 ;
        RECT 118.990 133.530 119.340 135.690 ;
        RECT 119.990 133.530 120.340 135.690 ;
        RECT 18.280 132.815 92.340 132.985 ;
      LAYER mcon ;
        RECT 18.425 206.255 18.595 206.425 ;
        RECT 18.885 206.255 19.055 206.425 ;
        RECT 19.345 206.255 19.515 206.425 ;
        RECT 19.805 206.255 19.975 206.425 ;
        RECT 20.265 206.255 20.435 206.425 ;
        RECT 20.725 206.255 20.895 206.425 ;
        RECT 21.185 206.255 21.355 206.425 ;
        RECT 21.645 206.255 21.815 206.425 ;
        RECT 22.105 206.255 22.275 206.425 ;
        RECT 22.565 206.255 22.735 206.425 ;
        RECT 23.025 206.255 23.195 206.425 ;
        RECT 23.485 206.255 23.655 206.425 ;
        RECT 23.945 206.255 24.115 206.425 ;
        RECT 24.405 206.255 24.575 206.425 ;
        RECT 24.865 206.255 25.035 206.425 ;
        RECT 25.325 206.255 25.495 206.425 ;
        RECT 25.785 206.255 25.955 206.425 ;
        RECT 26.245 206.255 26.415 206.425 ;
        RECT 26.705 206.255 26.875 206.425 ;
        RECT 27.165 206.255 27.335 206.425 ;
        RECT 27.625 206.255 27.795 206.425 ;
        RECT 28.085 206.255 28.255 206.425 ;
        RECT 28.545 206.255 28.715 206.425 ;
        RECT 29.005 206.255 29.175 206.425 ;
        RECT 29.465 206.255 29.635 206.425 ;
        RECT 29.925 206.255 30.095 206.425 ;
        RECT 30.385 206.255 30.555 206.425 ;
        RECT 30.845 206.255 31.015 206.425 ;
        RECT 31.305 206.255 31.475 206.425 ;
        RECT 31.765 206.255 31.935 206.425 ;
        RECT 32.225 206.255 32.395 206.425 ;
        RECT 32.685 206.255 32.855 206.425 ;
        RECT 33.145 206.255 33.315 206.425 ;
        RECT 33.605 206.255 33.775 206.425 ;
        RECT 34.065 206.255 34.235 206.425 ;
        RECT 34.525 206.255 34.695 206.425 ;
        RECT 34.985 206.255 35.155 206.425 ;
        RECT 35.445 206.255 35.615 206.425 ;
        RECT 35.905 206.255 36.075 206.425 ;
        RECT 36.365 206.255 36.535 206.425 ;
        RECT 36.825 206.255 36.995 206.425 ;
        RECT 37.285 206.255 37.455 206.425 ;
        RECT 37.745 206.255 37.915 206.425 ;
        RECT 38.205 206.255 38.375 206.425 ;
        RECT 38.665 206.255 38.835 206.425 ;
        RECT 39.125 206.255 39.295 206.425 ;
        RECT 39.585 206.255 39.755 206.425 ;
        RECT 40.045 206.255 40.215 206.425 ;
        RECT 40.505 206.255 40.675 206.425 ;
        RECT 40.965 206.255 41.135 206.425 ;
        RECT 41.425 206.255 41.595 206.425 ;
        RECT 41.885 206.255 42.055 206.425 ;
        RECT 42.345 206.255 42.515 206.425 ;
        RECT 42.805 206.255 42.975 206.425 ;
        RECT 43.265 206.255 43.435 206.425 ;
        RECT 43.725 206.255 43.895 206.425 ;
        RECT 44.185 206.255 44.355 206.425 ;
        RECT 44.645 206.255 44.815 206.425 ;
        RECT 45.105 206.255 45.275 206.425 ;
        RECT 45.565 206.255 45.735 206.425 ;
        RECT 46.025 206.255 46.195 206.425 ;
        RECT 46.485 206.255 46.655 206.425 ;
        RECT 46.945 206.255 47.115 206.425 ;
        RECT 47.405 206.255 47.575 206.425 ;
        RECT 47.865 206.255 48.035 206.425 ;
        RECT 48.325 206.255 48.495 206.425 ;
        RECT 48.785 206.255 48.955 206.425 ;
        RECT 49.245 206.255 49.415 206.425 ;
        RECT 49.705 206.255 49.875 206.425 ;
        RECT 50.165 206.255 50.335 206.425 ;
        RECT 50.625 206.255 50.795 206.425 ;
        RECT 51.085 206.255 51.255 206.425 ;
        RECT 51.545 206.255 51.715 206.425 ;
        RECT 52.005 206.255 52.175 206.425 ;
        RECT 52.465 206.255 52.635 206.425 ;
        RECT 52.925 206.255 53.095 206.425 ;
        RECT 53.385 206.255 53.555 206.425 ;
        RECT 53.845 206.255 54.015 206.425 ;
        RECT 54.305 206.255 54.475 206.425 ;
        RECT 54.765 206.255 54.935 206.425 ;
        RECT 55.225 206.255 55.395 206.425 ;
        RECT 55.685 206.255 55.855 206.425 ;
        RECT 56.145 206.255 56.315 206.425 ;
        RECT 56.605 206.255 56.775 206.425 ;
        RECT 57.065 206.255 57.235 206.425 ;
        RECT 57.525 206.255 57.695 206.425 ;
        RECT 57.985 206.255 58.155 206.425 ;
        RECT 58.445 206.255 58.615 206.425 ;
        RECT 58.905 206.255 59.075 206.425 ;
        RECT 59.365 206.255 59.535 206.425 ;
        RECT 59.825 206.255 59.995 206.425 ;
        RECT 60.285 206.255 60.455 206.425 ;
        RECT 60.745 206.255 60.915 206.425 ;
        RECT 61.205 206.255 61.375 206.425 ;
        RECT 61.665 206.255 61.835 206.425 ;
        RECT 62.125 206.255 62.295 206.425 ;
        RECT 62.585 206.255 62.755 206.425 ;
        RECT 63.045 206.255 63.215 206.425 ;
        RECT 63.505 206.255 63.675 206.425 ;
        RECT 63.965 206.255 64.135 206.425 ;
        RECT 64.425 206.255 64.595 206.425 ;
        RECT 64.885 206.255 65.055 206.425 ;
        RECT 65.345 206.255 65.515 206.425 ;
        RECT 65.805 206.255 65.975 206.425 ;
        RECT 66.265 206.255 66.435 206.425 ;
        RECT 66.725 206.255 66.895 206.425 ;
        RECT 67.185 206.255 67.355 206.425 ;
        RECT 67.645 206.255 67.815 206.425 ;
        RECT 68.105 206.255 68.275 206.425 ;
        RECT 68.565 206.255 68.735 206.425 ;
        RECT 69.025 206.255 69.195 206.425 ;
        RECT 69.485 206.255 69.655 206.425 ;
        RECT 69.945 206.255 70.115 206.425 ;
        RECT 70.405 206.255 70.575 206.425 ;
        RECT 70.865 206.255 71.035 206.425 ;
        RECT 71.325 206.255 71.495 206.425 ;
        RECT 71.785 206.255 71.955 206.425 ;
        RECT 72.245 206.255 72.415 206.425 ;
        RECT 72.705 206.255 72.875 206.425 ;
        RECT 73.165 206.255 73.335 206.425 ;
        RECT 73.625 206.255 73.795 206.425 ;
        RECT 74.085 206.255 74.255 206.425 ;
        RECT 74.545 206.255 74.715 206.425 ;
        RECT 75.005 206.255 75.175 206.425 ;
        RECT 75.465 206.255 75.635 206.425 ;
        RECT 75.925 206.255 76.095 206.425 ;
        RECT 76.385 206.255 76.555 206.425 ;
        RECT 76.845 206.255 77.015 206.425 ;
        RECT 77.305 206.255 77.475 206.425 ;
        RECT 77.765 206.255 77.935 206.425 ;
        RECT 78.225 206.255 78.395 206.425 ;
        RECT 78.685 206.255 78.855 206.425 ;
        RECT 79.145 206.255 79.315 206.425 ;
        RECT 79.605 206.255 79.775 206.425 ;
        RECT 80.065 206.255 80.235 206.425 ;
        RECT 80.525 206.255 80.695 206.425 ;
        RECT 80.985 206.255 81.155 206.425 ;
        RECT 81.445 206.255 81.615 206.425 ;
        RECT 81.905 206.255 82.075 206.425 ;
        RECT 82.365 206.255 82.535 206.425 ;
        RECT 82.825 206.255 82.995 206.425 ;
        RECT 83.285 206.255 83.455 206.425 ;
        RECT 83.745 206.255 83.915 206.425 ;
        RECT 84.205 206.255 84.375 206.425 ;
        RECT 84.665 206.255 84.835 206.425 ;
        RECT 85.125 206.255 85.295 206.425 ;
        RECT 85.585 206.255 85.755 206.425 ;
        RECT 86.045 206.255 86.215 206.425 ;
        RECT 86.505 206.255 86.675 206.425 ;
        RECT 86.965 206.255 87.135 206.425 ;
        RECT 87.425 206.255 87.595 206.425 ;
        RECT 87.885 206.255 88.055 206.425 ;
        RECT 88.345 206.255 88.515 206.425 ;
        RECT 88.805 206.255 88.975 206.425 ;
        RECT 89.265 206.255 89.435 206.425 ;
        RECT 89.725 206.255 89.895 206.425 ;
        RECT 90.185 206.255 90.355 206.425 ;
        RECT 90.645 206.255 90.815 206.425 ;
        RECT 91.105 206.255 91.275 206.425 ;
        RECT 91.565 206.255 91.735 206.425 ;
        RECT 92.025 206.255 92.195 206.425 ;
        RECT 27.625 204.725 27.795 204.895 ;
        RECT 26.245 204.045 26.415 204.215 ;
        RECT 28.545 204.045 28.715 204.215 ;
        RECT 33.605 204.725 33.775 204.895 ;
        RECT 34.525 204.385 34.695 204.555 ;
        RECT 40.045 204.725 40.215 204.895 ;
        RECT 40.965 204.725 41.135 204.895 ;
        RECT 46.025 205.745 46.195 205.915 ;
        RECT 46.025 204.725 46.195 204.895 ;
        RECT 47.405 204.725 47.575 204.895 ;
        RECT 47.865 204.725 48.035 204.895 ;
        RECT 44.645 204.045 44.815 204.215 ;
        RECT 48.785 204.045 48.955 204.215 ;
        RECT 52.465 204.725 52.635 204.895 ;
        RECT 53.385 204.045 53.555 204.215 ;
        RECT 59.365 205.745 59.535 205.915 ;
        RECT 58.905 205.065 59.075 205.235 ;
        RECT 57.525 204.725 57.695 204.895 ;
        RECT 60.285 204.045 60.455 204.215 ;
        RECT 61.665 204.725 61.835 204.895 ;
        RECT 65.345 205.745 65.515 205.915 ;
        RECT 60.745 204.045 60.915 204.215 ;
        RECT 64.885 205.065 65.055 205.235 ;
        RECT 66.265 204.725 66.435 204.895 ;
        RECT 66.725 204.725 66.895 204.895 ;
        RECT 63.505 204.045 63.675 204.215 ;
        RECT 67.645 204.045 67.815 204.215 ;
        RECT 73.165 205.745 73.335 205.915 ;
        RECT 73.625 205.065 73.795 205.235 ;
        RECT 75.005 204.725 75.175 204.895 ;
        RECT 75.465 204.725 75.635 204.895 ;
        RECT 72.245 204.045 72.415 204.215 ;
        RECT 76.385 204.045 76.555 204.215 ;
        RECT 78.225 204.725 78.395 204.895 ;
        RECT 79.145 204.045 79.315 204.215 ;
        RECT 81.445 204.725 81.615 204.895 ;
        RECT 82.365 204.725 82.535 204.895 ;
        RECT 84.665 204.725 84.835 204.895 ;
        RECT 81.905 204.045 82.075 204.215 ;
        RECT 85.585 204.045 85.755 204.215 ;
        RECT 89.725 205.405 89.895 205.575 ;
        RECT 90.645 204.725 90.815 204.895 ;
        RECT 18.425 203.535 18.595 203.705 ;
        RECT 18.885 203.535 19.055 203.705 ;
        RECT 19.345 203.535 19.515 203.705 ;
        RECT 19.805 203.535 19.975 203.705 ;
        RECT 20.265 203.535 20.435 203.705 ;
        RECT 20.725 203.535 20.895 203.705 ;
        RECT 21.185 203.535 21.355 203.705 ;
        RECT 21.645 203.535 21.815 203.705 ;
        RECT 22.105 203.535 22.275 203.705 ;
        RECT 22.565 203.535 22.735 203.705 ;
        RECT 23.025 203.535 23.195 203.705 ;
        RECT 23.485 203.535 23.655 203.705 ;
        RECT 23.945 203.535 24.115 203.705 ;
        RECT 24.405 203.535 24.575 203.705 ;
        RECT 24.865 203.535 25.035 203.705 ;
        RECT 25.325 203.535 25.495 203.705 ;
        RECT 25.785 203.535 25.955 203.705 ;
        RECT 26.245 203.535 26.415 203.705 ;
        RECT 26.705 203.535 26.875 203.705 ;
        RECT 27.165 203.535 27.335 203.705 ;
        RECT 27.625 203.535 27.795 203.705 ;
        RECT 28.085 203.535 28.255 203.705 ;
        RECT 28.545 203.535 28.715 203.705 ;
        RECT 29.005 203.535 29.175 203.705 ;
        RECT 29.465 203.535 29.635 203.705 ;
        RECT 29.925 203.535 30.095 203.705 ;
        RECT 30.385 203.535 30.555 203.705 ;
        RECT 30.845 203.535 31.015 203.705 ;
        RECT 31.305 203.535 31.475 203.705 ;
        RECT 31.765 203.535 31.935 203.705 ;
        RECT 32.225 203.535 32.395 203.705 ;
        RECT 32.685 203.535 32.855 203.705 ;
        RECT 33.145 203.535 33.315 203.705 ;
        RECT 33.605 203.535 33.775 203.705 ;
        RECT 34.065 203.535 34.235 203.705 ;
        RECT 34.525 203.535 34.695 203.705 ;
        RECT 34.985 203.535 35.155 203.705 ;
        RECT 35.445 203.535 35.615 203.705 ;
        RECT 35.905 203.535 36.075 203.705 ;
        RECT 36.365 203.535 36.535 203.705 ;
        RECT 36.825 203.535 36.995 203.705 ;
        RECT 37.285 203.535 37.455 203.705 ;
        RECT 37.745 203.535 37.915 203.705 ;
        RECT 38.205 203.535 38.375 203.705 ;
        RECT 38.665 203.535 38.835 203.705 ;
        RECT 39.125 203.535 39.295 203.705 ;
        RECT 39.585 203.535 39.755 203.705 ;
        RECT 40.045 203.535 40.215 203.705 ;
        RECT 40.505 203.535 40.675 203.705 ;
        RECT 40.965 203.535 41.135 203.705 ;
        RECT 41.425 203.535 41.595 203.705 ;
        RECT 41.885 203.535 42.055 203.705 ;
        RECT 42.345 203.535 42.515 203.705 ;
        RECT 42.805 203.535 42.975 203.705 ;
        RECT 43.265 203.535 43.435 203.705 ;
        RECT 43.725 203.535 43.895 203.705 ;
        RECT 44.185 203.535 44.355 203.705 ;
        RECT 44.645 203.535 44.815 203.705 ;
        RECT 45.105 203.535 45.275 203.705 ;
        RECT 45.565 203.535 45.735 203.705 ;
        RECT 46.025 203.535 46.195 203.705 ;
        RECT 46.485 203.535 46.655 203.705 ;
        RECT 46.945 203.535 47.115 203.705 ;
        RECT 47.405 203.535 47.575 203.705 ;
        RECT 47.865 203.535 48.035 203.705 ;
        RECT 48.325 203.535 48.495 203.705 ;
        RECT 48.785 203.535 48.955 203.705 ;
        RECT 49.245 203.535 49.415 203.705 ;
        RECT 49.705 203.535 49.875 203.705 ;
        RECT 50.165 203.535 50.335 203.705 ;
        RECT 50.625 203.535 50.795 203.705 ;
        RECT 51.085 203.535 51.255 203.705 ;
        RECT 51.545 203.535 51.715 203.705 ;
        RECT 52.005 203.535 52.175 203.705 ;
        RECT 52.465 203.535 52.635 203.705 ;
        RECT 52.925 203.535 53.095 203.705 ;
        RECT 53.385 203.535 53.555 203.705 ;
        RECT 53.845 203.535 54.015 203.705 ;
        RECT 54.305 203.535 54.475 203.705 ;
        RECT 54.765 203.535 54.935 203.705 ;
        RECT 55.225 203.535 55.395 203.705 ;
        RECT 55.685 203.535 55.855 203.705 ;
        RECT 56.145 203.535 56.315 203.705 ;
        RECT 56.605 203.535 56.775 203.705 ;
        RECT 57.065 203.535 57.235 203.705 ;
        RECT 57.525 203.535 57.695 203.705 ;
        RECT 57.985 203.535 58.155 203.705 ;
        RECT 58.445 203.535 58.615 203.705 ;
        RECT 58.905 203.535 59.075 203.705 ;
        RECT 59.365 203.535 59.535 203.705 ;
        RECT 59.825 203.535 59.995 203.705 ;
        RECT 60.285 203.535 60.455 203.705 ;
        RECT 60.745 203.535 60.915 203.705 ;
        RECT 61.205 203.535 61.375 203.705 ;
        RECT 61.665 203.535 61.835 203.705 ;
        RECT 62.125 203.535 62.295 203.705 ;
        RECT 62.585 203.535 62.755 203.705 ;
        RECT 63.045 203.535 63.215 203.705 ;
        RECT 63.505 203.535 63.675 203.705 ;
        RECT 63.965 203.535 64.135 203.705 ;
        RECT 64.425 203.535 64.595 203.705 ;
        RECT 64.885 203.535 65.055 203.705 ;
        RECT 65.345 203.535 65.515 203.705 ;
        RECT 65.805 203.535 65.975 203.705 ;
        RECT 66.265 203.535 66.435 203.705 ;
        RECT 66.725 203.535 66.895 203.705 ;
        RECT 67.185 203.535 67.355 203.705 ;
        RECT 67.645 203.535 67.815 203.705 ;
        RECT 68.105 203.535 68.275 203.705 ;
        RECT 68.565 203.535 68.735 203.705 ;
        RECT 69.025 203.535 69.195 203.705 ;
        RECT 69.485 203.535 69.655 203.705 ;
        RECT 69.945 203.535 70.115 203.705 ;
        RECT 70.405 203.535 70.575 203.705 ;
        RECT 70.865 203.535 71.035 203.705 ;
        RECT 71.325 203.535 71.495 203.705 ;
        RECT 71.785 203.535 71.955 203.705 ;
        RECT 72.245 203.535 72.415 203.705 ;
        RECT 72.705 203.535 72.875 203.705 ;
        RECT 73.165 203.535 73.335 203.705 ;
        RECT 73.625 203.535 73.795 203.705 ;
        RECT 74.085 203.535 74.255 203.705 ;
        RECT 74.545 203.535 74.715 203.705 ;
        RECT 75.005 203.535 75.175 203.705 ;
        RECT 75.465 203.535 75.635 203.705 ;
        RECT 75.925 203.535 76.095 203.705 ;
        RECT 76.385 203.535 76.555 203.705 ;
        RECT 76.845 203.535 77.015 203.705 ;
        RECT 77.305 203.535 77.475 203.705 ;
        RECT 77.765 203.535 77.935 203.705 ;
        RECT 78.225 203.535 78.395 203.705 ;
        RECT 78.685 203.535 78.855 203.705 ;
        RECT 79.145 203.535 79.315 203.705 ;
        RECT 79.605 203.535 79.775 203.705 ;
        RECT 80.065 203.535 80.235 203.705 ;
        RECT 80.525 203.535 80.695 203.705 ;
        RECT 80.985 203.535 81.155 203.705 ;
        RECT 81.445 203.535 81.615 203.705 ;
        RECT 81.905 203.535 82.075 203.705 ;
        RECT 82.365 203.535 82.535 203.705 ;
        RECT 82.825 203.535 82.995 203.705 ;
        RECT 83.285 203.535 83.455 203.705 ;
        RECT 83.745 203.535 83.915 203.705 ;
        RECT 84.205 203.535 84.375 203.705 ;
        RECT 84.665 203.535 84.835 203.705 ;
        RECT 85.125 203.535 85.295 203.705 ;
        RECT 85.585 203.535 85.755 203.705 ;
        RECT 86.045 203.535 86.215 203.705 ;
        RECT 86.505 203.535 86.675 203.705 ;
        RECT 86.965 203.535 87.135 203.705 ;
        RECT 87.425 203.535 87.595 203.705 ;
        RECT 87.885 203.535 88.055 203.705 ;
        RECT 88.345 203.535 88.515 203.705 ;
        RECT 88.805 203.535 88.975 203.705 ;
        RECT 89.265 203.535 89.435 203.705 ;
        RECT 89.725 203.535 89.895 203.705 ;
        RECT 90.185 203.535 90.355 203.705 ;
        RECT 90.645 203.535 90.815 203.705 ;
        RECT 91.105 203.535 91.275 203.705 ;
        RECT 91.565 203.535 91.735 203.705 ;
        RECT 92.025 203.535 92.195 203.705 ;
        RECT 24.405 202.005 24.575 202.175 ;
        RECT 24.870 202.345 25.040 202.515 ;
        RECT 25.785 202.685 25.955 202.855 ;
        RECT 25.275 201.665 25.445 201.835 ;
        RECT 26.705 202.345 26.875 202.515 ;
        RECT 28.065 202.685 28.235 202.855 ;
        RECT 28.425 202.685 28.595 202.855 ;
        RECT 27.165 201.665 27.335 201.835 ;
        RECT 30.285 202.345 30.455 202.515 ;
        RECT 31.665 202.685 31.835 202.855 ;
        RECT 31.365 202.370 31.535 202.540 ;
        RECT 33.145 203.025 33.315 203.195 ;
        RECT 30.285 201.665 30.455 201.835 ;
        RECT 34.525 202.685 34.695 202.855 ;
        RECT 35.445 201.665 35.615 201.835 ;
        RECT 36.825 202.005 36.995 202.175 ;
        RECT 37.310 201.665 37.480 201.835 ;
        RECT 37.705 202.005 37.875 202.175 ;
        RECT 38.160 202.345 38.330 202.515 ;
        RECT 38.895 202.005 39.065 202.175 ;
        RECT 39.410 201.665 39.580 201.835 ;
        RECT 40.980 201.665 41.150 201.835 ;
        RECT 41.415 202.005 41.585 202.175 ;
        RECT 45.105 203.025 45.275 203.195 ;
        RECT 43.725 201.325 43.895 201.495 ;
        RECT 46.945 202.005 47.115 202.175 ;
        RECT 47.405 202.005 47.575 202.175 ;
        RECT 48.785 202.345 48.955 202.515 ;
        RECT 48.325 201.325 48.495 201.495 ;
        RECT 50.625 203.025 50.795 203.195 ;
        RECT 49.705 201.325 49.875 201.495 ;
        RECT 52.935 202.005 53.105 202.175 ;
        RECT 53.370 201.665 53.540 201.835 ;
        RECT 55.455 202.005 55.625 202.175 ;
        RECT 54.940 201.665 55.110 201.835 ;
        RECT 56.245 202.345 56.415 202.515 ;
        RECT 56.645 202.005 56.815 202.175 ;
        RECT 60.285 203.025 60.455 203.195 ;
        RECT 57.525 202.345 57.695 202.515 ;
        RECT 57.040 201.665 57.210 201.835 ;
        RECT 62.595 202.005 62.765 202.175 ;
        RECT 63.030 201.665 63.200 201.835 ;
        RECT 65.115 202.005 65.285 202.175 ;
        RECT 64.600 201.665 64.770 201.835 ;
        RECT 65.905 202.345 66.075 202.515 ;
        RECT 66.305 202.005 66.475 202.175 ;
        RECT 70.405 203.025 70.575 203.195 ;
        RECT 67.185 202.345 67.355 202.515 ;
        RECT 66.700 201.665 66.870 201.835 ;
        RECT 72.715 202.005 72.885 202.175 ;
        RECT 73.150 201.665 73.320 201.835 ;
        RECT 75.235 202.005 75.405 202.175 ;
        RECT 74.720 201.665 74.890 201.835 ;
        RECT 75.970 202.345 76.140 202.515 ;
        RECT 76.425 202.005 76.595 202.175 ;
        RECT 81.905 203.025 82.075 203.195 ;
        RECT 77.305 202.345 77.475 202.515 ;
        RECT 79.475 202.345 79.645 202.515 ;
        RECT 80.065 202.345 80.235 202.515 ;
        RECT 80.525 202.345 80.695 202.515 ;
        RECT 80.985 202.345 81.155 202.515 ;
        RECT 76.820 201.665 76.990 201.835 ;
        RECT 82.365 202.345 82.535 202.515 ;
        RECT 82.830 201.665 83.000 201.835 ;
        RECT 83.290 202.685 83.460 202.855 ;
        RECT 83.745 202.005 83.915 202.175 ;
        RECT 84.690 202.685 84.860 202.855 ;
        RECT 86.530 202.685 86.700 202.855 ;
        RECT 85.150 201.665 85.320 201.835 ;
        RECT 86.530 201.665 86.700 201.835 ;
        RECT 90.645 202.345 90.815 202.515 ;
        RECT 18.425 200.815 18.595 200.985 ;
        RECT 18.885 200.815 19.055 200.985 ;
        RECT 19.345 200.815 19.515 200.985 ;
        RECT 19.805 200.815 19.975 200.985 ;
        RECT 20.265 200.815 20.435 200.985 ;
        RECT 20.725 200.815 20.895 200.985 ;
        RECT 21.185 200.815 21.355 200.985 ;
        RECT 21.645 200.815 21.815 200.985 ;
        RECT 22.105 200.815 22.275 200.985 ;
        RECT 22.565 200.815 22.735 200.985 ;
        RECT 23.025 200.815 23.195 200.985 ;
        RECT 23.485 200.815 23.655 200.985 ;
        RECT 23.945 200.815 24.115 200.985 ;
        RECT 24.405 200.815 24.575 200.985 ;
        RECT 24.865 200.815 25.035 200.985 ;
        RECT 25.325 200.815 25.495 200.985 ;
        RECT 25.785 200.815 25.955 200.985 ;
        RECT 26.245 200.815 26.415 200.985 ;
        RECT 26.705 200.815 26.875 200.985 ;
        RECT 27.165 200.815 27.335 200.985 ;
        RECT 27.625 200.815 27.795 200.985 ;
        RECT 28.085 200.815 28.255 200.985 ;
        RECT 28.545 200.815 28.715 200.985 ;
        RECT 29.005 200.815 29.175 200.985 ;
        RECT 29.465 200.815 29.635 200.985 ;
        RECT 29.925 200.815 30.095 200.985 ;
        RECT 30.385 200.815 30.555 200.985 ;
        RECT 30.845 200.815 31.015 200.985 ;
        RECT 31.305 200.815 31.475 200.985 ;
        RECT 31.765 200.815 31.935 200.985 ;
        RECT 32.225 200.815 32.395 200.985 ;
        RECT 32.685 200.815 32.855 200.985 ;
        RECT 33.145 200.815 33.315 200.985 ;
        RECT 33.605 200.815 33.775 200.985 ;
        RECT 34.065 200.815 34.235 200.985 ;
        RECT 34.525 200.815 34.695 200.985 ;
        RECT 34.985 200.815 35.155 200.985 ;
        RECT 35.445 200.815 35.615 200.985 ;
        RECT 35.905 200.815 36.075 200.985 ;
        RECT 36.365 200.815 36.535 200.985 ;
        RECT 36.825 200.815 36.995 200.985 ;
        RECT 37.285 200.815 37.455 200.985 ;
        RECT 37.745 200.815 37.915 200.985 ;
        RECT 38.205 200.815 38.375 200.985 ;
        RECT 38.665 200.815 38.835 200.985 ;
        RECT 39.125 200.815 39.295 200.985 ;
        RECT 39.585 200.815 39.755 200.985 ;
        RECT 40.045 200.815 40.215 200.985 ;
        RECT 40.505 200.815 40.675 200.985 ;
        RECT 40.965 200.815 41.135 200.985 ;
        RECT 41.425 200.815 41.595 200.985 ;
        RECT 41.885 200.815 42.055 200.985 ;
        RECT 42.345 200.815 42.515 200.985 ;
        RECT 42.805 200.815 42.975 200.985 ;
        RECT 43.265 200.815 43.435 200.985 ;
        RECT 43.725 200.815 43.895 200.985 ;
        RECT 44.185 200.815 44.355 200.985 ;
        RECT 44.645 200.815 44.815 200.985 ;
        RECT 45.105 200.815 45.275 200.985 ;
        RECT 45.565 200.815 45.735 200.985 ;
        RECT 46.025 200.815 46.195 200.985 ;
        RECT 46.485 200.815 46.655 200.985 ;
        RECT 46.945 200.815 47.115 200.985 ;
        RECT 47.405 200.815 47.575 200.985 ;
        RECT 47.865 200.815 48.035 200.985 ;
        RECT 48.325 200.815 48.495 200.985 ;
        RECT 48.785 200.815 48.955 200.985 ;
        RECT 49.245 200.815 49.415 200.985 ;
        RECT 49.705 200.815 49.875 200.985 ;
        RECT 50.165 200.815 50.335 200.985 ;
        RECT 50.625 200.815 50.795 200.985 ;
        RECT 51.085 200.815 51.255 200.985 ;
        RECT 51.545 200.815 51.715 200.985 ;
        RECT 52.005 200.815 52.175 200.985 ;
        RECT 52.465 200.815 52.635 200.985 ;
        RECT 52.925 200.815 53.095 200.985 ;
        RECT 53.385 200.815 53.555 200.985 ;
        RECT 53.845 200.815 54.015 200.985 ;
        RECT 54.305 200.815 54.475 200.985 ;
        RECT 54.765 200.815 54.935 200.985 ;
        RECT 55.225 200.815 55.395 200.985 ;
        RECT 55.685 200.815 55.855 200.985 ;
        RECT 56.145 200.815 56.315 200.985 ;
        RECT 56.605 200.815 56.775 200.985 ;
        RECT 57.065 200.815 57.235 200.985 ;
        RECT 57.525 200.815 57.695 200.985 ;
        RECT 57.985 200.815 58.155 200.985 ;
        RECT 58.445 200.815 58.615 200.985 ;
        RECT 58.905 200.815 59.075 200.985 ;
        RECT 59.365 200.815 59.535 200.985 ;
        RECT 59.825 200.815 59.995 200.985 ;
        RECT 60.285 200.815 60.455 200.985 ;
        RECT 60.745 200.815 60.915 200.985 ;
        RECT 61.205 200.815 61.375 200.985 ;
        RECT 61.665 200.815 61.835 200.985 ;
        RECT 62.125 200.815 62.295 200.985 ;
        RECT 62.585 200.815 62.755 200.985 ;
        RECT 63.045 200.815 63.215 200.985 ;
        RECT 63.505 200.815 63.675 200.985 ;
        RECT 63.965 200.815 64.135 200.985 ;
        RECT 64.425 200.815 64.595 200.985 ;
        RECT 64.885 200.815 65.055 200.985 ;
        RECT 65.345 200.815 65.515 200.985 ;
        RECT 65.805 200.815 65.975 200.985 ;
        RECT 66.265 200.815 66.435 200.985 ;
        RECT 66.725 200.815 66.895 200.985 ;
        RECT 67.185 200.815 67.355 200.985 ;
        RECT 67.645 200.815 67.815 200.985 ;
        RECT 68.105 200.815 68.275 200.985 ;
        RECT 68.565 200.815 68.735 200.985 ;
        RECT 69.025 200.815 69.195 200.985 ;
        RECT 69.485 200.815 69.655 200.985 ;
        RECT 69.945 200.815 70.115 200.985 ;
        RECT 70.405 200.815 70.575 200.985 ;
        RECT 70.865 200.815 71.035 200.985 ;
        RECT 71.325 200.815 71.495 200.985 ;
        RECT 71.785 200.815 71.955 200.985 ;
        RECT 72.245 200.815 72.415 200.985 ;
        RECT 72.705 200.815 72.875 200.985 ;
        RECT 73.165 200.815 73.335 200.985 ;
        RECT 73.625 200.815 73.795 200.985 ;
        RECT 74.085 200.815 74.255 200.985 ;
        RECT 74.545 200.815 74.715 200.985 ;
        RECT 75.005 200.815 75.175 200.985 ;
        RECT 75.465 200.815 75.635 200.985 ;
        RECT 75.925 200.815 76.095 200.985 ;
        RECT 76.385 200.815 76.555 200.985 ;
        RECT 76.845 200.815 77.015 200.985 ;
        RECT 77.305 200.815 77.475 200.985 ;
        RECT 77.765 200.815 77.935 200.985 ;
        RECT 78.225 200.815 78.395 200.985 ;
        RECT 78.685 200.815 78.855 200.985 ;
        RECT 79.145 200.815 79.315 200.985 ;
        RECT 79.605 200.815 79.775 200.985 ;
        RECT 80.065 200.815 80.235 200.985 ;
        RECT 80.525 200.815 80.695 200.985 ;
        RECT 80.985 200.815 81.155 200.985 ;
        RECT 81.445 200.815 81.615 200.985 ;
        RECT 81.905 200.815 82.075 200.985 ;
        RECT 82.365 200.815 82.535 200.985 ;
        RECT 82.825 200.815 82.995 200.985 ;
        RECT 83.285 200.815 83.455 200.985 ;
        RECT 83.745 200.815 83.915 200.985 ;
        RECT 84.205 200.815 84.375 200.985 ;
        RECT 84.665 200.815 84.835 200.985 ;
        RECT 85.125 200.815 85.295 200.985 ;
        RECT 85.585 200.815 85.755 200.985 ;
        RECT 86.045 200.815 86.215 200.985 ;
        RECT 86.505 200.815 86.675 200.985 ;
        RECT 86.965 200.815 87.135 200.985 ;
        RECT 87.425 200.815 87.595 200.985 ;
        RECT 87.885 200.815 88.055 200.985 ;
        RECT 88.345 200.815 88.515 200.985 ;
        RECT 88.805 200.815 88.975 200.985 ;
        RECT 89.265 200.815 89.435 200.985 ;
        RECT 89.725 200.815 89.895 200.985 ;
        RECT 90.185 200.815 90.355 200.985 ;
        RECT 90.645 200.815 90.815 200.985 ;
        RECT 91.105 200.815 91.275 200.985 ;
        RECT 91.565 200.815 91.735 200.985 ;
        RECT 92.025 200.815 92.195 200.985 ;
        RECT 29.005 199.285 29.175 199.455 ;
        RECT 28.545 198.945 28.715 199.115 ;
        RECT 33.630 199.965 33.800 200.135 ;
        RECT 33.145 199.285 33.315 199.455 ;
        RECT 34.025 199.625 34.195 199.795 ;
        RECT 34.480 199.285 34.650 199.455 ;
        RECT 35.730 199.965 35.900 200.135 ;
        RECT 35.215 199.625 35.385 199.795 ;
        RECT 37.300 199.965 37.470 200.135 ;
        RECT 37.735 199.625 37.905 199.795 ;
        RECT 40.045 199.965 40.215 200.135 ;
        RECT 43.265 199.285 43.435 199.455 ;
        RECT 44.185 199.285 44.355 199.455 ;
        RECT 44.645 199.285 44.815 199.455 ;
        RECT 46.485 198.605 46.655 198.775 ;
        RECT 49.245 200.305 49.415 200.475 ;
        RECT 48.325 199.285 48.495 199.455 ;
        RECT 49.705 199.285 49.875 199.455 ;
        RECT 46.945 198.605 47.115 198.775 ;
        RECT 57.525 200.305 57.695 200.475 ;
        RECT 58.445 199.285 58.615 199.455 ;
        RECT 58.905 199.285 59.075 199.455 ;
        RECT 60.745 199.625 60.915 199.795 ;
        RECT 63.505 199.625 63.675 199.795 ;
        RECT 65.345 199.285 65.515 199.455 ;
        RECT 65.805 199.625 65.975 199.795 ;
        RECT 66.725 200.305 66.895 200.475 ;
        RECT 72.245 199.625 72.415 199.795 ;
        RECT 74.085 199.625 74.255 199.795 ;
        RECT 75.465 200.305 75.635 200.475 ;
        RECT 74.545 199.285 74.715 199.455 ;
        RECT 81.445 200.305 81.615 200.475 ;
        RECT 80.525 199.285 80.695 199.455 ;
        RECT 83.285 200.305 83.455 200.475 ;
        RECT 81.445 199.285 81.615 199.455 ;
        RECT 83.285 198.945 83.455 199.115 ;
        RECT 84.205 199.285 84.375 199.455 ;
        RECT 84.665 199.285 84.835 199.455 ;
        RECT 86.045 198.605 86.215 198.775 ;
        RECT 89.265 199.625 89.435 199.795 ;
        RECT 18.425 198.095 18.595 198.265 ;
        RECT 18.885 198.095 19.055 198.265 ;
        RECT 19.345 198.095 19.515 198.265 ;
        RECT 19.805 198.095 19.975 198.265 ;
        RECT 20.265 198.095 20.435 198.265 ;
        RECT 20.725 198.095 20.895 198.265 ;
        RECT 21.185 198.095 21.355 198.265 ;
        RECT 21.645 198.095 21.815 198.265 ;
        RECT 22.105 198.095 22.275 198.265 ;
        RECT 22.565 198.095 22.735 198.265 ;
        RECT 23.025 198.095 23.195 198.265 ;
        RECT 23.485 198.095 23.655 198.265 ;
        RECT 23.945 198.095 24.115 198.265 ;
        RECT 24.405 198.095 24.575 198.265 ;
        RECT 24.865 198.095 25.035 198.265 ;
        RECT 25.325 198.095 25.495 198.265 ;
        RECT 25.785 198.095 25.955 198.265 ;
        RECT 26.245 198.095 26.415 198.265 ;
        RECT 26.705 198.095 26.875 198.265 ;
        RECT 27.165 198.095 27.335 198.265 ;
        RECT 27.625 198.095 27.795 198.265 ;
        RECT 28.085 198.095 28.255 198.265 ;
        RECT 28.545 198.095 28.715 198.265 ;
        RECT 29.005 198.095 29.175 198.265 ;
        RECT 29.465 198.095 29.635 198.265 ;
        RECT 29.925 198.095 30.095 198.265 ;
        RECT 30.385 198.095 30.555 198.265 ;
        RECT 30.845 198.095 31.015 198.265 ;
        RECT 31.305 198.095 31.475 198.265 ;
        RECT 31.765 198.095 31.935 198.265 ;
        RECT 32.225 198.095 32.395 198.265 ;
        RECT 32.685 198.095 32.855 198.265 ;
        RECT 33.145 198.095 33.315 198.265 ;
        RECT 33.605 198.095 33.775 198.265 ;
        RECT 34.065 198.095 34.235 198.265 ;
        RECT 34.525 198.095 34.695 198.265 ;
        RECT 34.985 198.095 35.155 198.265 ;
        RECT 35.445 198.095 35.615 198.265 ;
        RECT 35.905 198.095 36.075 198.265 ;
        RECT 36.365 198.095 36.535 198.265 ;
        RECT 36.825 198.095 36.995 198.265 ;
        RECT 37.285 198.095 37.455 198.265 ;
        RECT 37.745 198.095 37.915 198.265 ;
        RECT 38.205 198.095 38.375 198.265 ;
        RECT 38.665 198.095 38.835 198.265 ;
        RECT 39.125 198.095 39.295 198.265 ;
        RECT 39.585 198.095 39.755 198.265 ;
        RECT 40.045 198.095 40.215 198.265 ;
        RECT 40.505 198.095 40.675 198.265 ;
        RECT 40.965 198.095 41.135 198.265 ;
        RECT 41.425 198.095 41.595 198.265 ;
        RECT 41.885 198.095 42.055 198.265 ;
        RECT 42.345 198.095 42.515 198.265 ;
        RECT 42.805 198.095 42.975 198.265 ;
        RECT 43.265 198.095 43.435 198.265 ;
        RECT 43.725 198.095 43.895 198.265 ;
        RECT 44.185 198.095 44.355 198.265 ;
        RECT 44.645 198.095 44.815 198.265 ;
        RECT 45.105 198.095 45.275 198.265 ;
        RECT 45.565 198.095 45.735 198.265 ;
        RECT 46.025 198.095 46.195 198.265 ;
        RECT 46.485 198.095 46.655 198.265 ;
        RECT 46.945 198.095 47.115 198.265 ;
        RECT 47.405 198.095 47.575 198.265 ;
        RECT 47.865 198.095 48.035 198.265 ;
        RECT 48.325 198.095 48.495 198.265 ;
        RECT 48.785 198.095 48.955 198.265 ;
        RECT 49.245 198.095 49.415 198.265 ;
        RECT 49.705 198.095 49.875 198.265 ;
        RECT 50.165 198.095 50.335 198.265 ;
        RECT 50.625 198.095 50.795 198.265 ;
        RECT 51.085 198.095 51.255 198.265 ;
        RECT 51.545 198.095 51.715 198.265 ;
        RECT 52.005 198.095 52.175 198.265 ;
        RECT 52.465 198.095 52.635 198.265 ;
        RECT 52.925 198.095 53.095 198.265 ;
        RECT 53.385 198.095 53.555 198.265 ;
        RECT 53.845 198.095 54.015 198.265 ;
        RECT 54.305 198.095 54.475 198.265 ;
        RECT 54.765 198.095 54.935 198.265 ;
        RECT 55.225 198.095 55.395 198.265 ;
        RECT 55.685 198.095 55.855 198.265 ;
        RECT 56.145 198.095 56.315 198.265 ;
        RECT 56.605 198.095 56.775 198.265 ;
        RECT 57.065 198.095 57.235 198.265 ;
        RECT 57.525 198.095 57.695 198.265 ;
        RECT 57.985 198.095 58.155 198.265 ;
        RECT 58.445 198.095 58.615 198.265 ;
        RECT 58.905 198.095 59.075 198.265 ;
        RECT 59.365 198.095 59.535 198.265 ;
        RECT 59.825 198.095 59.995 198.265 ;
        RECT 60.285 198.095 60.455 198.265 ;
        RECT 60.745 198.095 60.915 198.265 ;
        RECT 61.205 198.095 61.375 198.265 ;
        RECT 61.665 198.095 61.835 198.265 ;
        RECT 62.125 198.095 62.295 198.265 ;
        RECT 62.585 198.095 62.755 198.265 ;
        RECT 63.045 198.095 63.215 198.265 ;
        RECT 63.505 198.095 63.675 198.265 ;
        RECT 63.965 198.095 64.135 198.265 ;
        RECT 64.425 198.095 64.595 198.265 ;
        RECT 64.885 198.095 65.055 198.265 ;
        RECT 65.345 198.095 65.515 198.265 ;
        RECT 65.805 198.095 65.975 198.265 ;
        RECT 66.265 198.095 66.435 198.265 ;
        RECT 66.725 198.095 66.895 198.265 ;
        RECT 67.185 198.095 67.355 198.265 ;
        RECT 67.645 198.095 67.815 198.265 ;
        RECT 68.105 198.095 68.275 198.265 ;
        RECT 68.565 198.095 68.735 198.265 ;
        RECT 69.025 198.095 69.195 198.265 ;
        RECT 69.485 198.095 69.655 198.265 ;
        RECT 69.945 198.095 70.115 198.265 ;
        RECT 70.405 198.095 70.575 198.265 ;
        RECT 70.865 198.095 71.035 198.265 ;
        RECT 71.325 198.095 71.495 198.265 ;
        RECT 71.785 198.095 71.955 198.265 ;
        RECT 72.245 198.095 72.415 198.265 ;
        RECT 72.705 198.095 72.875 198.265 ;
        RECT 73.165 198.095 73.335 198.265 ;
        RECT 73.625 198.095 73.795 198.265 ;
        RECT 74.085 198.095 74.255 198.265 ;
        RECT 74.545 198.095 74.715 198.265 ;
        RECT 75.005 198.095 75.175 198.265 ;
        RECT 75.465 198.095 75.635 198.265 ;
        RECT 75.925 198.095 76.095 198.265 ;
        RECT 76.385 198.095 76.555 198.265 ;
        RECT 76.845 198.095 77.015 198.265 ;
        RECT 77.305 198.095 77.475 198.265 ;
        RECT 77.765 198.095 77.935 198.265 ;
        RECT 78.225 198.095 78.395 198.265 ;
        RECT 78.685 198.095 78.855 198.265 ;
        RECT 79.145 198.095 79.315 198.265 ;
        RECT 79.605 198.095 79.775 198.265 ;
        RECT 80.065 198.095 80.235 198.265 ;
        RECT 80.525 198.095 80.695 198.265 ;
        RECT 80.985 198.095 81.155 198.265 ;
        RECT 81.445 198.095 81.615 198.265 ;
        RECT 81.905 198.095 82.075 198.265 ;
        RECT 82.365 198.095 82.535 198.265 ;
        RECT 82.825 198.095 82.995 198.265 ;
        RECT 83.285 198.095 83.455 198.265 ;
        RECT 83.745 198.095 83.915 198.265 ;
        RECT 84.205 198.095 84.375 198.265 ;
        RECT 84.665 198.095 84.835 198.265 ;
        RECT 85.125 198.095 85.295 198.265 ;
        RECT 85.585 198.095 85.755 198.265 ;
        RECT 86.045 198.095 86.215 198.265 ;
        RECT 86.505 198.095 86.675 198.265 ;
        RECT 86.965 198.095 87.135 198.265 ;
        RECT 87.425 198.095 87.595 198.265 ;
        RECT 87.885 198.095 88.055 198.265 ;
        RECT 88.345 198.095 88.515 198.265 ;
        RECT 88.805 198.095 88.975 198.265 ;
        RECT 89.265 198.095 89.435 198.265 ;
        RECT 89.725 198.095 89.895 198.265 ;
        RECT 90.185 198.095 90.355 198.265 ;
        RECT 90.645 198.095 90.815 198.265 ;
        RECT 91.105 198.095 91.275 198.265 ;
        RECT 91.565 198.095 91.735 198.265 ;
        RECT 92.025 198.095 92.195 198.265 ;
        RECT 47.865 196.905 48.035 197.075 ;
        RECT 48.325 195.885 48.495 196.055 ;
        RECT 53.385 195.885 53.555 196.055 ;
        RECT 54.305 196.565 54.475 196.735 ;
        RECT 54.765 196.905 54.935 197.075 ;
        RECT 56.605 197.585 56.775 197.755 ;
        RECT 57.065 197.585 57.235 197.755 ;
        RECT 59.825 196.905 59.995 197.075 ;
        RECT 58.445 196.565 58.615 196.735 ;
        RECT 59.365 195.885 59.535 196.055 ;
        RECT 64.885 196.905 65.055 197.075 ;
        RECT 63.965 195.885 64.135 196.055 ;
        RECT 65.345 196.905 65.515 197.075 ;
        RECT 67.185 196.565 67.355 196.735 ;
        RECT 71.785 196.565 71.955 196.735 ;
        RECT 73.625 196.905 73.795 197.075 ;
        RECT 74.085 196.565 74.255 196.735 ;
        RECT 81.445 197.585 81.615 197.755 ;
        RECT 75.005 195.885 75.175 196.055 ;
        RECT 81.905 196.905 82.075 197.075 ;
        RECT 80.525 195.885 80.695 196.055 ;
        RECT 81.445 196.565 81.615 196.735 ;
        RECT 82.825 196.905 82.995 197.075 ;
        RECT 83.285 196.905 83.455 197.075 ;
        RECT 83.745 196.905 83.915 197.075 ;
        RECT 85.585 196.905 85.755 197.075 ;
        RECT 86.505 196.905 86.675 197.075 ;
        RECT 85.125 195.885 85.295 196.055 ;
        RECT 87.425 195.885 87.595 196.055 ;
        RECT 18.425 195.375 18.595 195.545 ;
        RECT 18.885 195.375 19.055 195.545 ;
        RECT 19.345 195.375 19.515 195.545 ;
        RECT 19.805 195.375 19.975 195.545 ;
        RECT 20.265 195.375 20.435 195.545 ;
        RECT 20.725 195.375 20.895 195.545 ;
        RECT 21.185 195.375 21.355 195.545 ;
        RECT 21.645 195.375 21.815 195.545 ;
        RECT 22.105 195.375 22.275 195.545 ;
        RECT 22.565 195.375 22.735 195.545 ;
        RECT 23.025 195.375 23.195 195.545 ;
        RECT 23.485 195.375 23.655 195.545 ;
        RECT 23.945 195.375 24.115 195.545 ;
        RECT 24.405 195.375 24.575 195.545 ;
        RECT 24.865 195.375 25.035 195.545 ;
        RECT 25.325 195.375 25.495 195.545 ;
        RECT 25.785 195.375 25.955 195.545 ;
        RECT 26.245 195.375 26.415 195.545 ;
        RECT 26.705 195.375 26.875 195.545 ;
        RECT 27.165 195.375 27.335 195.545 ;
        RECT 27.625 195.375 27.795 195.545 ;
        RECT 28.085 195.375 28.255 195.545 ;
        RECT 28.545 195.375 28.715 195.545 ;
        RECT 29.005 195.375 29.175 195.545 ;
        RECT 29.465 195.375 29.635 195.545 ;
        RECT 29.925 195.375 30.095 195.545 ;
        RECT 30.385 195.375 30.555 195.545 ;
        RECT 30.845 195.375 31.015 195.545 ;
        RECT 31.305 195.375 31.475 195.545 ;
        RECT 31.765 195.375 31.935 195.545 ;
        RECT 32.225 195.375 32.395 195.545 ;
        RECT 32.685 195.375 32.855 195.545 ;
        RECT 33.145 195.375 33.315 195.545 ;
        RECT 33.605 195.375 33.775 195.545 ;
        RECT 34.065 195.375 34.235 195.545 ;
        RECT 34.525 195.375 34.695 195.545 ;
        RECT 34.985 195.375 35.155 195.545 ;
        RECT 35.445 195.375 35.615 195.545 ;
        RECT 35.905 195.375 36.075 195.545 ;
        RECT 36.365 195.375 36.535 195.545 ;
        RECT 36.825 195.375 36.995 195.545 ;
        RECT 37.285 195.375 37.455 195.545 ;
        RECT 37.745 195.375 37.915 195.545 ;
        RECT 38.205 195.375 38.375 195.545 ;
        RECT 38.665 195.375 38.835 195.545 ;
        RECT 39.125 195.375 39.295 195.545 ;
        RECT 39.585 195.375 39.755 195.545 ;
        RECT 40.045 195.375 40.215 195.545 ;
        RECT 40.505 195.375 40.675 195.545 ;
        RECT 40.965 195.375 41.135 195.545 ;
        RECT 41.425 195.375 41.595 195.545 ;
        RECT 41.885 195.375 42.055 195.545 ;
        RECT 42.345 195.375 42.515 195.545 ;
        RECT 42.805 195.375 42.975 195.545 ;
        RECT 43.265 195.375 43.435 195.545 ;
        RECT 43.725 195.375 43.895 195.545 ;
        RECT 44.185 195.375 44.355 195.545 ;
        RECT 44.645 195.375 44.815 195.545 ;
        RECT 45.105 195.375 45.275 195.545 ;
        RECT 45.565 195.375 45.735 195.545 ;
        RECT 46.025 195.375 46.195 195.545 ;
        RECT 46.485 195.375 46.655 195.545 ;
        RECT 46.945 195.375 47.115 195.545 ;
        RECT 47.405 195.375 47.575 195.545 ;
        RECT 47.865 195.375 48.035 195.545 ;
        RECT 48.325 195.375 48.495 195.545 ;
        RECT 48.785 195.375 48.955 195.545 ;
        RECT 49.245 195.375 49.415 195.545 ;
        RECT 49.705 195.375 49.875 195.545 ;
        RECT 50.165 195.375 50.335 195.545 ;
        RECT 50.625 195.375 50.795 195.545 ;
        RECT 51.085 195.375 51.255 195.545 ;
        RECT 51.545 195.375 51.715 195.545 ;
        RECT 52.005 195.375 52.175 195.545 ;
        RECT 52.465 195.375 52.635 195.545 ;
        RECT 52.925 195.375 53.095 195.545 ;
        RECT 53.385 195.375 53.555 195.545 ;
        RECT 53.845 195.375 54.015 195.545 ;
        RECT 54.305 195.375 54.475 195.545 ;
        RECT 54.765 195.375 54.935 195.545 ;
        RECT 55.225 195.375 55.395 195.545 ;
        RECT 55.685 195.375 55.855 195.545 ;
        RECT 56.145 195.375 56.315 195.545 ;
        RECT 56.605 195.375 56.775 195.545 ;
        RECT 57.065 195.375 57.235 195.545 ;
        RECT 57.525 195.375 57.695 195.545 ;
        RECT 57.985 195.375 58.155 195.545 ;
        RECT 58.445 195.375 58.615 195.545 ;
        RECT 58.905 195.375 59.075 195.545 ;
        RECT 59.365 195.375 59.535 195.545 ;
        RECT 59.825 195.375 59.995 195.545 ;
        RECT 60.285 195.375 60.455 195.545 ;
        RECT 60.745 195.375 60.915 195.545 ;
        RECT 61.205 195.375 61.375 195.545 ;
        RECT 61.665 195.375 61.835 195.545 ;
        RECT 62.125 195.375 62.295 195.545 ;
        RECT 62.585 195.375 62.755 195.545 ;
        RECT 63.045 195.375 63.215 195.545 ;
        RECT 63.505 195.375 63.675 195.545 ;
        RECT 63.965 195.375 64.135 195.545 ;
        RECT 64.425 195.375 64.595 195.545 ;
        RECT 64.885 195.375 65.055 195.545 ;
        RECT 65.345 195.375 65.515 195.545 ;
        RECT 65.805 195.375 65.975 195.545 ;
        RECT 66.265 195.375 66.435 195.545 ;
        RECT 66.725 195.375 66.895 195.545 ;
        RECT 67.185 195.375 67.355 195.545 ;
        RECT 67.645 195.375 67.815 195.545 ;
        RECT 68.105 195.375 68.275 195.545 ;
        RECT 68.565 195.375 68.735 195.545 ;
        RECT 69.025 195.375 69.195 195.545 ;
        RECT 69.485 195.375 69.655 195.545 ;
        RECT 69.945 195.375 70.115 195.545 ;
        RECT 70.405 195.375 70.575 195.545 ;
        RECT 70.865 195.375 71.035 195.545 ;
        RECT 71.325 195.375 71.495 195.545 ;
        RECT 71.785 195.375 71.955 195.545 ;
        RECT 72.245 195.375 72.415 195.545 ;
        RECT 72.705 195.375 72.875 195.545 ;
        RECT 73.165 195.375 73.335 195.545 ;
        RECT 73.625 195.375 73.795 195.545 ;
        RECT 74.085 195.375 74.255 195.545 ;
        RECT 74.545 195.375 74.715 195.545 ;
        RECT 75.005 195.375 75.175 195.545 ;
        RECT 75.465 195.375 75.635 195.545 ;
        RECT 75.925 195.375 76.095 195.545 ;
        RECT 76.385 195.375 76.555 195.545 ;
        RECT 76.845 195.375 77.015 195.545 ;
        RECT 77.305 195.375 77.475 195.545 ;
        RECT 77.765 195.375 77.935 195.545 ;
        RECT 78.225 195.375 78.395 195.545 ;
        RECT 78.685 195.375 78.855 195.545 ;
        RECT 79.145 195.375 79.315 195.545 ;
        RECT 79.605 195.375 79.775 195.545 ;
        RECT 80.065 195.375 80.235 195.545 ;
        RECT 80.525 195.375 80.695 195.545 ;
        RECT 80.985 195.375 81.155 195.545 ;
        RECT 81.445 195.375 81.615 195.545 ;
        RECT 81.905 195.375 82.075 195.545 ;
        RECT 82.365 195.375 82.535 195.545 ;
        RECT 82.825 195.375 82.995 195.545 ;
        RECT 83.285 195.375 83.455 195.545 ;
        RECT 83.745 195.375 83.915 195.545 ;
        RECT 84.205 195.375 84.375 195.545 ;
        RECT 84.665 195.375 84.835 195.545 ;
        RECT 85.125 195.375 85.295 195.545 ;
        RECT 85.585 195.375 85.755 195.545 ;
        RECT 86.045 195.375 86.215 195.545 ;
        RECT 86.505 195.375 86.675 195.545 ;
        RECT 86.965 195.375 87.135 195.545 ;
        RECT 87.425 195.375 87.595 195.545 ;
        RECT 87.885 195.375 88.055 195.545 ;
        RECT 88.345 195.375 88.515 195.545 ;
        RECT 88.805 195.375 88.975 195.545 ;
        RECT 89.265 195.375 89.435 195.545 ;
        RECT 89.725 195.375 89.895 195.545 ;
        RECT 90.185 195.375 90.355 195.545 ;
        RECT 90.645 195.375 90.815 195.545 ;
        RECT 91.105 195.375 91.275 195.545 ;
        RECT 91.565 195.375 91.735 195.545 ;
        RECT 92.025 195.375 92.195 195.545 ;
        RECT 33.170 194.525 33.340 194.695 ;
        RECT 32.685 193.845 32.855 194.015 ;
        RECT 33.565 194.185 33.735 194.355 ;
        RECT 34.020 193.505 34.190 193.675 ;
        RECT 35.270 194.525 35.440 194.695 ;
        RECT 34.755 194.185 34.925 194.355 ;
        RECT 36.840 194.525 37.010 194.695 ;
        RECT 37.275 194.185 37.445 194.355 ;
        RECT 43.265 194.865 43.435 195.035 ;
        RECT 41.885 193.845 42.055 194.015 ;
        RECT 39.585 193.165 39.755 193.335 ;
        RECT 44.645 193.845 44.815 194.015 ;
        RECT 46.025 194.525 46.195 194.695 ;
        RECT 44.185 193.165 44.355 193.335 ;
        RECT 46.945 193.165 47.115 193.335 ;
        RECT 48.325 193.165 48.495 193.335 ;
        RECT 50.635 194.185 50.805 194.355 ;
        RECT 51.070 194.525 51.240 194.695 ;
        RECT 52.640 194.525 52.810 194.695 ;
        RECT 53.155 194.185 53.325 194.355 ;
        RECT 53.890 193.845 54.060 194.015 ;
        RECT 54.345 194.185 54.515 194.355 ;
        RECT 54.740 194.525 54.910 194.695 ;
        RECT 55.225 194.185 55.395 194.355 ;
        RECT 59.825 193.845 59.995 194.015 ;
        RECT 59.365 193.165 59.535 193.335 ;
        RECT 60.285 193.165 60.455 193.335 ;
        RECT 62.595 194.185 62.765 194.355 ;
        RECT 63.030 194.525 63.200 194.695 ;
        RECT 64.600 194.525 64.770 194.695 ;
        RECT 65.115 194.185 65.285 194.355 ;
        RECT 65.850 193.505 66.020 193.675 ;
        RECT 66.305 194.185 66.475 194.355 ;
        RECT 66.700 194.525 66.870 194.695 ;
        RECT 67.185 194.185 67.355 194.355 ;
        RECT 69.485 193.165 69.655 193.335 ;
        RECT 71.795 194.185 71.965 194.355 ;
        RECT 72.230 194.525 72.400 194.695 ;
        RECT 73.800 194.525 73.970 194.695 ;
        RECT 74.315 194.185 74.485 194.355 ;
        RECT 75.050 193.505 75.220 193.675 ;
        RECT 75.505 194.185 75.675 194.355 ;
        RECT 75.900 194.525 76.070 194.695 ;
        RECT 76.385 193.845 76.555 194.015 ;
        RECT 79.145 193.845 79.315 194.015 ;
        RECT 80.065 193.165 80.235 193.335 ;
        RECT 80.525 194.865 80.695 195.035 ;
        RECT 83.285 194.865 83.455 195.035 ;
        RECT 81.445 193.845 81.615 194.015 ;
        RECT 82.365 193.845 82.535 194.015 ;
        RECT 84.205 193.845 84.375 194.015 ;
        RECT 84.665 193.505 84.835 193.675 ;
        RECT 85.125 193.845 85.295 194.015 ;
        RECT 86.045 193.845 86.215 194.015 ;
        RECT 86.505 193.895 86.675 194.065 ;
        RECT 86.995 193.845 87.165 194.015 ;
        RECT 87.885 193.845 88.055 194.015 ;
        RECT 87.425 193.165 87.595 193.335 ;
        RECT 18.425 192.655 18.595 192.825 ;
        RECT 18.885 192.655 19.055 192.825 ;
        RECT 19.345 192.655 19.515 192.825 ;
        RECT 19.805 192.655 19.975 192.825 ;
        RECT 20.265 192.655 20.435 192.825 ;
        RECT 20.725 192.655 20.895 192.825 ;
        RECT 21.185 192.655 21.355 192.825 ;
        RECT 21.645 192.655 21.815 192.825 ;
        RECT 22.105 192.655 22.275 192.825 ;
        RECT 22.565 192.655 22.735 192.825 ;
        RECT 23.025 192.655 23.195 192.825 ;
        RECT 23.485 192.655 23.655 192.825 ;
        RECT 23.945 192.655 24.115 192.825 ;
        RECT 24.405 192.655 24.575 192.825 ;
        RECT 24.865 192.655 25.035 192.825 ;
        RECT 25.325 192.655 25.495 192.825 ;
        RECT 25.785 192.655 25.955 192.825 ;
        RECT 26.245 192.655 26.415 192.825 ;
        RECT 26.705 192.655 26.875 192.825 ;
        RECT 27.165 192.655 27.335 192.825 ;
        RECT 27.625 192.655 27.795 192.825 ;
        RECT 28.085 192.655 28.255 192.825 ;
        RECT 28.545 192.655 28.715 192.825 ;
        RECT 29.005 192.655 29.175 192.825 ;
        RECT 29.465 192.655 29.635 192.825 ;
        RECT 29.925 192.655 30.095 192.825 ;
        RECT 30.385 192.655 30.555 192.825 ;
        RECT 30.845 192.655 31.015 192.825 ;
        RECT 31.305 192.655 31.475 192.825 ;
        RECT 31.765 192.655 31.935 192.825 ;
        RECT 32.225 192.655 32.395 192.825 ;
        RECT 32.685 192.655 32.855 192.825 ;
        RECT 33.145 192.655 33.315 192.825 ;
        RECT 33.605 192.655 33.775 192.825 ;
        RECT 34.065 192.655 34.235 192.825 ;
        RECT 34.525 192.655 34.695 192.825 ;
        RECT 34.985 192.655 35.155 192.825 ;
        RECT 35.445 192.655 35.615 192.825 ;
        RECT 35.905 192.655 36.075 192.825 ;
        RECT 36.365 192.655 36.535 192.825 ;
        RECT 36.825 192.655 36.995 192.825 ;
        RECT 37.285 192.655 37.455 192.825 ;
        RECT 37.745 192.655 37.915 192.825 ;
        RECT 38.205 192.655 38.375 192.825 ;
        RECT 38.665 192.655 38.835 192.825 ;
        RECT 39.125 192.655 39.295 192.825 ;
        RECT 39.585 192.655 39.755 192.825 ;
        RECT 40.045 192.655 40.215 192.825 ;
        RECT 40.505 192.655 40.675 192.825 ;
        RECT 40.965 192.655 41.135 192.825 ;
        RECT 41.425 192.655 41.595 192.825 ;
        RECT 41.885 192.655 42.055 192.825 ;
        RECT 42.345 192.655 42.515 192.825 ;
        RECT 42.805 192.655 42.975 192.825 ;
        RECT 43.265 192.655 43.435 192.825 ;
        RECT 43.725 192.655 43.895 192.825 ;
        RECT 44.185 192.655 44.355 192.825 ;
        RECT 44.645 192.655 44.815 192.825 ;
        RECT 45.105 192.655 45.275 192.825 ;
        RECT 45.565 192.655 45.735 192.825 ;
        RECT 46.025 192.655 46.195 192.825 ;
        RECT 46.485 192.655 46.655 192.825 ;
        RECT 46.945 192.655 47.115 192.825 ;
        RECT 47.405 192.655 47.575 192.825 ;
        RECT 47.865 192.655 48.035 192.825 ;
        RECT 48.325 192.655 48.495 192.825 ;
        RECT 48.785 192.655 48.955 192.825 ;
        RECT 49.245 192.655 49.415 192.825 ;
        RECT 49.705 192.655 49.875 192.825 ;
        RECT 50.165 192.655 50.335 192.825 ;
        RECT 50.625 192.655 50.795 192.825 ;
        RECT 51.085 192.655 51.255 192.825 ;
        RECT 51.545 192.655 51.715 192.825 ;
        RECT 52.005 192.655 52.175 192.825 ;
        RECT 52.465 192.655 52.635 192.825 ;
        RECT 52.925 192.655 53.095 192.825 ;
        RECT 53.385 192.655 53.555 192.825 ;
        RECT 53.845 192.655 54.015 192.825 ;
        RECT 54.305 192.655 54.475 192.825 ;
        RECT 54.765 192.655 54.935 192.825 ;
        RECT 55.225 192.655 55.395 192.825 ;
        RECT 55.685 192.655 55.855 192.825 ;
        RECT 56.145 192.655 56.315 192.825 ;
        RECT 56.605 192.655 56.775 192.825 ;
        RECT 57.065 192.655 57.235 192.825 ;
        RECT 57.525 192.655 57.695 192.825 ;
        RECT 57.985 192.655 58.155 192.825 ;
        RECT 58.445 192.655 58.615 192.825 ;
        RECT 58.905 192.655 59.075 192.825 ;
        RECT 59.365 192.655 59.535 192.825 ;
        RECT 59.825 192.655 59.995 192.825 ;
        RECT 60.285 192.655 60.455 192.825 ;
        RECT 60.745 192.655 60.915 192.825 ;
        RECT 61.205 192.655 61.375 192.825 ;
        RECT 61.665 192.655 61.835 192.825 ;
        RECT 62.125 192.655 62.295 192.825 ;
        RECT 62.585 192.655 62.755 192.825 ;
        RECT 63.045 192.655 63.215 192.825 ;
        RECT 63.505 192.655 63.675 192.825 ;
        RECT 63.965 192.655 64.135 192.825 ;
        RECT 64.425 192.655 64.595 192.825 ;
        RECT 64.885 192.655 65.055 192.825 ;
        RECT 65.345 192.655 65.515 192.825 ;
        RECT 65.805 192.655 65.975 192.825 ;
        RECT 66.265 192.655 66.435 192.825 ;
        RECT 66.725 192.655 66.895 192.825 ;
        RECT 67.185 192.655 67.355 192.825 ;
        RECT 67.645 192.655 67.815 192.825 ;
        RECT 68.105 192.655 68.275 192.825 ;
        RECT 68.565 192.655 68.735 192.825 ;
        RECT 69.025 192.655 69.195 192.825 ;
        RECT 69.485 192.655 69.655 192.825 ;
        RECT 69.945 192.655 70.115 192.825 ;
        RECT 70.405 192.655 70.575 192.825 ;
        RECT 70.865 192.655 71.035 192.825 ;
        RECT 71.325 192.655 71.495 192.825 ;
        RECT 71.785 192.655 71.955 192.825 ;
        RECT 72.245 192.655 72.415 192.825 ;
        RECT 72.705 192.655 72.875 192.825 ;
        RECT 73.165 192.655 73.335 192.825 ;
        RECT 73.625 192.655 73.795 192.825 ;
        RECT 74.085 192.655 74.255 192.825 ;
        RECT 74.545 192.655 74.715 192.825 ;
        RECT 75.005 192.655 75.175 192.825 ;
        RECT 75.465 192.655 75.635 192.825 ;
        RECT 75.925 192.655 76.095 192.825 ;
        RECT 76.385 192.655 76.555 192.825 ;
        RECT 76.845 192.655 77.015 192.825 ;
        RECT 77.305 192.655 77.475 192.825 ;
        RECT 77.765 192.655 77.935 192.825 ;
        RECT 78.225 192.655 78.395 192.825 ;
        RECT 78.685 192.655 78.855 192.825 ;
        RECT 79.145 192.655 79.315 192.825 ;
        RECT 79.605 192.655 79.775 192.825 ;
        RECT 80.065 192.655 80.235 192.825 ;
        RECT 80.525 192.655 80.695 192.825 ;
        RECT 80.985 192.655 81.155 192.825 ;
        RECT 81.445 192.655 81.615 192.825 ;
        RECT 81.905 192.655 82.075 192.825 ;
        RECT 82.365 192.655 82.535 192.825 ;
        RECT 82.825 192.655 82.995 192.825 ;
        RECT 83.285 192.655 83.455 192.825 ;
        RECT 83.745 192.655 83.915 192.825 ;
        RECT 84.205 192.655 84.375 192.825 ;
        RECT 84.665 192.655 84.835 192.825 ;
        RECT 85.125 192.655 85.295 192.825 ;
        RECT 85.585 192.655 85.755 192.825 ;
        RECT 86.045 192.655 86.215 192.825 ;
        RECT 86.505 192.655 86.675 192.825 ;
        RECT 86.965 192.655 87.135 192.825 ;
        RECT 87.425 192.655 87.595 192.825 ;
        RECT 87.885 192.655 88.055 192.825 ;
        RECT 88.345 192.655 88.515 192.825 ;
        RECT 88.805 192.655 88.975 192.825 ;
        RECT 89.265 192.655 89.435 192.825 ;
        RECT 89.725 192.655 89.895 192.825 ;
        RECT 90.185 192.655 90.355 192.825 ;
        RECT 90.645 192.655 90.815 192.825 ;
        RECT 91.105 192.655 91.275 192.825 ;
        RECT 91.565 192.655 91.735 192.825 ;
        RECT 92.025 192.655 92.195 192.825 ;
        RECT 26.245 191.125 26.415 191.295 ;
        RECT 26.730 190.785 26.900 190.955 ;
        RECT 27.125 191.125 27.295 191.295 ;
        RECT 27.580 191.805 27.750 191.975 ;
        RECT 28.315 191.125 28.485 191.295 ;
        RECT 28.830 190.785 29.000 190.955 ;
        RECT 30.400 190.785 30.570 190.955 ;
        RECT 30.835 191.125 31.005 191.295 ;
        RECT 34.525 191.805 34.695 191.975 ;
        RECT 34.065 191.465 34.235 191.635 ;
        RECT 34.985 191.465 35.155 191.635 ;
        RECT 33.145 190.785 33.315 190.955 ;
        RECT 36.825 191.465 36.995 191.635 ;
        RECT 37.285 190.785 37.455 190.955 ;
        RECT 40.045 191.125 40.215 191.295 ;
        RECT 46.485 191.805 46.655 191.975 ;
        RECT 45.105 191.465 45.275 191.635 ;
        RECT 46.945 191.465 47.115 191.635 ;
        RECT 47.635 191.465 47.805 191.635 ;
        RECT 43.265 190.445 43.435 190.615 ;
        RECT 51.545 191.465 51.715 191.635 ;
        RECT 52.925 191.465 53.095 191.635 ;
        RECT 53.385 191.465 53.555 191.635 ;
        RECT 48.325 190.445 48.495 190.615 ;
        RECT 52.005 190.445 52.175 190.615 ;
        RECT 64.885 192.145 65.055 192.315 ;
        RECT 54.305 190.445 54.475 190.615 ;
        RECT 63.045 191.465 63.215 191.635 ;
        RECT 63.505 191.125 63.675 191.295 ;
        RECT 71.325 192.145 71.495 192.315 ;
        RECT 63.045 190.445 63.215 190.615 ;
        RECT 74.085 191.465 74.255 191.635 ;
        RECT 72.705 191.125 72.875 191.295 ;
        RECT 72.705 190.445 72.875 190.615 ;
        RECT 82.365 191.465 82.535 191.635 ;
        RECT 82.830 190.785 83.000 190.955 ;
        RECT 83.290 191.805 83.460 191.975 ;
        RECT 83.745 191.465 83.915 191.635 ;
        RECT 84.690 191.805 84.860 191.975 ;
        RECT 86.530 191.805 86.700 191.975 ;
        RECT 85.150 190.785 85.320 190.955 ;
        RECT 86.530 190.785 86.700 190.955 ;
        RECT 90.645 191.805 90.815 191.975 ;
        RECT 18.425 189.935 18.595 190.105 ;
        RECT 18.885 189.935 19.055 190.105 ;
        RECT 19.345 189.935 19.515 190.105 ;
        RECT 19.805 189.935 19.975 190.105 ;
        RECT 20.265 189.935 20.435 190.105 ;
        RECT 20.725 189.935 20.895 190.105 ;
        RECT 21.185 189.935 21.355 190.105 ;
        RECT 21.645 189.935 21.815 190.105 ;
        RECT 22.105 189.935 22.275 190.105 ;
        RECT 22.565 189.935 22.735 190.105 ;
        RECT 23.025 189.935 23.195 190.105 ;
        RECT 23.485 189.935 23.655 190.105 ;
        RECT 23.945 189.935 24.115 190.105 ;
        RECT 24.405 189.935 24.575 190.105 ;
        RECT 24.865 189.935 25.035 190.105 ;
        RECT 25.325 189.935 25.495 190.105 ;
        RECT 25.785 189.935 25.955 190.105 ;
        RECT 26.245 189.935 26.415 190.105 ;
        RECT 26.705 189.935 26.875 190.105 ;
        RECT 27.165 189.935 27.335 190.105 ;
        RECT 27.625 189.935 27.795 190.105 ;
        RECT 28.085 189.935 28.255 190.105 ;
        RECT 28.545 189.935 28.715 190.105 ;
        RECT 29.005 189.935 29.175 190.105 ;
        RECT 29.465 189.935 29.635 190.105 ;
        RECT 29.925 189.935 30.095 190.105 ;
        RECT 30.385 189.935 30.555 190.105 ;
        RECT 30.845 189.935 31.015 190.105 ;
        RECT 31.305 189.935 31.475 190.105 ;
        RECT 31.765 189.935 31.935 190.105 ;
        RECT 32.225 189.935 32.395 190.105 ;
        RECT 32.685 189.935 32.855 190.105 ;
        RECT 33.145 189.935 33.315 190.105 ;
        RECT 33.605 189.935 33.775 190.105 ;
        RECT 34.065 189.935 34.235 190.105 ;
        RECT 34.525 189.935 34.695 190.105 ;
        RECT 34.985 189.935 35.155 190.105 ;
        RECT 35.445 189.935 35.615 190.105 ;
        RECT 35.905 189.935 36.075 190.105 ;
        RECT 36.365 189.935 36.535 190.105 ;
        RECT 36.825 189.935 36.995 190.105 ;
        RECT 37.285 189.935 37.455 190.105 ;
        RECT 37.745 189.935 37.915 190.105 ;
        RECT 38.205 189.935 38.375 190.105 ;
        RECT 38.665 189.935 38.835 190.105 ;
        RECT 39.125 189.935 39.295 190.105 ;
        RECT 39.585 189.935 39.755 190.105 ;
        RECT 40.045 189.935 40.215 190.105 ;
        RECT 40.505 189.935 40.675 190.105 ;
        RECT 40.965 189.935 41.135 190.105 ;
        RECT 41.425 189.935 41.595 190.105 ;
        RECT 41.885 189.935 42.055 190.105 ;
        RECT 42.345 189.935 42.515 190.105 ;
        RECT 42.805 189.935 42.975 190.105 ;
        RECT 43.265 189.935 43.435 190.105 ;
        RECT 43.725 189.935 43.895 190.105 ;
        RECT 44.185 189.935 44.355 190.105 ;
        RECT 44.645 189.935 44.815 190.105 ;
        RECT 45.105 189.935 45.275 190.105 ;
        RECT 45.565 189.935 45.735 190.105 ;
        RECT 46.025 189.935 46.195 190.105 ;
        RECT 46.485 189.935 46.655 190.105 ;
        RECT 46.945 189.935 47.115 190.105 ;
        RECT 47.405 189.935 47.575 190.105 ;
        RECT 47.865 189.935 48.035 190.105 ;
        RECT 48.325 189.935 48.495 190.105 ;
        RECT 48.785 189.935 48.955 190.105 ;
        RECT 49.245 189.935 49.415 190.105 ;
        RECT 49.705 189.935 49.875 190.105 ;
        RECT 50.165 189.935 50.335 190.105 ;
        RECT 50.625 189.935 50.795 190.105 ;
        RECT 51.085 189.935 51.255 190.105 ;
        RECT 51.545 189.935 51.715 190.105 ;
        RECT 52.005 189.935 52.175 190.105 ;
        RECT 52.465 189.935 52.635 190.105 ;
        RECT 52.925 189.935 53.095 190.105 ;
        RECT 53.385 189.935 53.555 190.105 ;
        RECT 53.845 189.935 54.015 190.105 ;
        RECT 54.305 189.935 54.475 190.105 ;
        RECT 54.765 189.935 54.935 190.105 ;
        RECT 55.225 189.935 55.395 190.105 ;
        RECT 55.685 189.935 55.855 190.105 ;
        RECT 56.145 189.935 56.315 190.105 ;
        RECT 56.605 189.935 56.775 190.105 ;
        RECT 57.065 189.935 57.235 190.105 ;
        RECT 57.525 189.935 57.695 190.105 ;
        RECT 57.985 189.935 58.155 190.105 ;
        RECT 58.445 189.935 58.615 190.105 ;
        RECT 58.905 189.935 59.075 190.105 ;
        RECT 59.365 189.935 59.535 190.105 ;
        RECT 59.825 189.935 59.995 190.105 ;
        RECT 60.285 189.935 60.455 190.105 ;
        RECT 60.745 189.935 60.915 190.105 ;
        RECT 61.205 189.935 61.375 190.105 ;
        RECT 61.665 189.935 61.835 190.105 ;
        RECT 62.125 189.935 62.295 190.105 ;
        RECT 62.585 189.935 62.755 190.105 ;
        RECT 63.045 189.935 63.215 190.105 ;
        RECT 63.505 189.935 63.675 190.105 ;
        RECT 63.965 189.935 64.135 190.105 ;
        RECT 64.425 189.935 64.595 190.105 ;
        RECT 64.885 189.935 65.055 190.105 ;
        RECT 65.345 189.935 65.515 190.105 ;
        RECT 65.805 189.935 65.975 190.105 ;
        RECT 66.265 189.935 66.435 190.105 ;
        RECT 66.725 189.935 66.895 190.105 ;
        RECT 67.185 189.935 67.355 190.105 ;
        RECT 67.645 189.935 67.815 190.105 ;
        RECT 68.105 189.935 68.275 190.105 ;
        RECT 68.565 189.935 68.735 190.105 ;
        RECT 69.025 189.935 69.195 190.105 ;
        RECT 69.485 189.935 69.655 190.105 ;
        RECT 69.945 189.935 70.115 190.105 ;
        RECT 70.405 189.935 70.575 190.105 ;
        RECT 70.865 189.935 71.035 190.105 ;
        RECT 71.325 189.935 71.495 190.105 ;
        RECT 71.785 189.935 71.955 190.105 ;
        RECT 72.245 189.935 72.415 190.105 ;
        RECT 72.705 189.935 72.875 190.105 ;
        RECT 73.165 189.935 73.335 190.105 ;
        RECT 73.625 189.935 73.795 190.105 ;
        RECT 74.085 189.935 74.255 190.105 ;
        RECT 74.545 189.935 74.715 190.105 ;
        RECT 75.005 189.935 75.175 190.105 ;
        RECT 75.465 189.935 75.635 190.105 ;
        RECT 75.925 189.935 76.095 190.105 ;
        RECT 76.385 189.935 76.555 190.105 ;
        RECT 76.845 189.935 77.015 190.105 ;
        RECT 77.305 189.935 77.475 190.105 ;
        RECT 77.765 189.935 77.935 190.105 ;
        RECT 78.225 189.935 78.395 190.105 ;
        RECT 78.685 189.935 78.855 190.105 ;
        RECT 79.145 189.935 79.315 190.105 ;
        RECT 79.605 189.935 79.775 190.105 ;
        RECT 80.065 189.935 80.235 190.105 ;
        RECT 80.525 189.935 80.695 190.105 ;
        RECT 80.985 189.935 81.155 190.105 ;
        RECT 81.445 189.935 81.615 190.105 ;
        RECT 81.905 189.935 82.075 190.105 ;
        RECT 82.365 189.935 82.535 190.105 ;
        RECT 82.825 189.935 82.995 190.105 ;
        RECT 83.285 189.935 83.455 190.105 ;
        RECT 83.745 189.935 83.915 190.105 ;
        RECT 84.205 189.935 84.375 190.105 ;
        RECT 84.665 189.935 84.835 190.105 ;
        RECT 85.125 189.935 85.295 190.105 ;
        RECT 85.585 189.935 85.755 190.105 ;
        RECT 86.045 189.935 86.215 190.105 ;
        RECT 86.505 189.935 86.675 190.105 ;
        RECT 86.965 189.935 87.135 190.105 ;
        RECT 87.425 189.935 87.595 190.105 ;
        RECT 87.885 189.935 88.055 190.105 ;
        RECT 88.345 189.935 88.515 190.105 ;
        RECT 88.805 189.935 88.975 190.105 ;
        RECT 89.265 189.935 89.435 190.105 ;
        RECT 89.725 189.935 89.895 190.105 ;
        RECT 90.185 189.935 90.355 190.105 ;
        RECT 90.645 189.935 90.815 190.105 ;
        RECT 91.105 189.935 91.275 190.105 ;
        RECT 91.565 189.935 91.735 190.105 ;
        RECT 92.025 189.935 92.195 190.105 ;
        RECT 28.085 189.425 28.255 189.595 ;
        RECT 28.085 188.405 28.255 188.575 ;
        RECT 29.005 188.405 29.175 188.575 ;
        RECT 33.145 188.745 33.315 188.915 ;
        RECT 34.525 188.745 34.695 188.915 ;
        RECT 34.065 188.405 34.235 188.575 ;
        RECT 34.985 188.405 35.155 188.575 ;
        RECT 35.445 188.405 35.615 188.575 ;
        RECT 37.745 189.085 37.915 189.255 ;
        RECT 36.365 188.405 36.535 188.575 ;
        RECT 38.665 187.725 38.835 187.895 ;
        RECT 39.125 187.725 39.295 187.895 ;
        RECT 40.505 188.405 40.675 188.575 ;
        RECT 39.585 187.725 39.755 187.895 ;
        RECT 43.725 189.425 43.895 189.595 ;
        RECT 42.805 189.085 42.975 189.255 ;
        RECT 44.645 189.425 44.815 189.595 ;
        RECT 44.185 188.405 44.355 188.575 ;
        RECT 48.325 188.405 48.495 188.575 ;
        RECT 56.605 189.425 56.775 189.595 ;
        RECT 53.385 188.405 53.555 188.575 ;
        RECT 53.850 188.405 54.020 188.575 ;
        RECT 47.405 187.725 47.575 187.895 ;
        RECT 54.765 188.065 54.935 188.235 ;
        RECT 55.915 188.405 56.085 188.575 ;
        RECT 55.225 188.065 55.395 188.235 ;
        RECT 57.525 188.405 57.695 188.575 ;
        RECT 58.905 188.405 59.075 188.575 ;
        RECT 59.365 189.085 59.535 189.255 ;
        RECT 59.825 189.425 59.995 189.595 ;
        RECT 57.985 187.725 58.155 187.895 ;
        RECT 61.205 187.725 61.375 187.895 ;
        RECT 61.665 189.085 61.835 189.255 ;
        RECT 62.585 188.745 62.755 188.915 ;
        RECT 63.045 188.405 63.215 188.575 ;
        RECT 64.425 188.745 64.595 188.915 ;
        RECT 64.885 188.065 65.055 188.235 ;
        RECT 65.805 189.085 65.975 189.255 ;
        RECT 65.345 187.725 65.515 187.895 ;
        RECT 67.645 188.065 67.815 188.235 ;
        RECT 70.405 189.085 70.575 189.255 ;
        RECT 75.005 189.425 75.175 189.595 ;
        RECT 71.325 187.725 71.495 187.895 ;
        RECT 72.705 188.405 72.875 188.575 ;
        RECT 72.245 187.725 72.415 187.895 ;
        RECT 75.925 188.405 76.095 188.575 ;
        RECT 73.625 187.725 73.795 187.895 ;
        RECT 18.425 187.215 18.595 187.385 ;
        RECT 18.885 187.215 19.055 187.385 ;
        RECT 19.345 187.215 19.515 187.385 ;
        RECT 19.805 187.215 19.975 187.385 ;
        RECT 20.265 187.215 20.435 187.385 ;
        RECT 20.725 187.215 20.895 187.385 ;
        RECT 21.185 187.215 21.355 187.385 ;
        RECT 21.645 187.215 21.815 187.385 ;
        RECT 22.105 187.215 22.275 187.385 ;
        RECT 22.565 187.215 22.735 187.385 ;
        RECT 23.025 187.215 23.195 187.385 ;
        RECT 23.485 187.215 23.655 187.385 ;
        RECT 23.945 187.215 24.115 187.385 ;
        RECT 24.405 187.215 24.575 187.385 ;
        RECT 24.865 187.215 25.035 187.385 ;
        RECT 25.325 187.215 25.495 187.385 ;
        RECT 25.785 187.215 25.955 187.385 ;
        RECT 26.245 187.215 26.415 187.385 ;
        RECT 26.705 187.215 26.875 187.385 ;
        RECT 27.165 187.215 27.335 187.385 ;
        RECT 27.625 187.215 27.795 187.385 ;
        RECT 28.085 187.215 28.255 187.385 ;
        RECT 28.545 187.215 28.715 187.385 ;
        RECT 29.005 187.215 29.175 187.385 ;
        RECT 29.465 187.215 29.635 187.385 ;
        RECT 29.925 187.215 30.095 187.385 ;
        RECT 30.385 187.215 30.555 187.385 ;
        RECT 30.845 187.215 31.015 187.385 ;
        RECT 31.305 187.215 31.475 187.385 ;
        RECT 31.765 187.215 31.935 187.385 ;
        RECT 32.225 187.215 32.395 187.385 ;
        RECT 32.685 187.215 32.855 187.385 ;
        RECT 33.145 187.215 33.315 187.385 ;
        RECT 33.605 187.215 33.775 187.385 ;
        RECT 34.065 187.215 34.235 187.385 ;
        RECT 34.525 187.215 34.695 187.385 ;
        RECT 34.985 187.215 35.155 187.385 ;
        RECT 35.445 187.215 35.615 187.385 ;
        RECT 35.905 187.215 36.075 187.385 ;
        RECT 36.365 187.215 36.535 187.385 ;
        RECT 36.825 187.215 36.995 187.385 ;
        RECT 37.285 187.215 37.455 187.385 ;
        RECT 37.745 187.215 37.915 187.385 ;
        RECT 38.205 187.215 38.375 187.385 ;
        RECT 38.665 187.215 38.835 187.385 ;
        RECT 39.125 187.215 39.295 187.385 ;
        RECT 39.585 187.215 39.755 187.385 ;
        RECT 40.045 187.215 40.215 187.385 ;
        RECT 40.505 187.215 40.675 187.385 ;
        RECT 40.965 187.215 41.135 187.385 ;
        RECT 41.425 187.215 41.595 187.385 ;
        RECT 41.885 187.215 42.055 187.385 ;
        RECT 42.345 187.215 42.515 187.385 ;
        RECT 42.805 187.215 42.975 187.385 ;
        RECT 43.265 187.215 43.435 187.385 ;
        RECT 43.725 187.215 43.895 187.385 ;
        RECT 44.185 187.215 44.355 187.385 ;
        RECT 44.645 187.215 44.815 187.385 ;
        RECT 45.105 187.215 45.275 187.385 ;
        RECT 45.565 187.215 45.735 187.385 ;
        RECT 46.025 187.215 46.195 187.385 ;
        RECT 46.485 187.215 46.655 187.385 ;
        RECT 46.945 187.215 47.115 187.385 ;
        RECT 47.405 187.215 47.575 187.385 ;
        RECT 47.865 187.215 48.035 187.385 ;
        RECT 48.325 187.215 48.495 187.385 ;
        RECT 48.785 187.215 48.955 187.385 ;
        RECT 49.245 187.215 49.415 187.385 ;
        RECT 49.705 187.215 49.875 187.385 ;
        RECT 50.165 187.215 50.335 187.385 ;
        RECT 50.625 187.215 50.795 187.385 ;
        RECT 51.085 187.215 51.255 187.385 ;
        RECT 51.545 187.215 51.715 187.385 ;
        RECT 52.005 187.215 52.175 187.385 ;
        RECT 52.465 187.215 52.635 187.385 ;
        RECT 52.925 187.215 53.095 187.385 ;
        RECT 53.385 187.215 53.555 187.385 ;
        RECT 53.845 187.215 54.015 187.385 ;
        RECT 54.305 187.215 54.475 187.385 ;
        RECT 54.765 187.215 54.935 187.385 ;
        RECT 55.225 187.215 55.395 187.385 ;
        RECT 55.685 187.215 55.855 187.385 ;
        RECT 56.145 187.215 56.315 187.385 ;
        RECT 56.605 187.215 56.775 187.385 ;
        RECT 57.065 187.215 57.235 187.385 ;
        RECT 57.525 187.215 57.695 187.385 ;
        RECT 57.985 187.215 58.155 187.385 ;
        RECT 58.445 187.215 58.615 187.385 ;
        RECT 58.905 187.215 59.075 187.385 ;
        RECT 59.365 187.215 59.535 187.385 ;
        RECT 59.825 187.215 59.995 187.385 ;
        RECT 60.285 187.215 60.455 187.385 ;
        RECT 60.745 187.215 60.915 187.385 ;
        RECT 61.205 187.215 61.375 187.385 ;
        RECT 61.665 187.215 61.835 187.385 ;
        RECT 62.125 187.215 62.295 187.385 ;
        RECT 62.585 187.215 62.755 187.385 ;
        RECT 63.045 187.215 63.215 187.385 ;
        RECT 63.505 187.215 63.675 187.385 ;
        RECT 63.965 187.215 64.135 187.385 ;
        RECT 64.425 187.215 64.595 187.385 ;
        RECT 64.885 187.215 65.055 187.385 ;
        RECT 65.345 187.215 65.515 187.385 ;
        RECT 65.805 187.215 65.975 187.385 ;
        RECT 66.265 187.215 66.435 187.385 ;
        RECT 66.725 187.215 66.895 187.385 ;
        RECT 67.185 187.215 67.355 187.385 ;
        RECT 67.645 187.215 67.815 187.385 ;
        RECT 68.105 187.215 68.275 187.385 ;
        RECT 68.565 187.215 68.735 187.385 ;
        RECT 69.025 187.215 69.195 187.385 ;
        RECT 69.485 187.215 69.655 187.385 ;
        RECT 69.945 187.215 70.115 187.385 ;
        RECT 70.405 187.215 70.575 187.385 ;
        RECT 70.865 187.215 71.035 187.385 ;
        RECT 71.325 187.215 71.495 187.385 ;
        RECT 71.785 187.215 71.955 187.385 ;
        RECT 72.245 187.215 72.415 187.385 ;
        RECT 72.705 187.215 72.875 187.385 ;
        RECT 73.165 187.215 73.335 187.385 ;
        RECT 73.625 187.215 73.795 187.385 ;
        RECT 74.085 187.215 74.255 187.385 ;
        RECT 74.545 187.215 74.715 187.385 ;
        RECT 75.005 187.215 75.175 187.385 ;
        RECT 75.465 187.215 75.635 187.385 ;
        RECT 75.925 187.215 76.095 187.385 ;
        RECT 76.385 187.215 76.555 187.385 ;
        RECT 76.845 187.215 77.015 187.385 ;
        RECT 77.305 187.215 77.475 187.385 ;
        RECT 77.765 187.215 77.935 187.385 ;
        RECT 78.225 187.215 78.395 187.385 ;
        RECT 78.685 187.215 78.855 187.385 ;
        RECT 79.145 187.215 79.315 187.385 ;
        RECT 79.605 187.215 79.775 187.385 ;
        RECT 80.065 187.215 80.235 187.385 ;
        RECT 80.525 187.215 80.695 187.385 ;
        RECT 80.985 187.215 81.155 187.385 ;
        RECT 81.445 187.215 81.615 187.385 ;
        RECT 81.905 187.215 82.075 187.385 ;
        RECT 82.365 187.215 82.535 187.385 ;
        RECT 82.825 187.215 82.995 187.385 ;
        RECT 83.285 187.215 83.455 187.385 ;
        RECT 83.745 187.215 83.915 187.385 ;
        RECT 84.205 187.215 84.375 187.385 ;
        RECT 84.665 187.215 84.835 187.385 ;
        RECT 85.125 187.215 85.295 187.385 ;
        RECT 85.585 187.215 85.755 187.385 ;
        RECT 86.045 187.215 86.215 187.385 ;
        RECT 86.505 187.215 86.675 187.385 ;
        RECT 86.965 187.215 87.135 187.385 ;
        RECT 87.425 187.215 87.595 187.385 ;
        RECT 87.885 187.215 88.055 187.385 ;
        RECT 88.345 187.215 88.515 187.385 ;
        RECT 88.805 187.215 88.975 187.385 ;
        RECT 89.265 187.215 89.435 187.385 ;
        RECT 89.725 187.215 89.895 187.385 ;
        RECT 90.185 187.215 90.355 187.385 ;
        RECT 90.645 187.215 90.815 187.385 ;
        RECT 91.105 187.215 91.275 187.385 ;
        RECT 91.565 187.215 91.735 187.385 ;
        RECT 92.025 187.215 92.195 187.385 ;
        RECT 20.725 185.005 20.895 185.175 ;
        RECT 23.035 185.685 23.205 185.855 ;
        RECT 23.470 185.345 23.640 185.515 ;
        RECT 25.555 185.685 25.725 185.855 ;
        RECT 25.040 185.345 25.210 185.515 ;
        RECT 26.290 186.025 26.460 186.195 ;
        RECT 26.745 185.685 26.915 185.855 ;
        RECT 27.625 186.025 27.795 186.195 ;
        RECT 27.140 185.345 27.310 185.515 ;
        RECT 28.085 185.005 28.255 185.175 ;
        RECT 36.365 186.705 36.535 186.875 ;
        RECT 40.535 186.705 40.705 186.875 ;
        RECT 32.685 186.025 32.855 186.195 ;
        RECT 33.145 186.025 33.315 186.195 ;
        RECT 34.065 186.025 34.235 186.195 ;
        RECT 34.525 186.025 34.695 186.195 ;
        RECT 34.985 186.025 35.155 186.195 ;
        RECT 35.905 186.025 36.075 186.195 ;
        RECT 37.285 186.025 37.455 186.195 ;
        RECT 31.765 185.005 31.935 185.175 ;
        RECT 34.985 185.005 35.155 185.175 ;
        RECT 38.205 185.685 38.375 185.855 ;
        RECT 38.665 185.685 38.835 185.855 ;
        RECT 37.745 185.345 37.915 185.515 ;
        RECT 39.540 186.025 39.710 186.195 ;
        RECT 40.045 186.195 40.215 186.365 ;
        RECT 40.965 186.705 41.135 186.875 ;
        RECT 41.425 186.025 41.595 186.195 ;
        RECT 42.805 186.025 42.975 186.195 ;
        RECT 42.345 185.005 42.515 185.175 ;
        RECT 45.565 185.685 45.735 185.855 ;
        RECT 46.050 185.345 46.220 185.515 ;
        RECT 46.445 185.685 46.615 185.855 ;
        RECT 46.900 186.365 47.070 186.535 ;
        RECT 47.635 185.685 47.805 185.855 ;
        RECT 48.150 185.345 48.320 185.515 ;
        RECT 49.720 185.345 49.890 185.515 ;
        RECT 50.155 185.685 50.325 185.855 ;
        RECT 52.465 185.005 52.635 185.175 ;
        RECT 60.285 186.025 60.455 186.195 ;
        RECT 61.665 186.025 61.835 186.195 ;
        RECT 62.125 186.025 62.295 186.195 ;
        RECT 60.745 185.685 60.915 185.855 ;
        RECT 63.045 185.345 63.215 185.515 ;
        RECT 64.425 186.025 64.595 186.195 ;
        RECT 63.505 185.005 63.675 185.175 ;
        RECT 64.885 185.345 65.055 185.515 ;
        RECT 65.345 186.025 65.515 186.195 ;
        RECT 65.805 186.025 65.975 186.195 ;
        RECT 67.185 186.025 67.355 186.195 ;
        RECT 70.405 186.705 70.575 186.875 ;
        RECT 69.485 185.685 69.655 185.855 ;
        RECT 68.565 185.005 68.735 185.175 ;
        RECT 71.325 186.025 71.495 186.195 ;
        RECT 73.165 186.025 73.335 186.195 ;
        RECT 71.325 185.005 71.495 185.175 ;
        RECT 75.465 186.025 75.635 186.195 ;
        RECT 75.005 185.685 75.175 185.855 ;
        RECT 77.765 186.365 77.935 186.535 ;
        RECT 77.305 186.025 77.475 186.195 ;
        RECT 78.225 186.025 78.395 186.195 ;
        RECT 78.685 186.025 78.855 186.195 ;
        RECT 80.065 186.025 80.235 186.195 ;
        RECT 80.525 186.025 80.695 186.195 ;
        RECT 73.625 185.005 73.795 185.175 ;
        RECT 82.365 186.025 82.535 186.195 ;
        RECT 81.905 185.005 82.075 185.175 ;
        RECT 82.830 185.345 83.000 185.515 ;
        RECT 83.290 186.365 83.460 186.535 ;
        RECT 83.745 185.685 83.915 185.855 ;
        RECT 84.690 186.365 84.860 186.535 ;
        RECT 86.530 186.365 86.700 186.535 ;
        RECT 85.150 185.345 85.320 185.515 ;
        RECT 86.530 185.345 86.700 185.515 ;
        RECT 90.185 185.005 90.355 185.175 ;
        RECT 18.425 184.495 18.595 184.665 ;
        RECT 18.885 184.495 19.055 184.665 ;
        RECT 19.345 184.495 19.515 184.665 ;
        RECT 19.805 184.495 19.975 184.665 ;
        RECT 20.265 184.495 20.435 184.665 ;
        RECT 20.725 184.495 20.895 184.665 ;
        RECT 21.185 184.495 21.355 184.665 ;
        RECT 21.645 184.495 21.815 184.665 ;
        RECT 22.105 184.495 22.275 184.665 ;
        RECT 22.565 184.495 22.735 184.665 ;
        RECT 23.025 184.495 23.195 184.665 ;
        RECT 23.485 184.495 23.655 184.665 ;
        RECT 23.945 184.495 24.115 184.665 ;
        RECT 24.405 184.495 24.575 184.665 ;
        RECT 24.865 184.495 25.035 184.665 ;
        RECT 25.325 184.495 25.495 184.665 ;
        RECT 25.785 184.495 25.955 184.665 ;
        RECT 26.245 184.495 26.415 184.665 ;
        RECT 26.705 184.495 26.875 184.665 ;
        RECT 27.165 184.495 27.335 184.665 ;
        RECT 27.625 184.495 27.795 184.665 ;
        RECT 28.085 184.495 28.255 184.665 ;
        RECT 28.545 184.495 28.715 184.665 ;
        RECT 29.005 184.495 29.175 184.665 ;
        RECT 29.465 184.495 29.635 184.665 ;
        RECT 29.925 184.495 30.095 184.665 ;
        RECT 30.385 184.495 30.555 184.665 ;
        RECT 30.845 184.495 31.015 184.665 ;
        RECT 31.305 184.495 31.475 184.665 ;
        RECT 31.765 184.495 31.935 184.665 ;
        RECT 32.225 184.495 32.395 184.665 ;
        RECT 32.685 184.495 32.855 184.665 ;
        RECT 33.145 184.495 33.315 184.665 ;
        RECT 33.605 184.495 33.775 184.665 ;
        RECT 34.065 184.495 34.235 184.665 ;
        RECT 34.525 184.495 34.695 184.665 ;
        RECT 34.985 184.495 35.155 184.665 ;
        RECT 35.445 184.495 35.615 184.665 ;
        RECT 35.905 184.495 36.075 184.665 ;
        RECT 36.365 184.495 36.535 184.665 ;
        RECT 36.825 184.495 36.995 184.665 ;
        RECT 37.285 184.495 37.455 184.665 ;
        RECT 37.745 184.495 37.915 184.665 ;
        RECT 38.205 184.495 38.375 184.665 ;
        RECT 38.665 184.495 38.835 184.665 ;
        RECT 39.125 184.495 39.295 184.665 ;
        RECT 39.585 184.495 39.755 184.665 ;
        RECT 40.045 184.495 40.215 184.665 ;
        RECT 40.505 184.495 40.675 184.665 ;
        RECT 40.965 184.495 41.135 184.665 ;
        RECT 41.425 184.495 41.595 184.665 ;
        RECT 41.885 184.495 42.055 184.665 ;
        RECT 42.345 184.495 42.515 184.665 ;
        RECT 42.805 184.495 42.975 184.665 ;
        RECT 43.265 184.495 43.435 184.665 ;
        RECT 43.725 184.495 43.895 184.665 ;
        RECT 44.185 184.495 44.355 184.665 ;
        RECT 44.645 184.495 44.815 184.665 ;
        RECT 45.105 184.495 45.275 184.665 ;
        RECT 45.565 184.495 45.735 184.665 ;
        RECT 46.025 184.495 46.195 184.665 ;
        RECT 46.485 184.495 46.655 184.665 ;
        RECT 46.945 184.495 47.115 184.665 ;
        RECT 47.405 184.495 47.575 184.665 ;
        RECT 47.865 184.495 48.035 184.665 ;
        RECT 48.325 184.495 48.495 184.665 ;
        RECT 48.785 184.495 48.955 184.665 ;
        RECT 49.245 184.495 49.415 184.665 ;
        RECT 49.705 184.495 49.875 184.665 ;
        RECT 50.165 184.495 50.335 184.665 ;
        RECT 50.625 184.495 50.795 184.665 ;
        RECT 51.085 184.495 51.255 184.665 ;
        RECT 51.545 184.495 51.715 184.665 ;
        RECT 52.005 184.495 52.175 184.665 ;
        RECT 52.465 184.495 52.635 184.665 ;
        RECT 52.925 184.495 53.095 184.665 ;
        RECT 53.385 184.495 53.555 184.665 ;
        RECT 53.845 184.495 54.015 184.665 ;
        RECT 54.305 184.495 54.475 184.665 ;
        RECT 54.765 184.495 54.935 184.665 ;
        RECT 55.225 184.495 55.395 184.665 ;
        RECT 55.685 184.495 55.855 184.665 ;
        RECT 56.145 184.495 56.315 184.665 ;
        RECT 56.605 184.495 56.775 184.665 ;
        RECT 57.065 184.495 57.235 184.665 ;
        RECT 57.525 184.495 57.695 184.665 ;
        RECT 57.985 184.495 58.155 184.665 ;
        RECT 58.445 184.495 58.615 184.665 ;
        RECT 58.905 184.495 59.075 184.665 ;
        RECT 59.365 184.495 59.535 184.665 ;
        RECT 59.825 184.495 59.995 184.665 ;
        RECT 60.285 184.495 60.455 184.665 ;
        RECT 60.745 184.495 60.915 184.665 ;
        RECT 61.205 184.495 61.375 184.665 ;
        RECT 61.665 184.495 61.835 184.665 ;
        RECT 62.125 184.495 62.295 184.665 ;
        RECT 62.585 184.495 62.755 184.665 ;
        RECT 63.045 184.495 63.215 184.665 ;
        RECT 63.505 184.495 63.675 184.665 ;
        RECT 63.965 184.495 64.135 184.665 ;
        RECT 64.425 184.495 64.595 184.665 ;
        RECT 64.885 184.495 65.055 184.665 ;
        RECT 65.345 184.495 65.515 184.665 ;
        RECT 65.805 184.495 65.975 184.665 ;
        RECT 66.265 184.495 66.435 184.665 ;
        RECT 66.725 184.495 66.895 184.665 ;
        RECT 67.185 184.495 67.355 184.665 ;
        RECT 67.645 184.495 67.815 184.665 ;
        RECT 68.105 184.495 68.275 184.665 ;
        RECT 68.565 184.495 68.735 184.665 ;
        RECT 69.025 184.495 69.195 184.665 ;
        RECT 69.485 184.495 69.655 184.665 ;
        RECT 69.945 184.495 70.115 184.665 ;
        RECT 70.405 184.495 70.575 184.665 ;
        RECT 70.865 184.495 71.035 184.665 ;
        RECT 71.325 184.495 71.495 184.665 ;
        RECT 71.785 184.495 71.955 184.665 ;
        RECT 72.245 184.495 72.415 184.665 ;
        RECT 72.705 184.495 72.875 184.665 ;
        RECT 73.165 184.495 73.335 184.665 ;
        RECT 73.625 184.495 73.795 184.665 ;
        RECT 74.085 184.495 74.255 184.665 ;
        RECT 74.545 184.495 74.715 184.665 ;
        RECT 75.005 184.495 75.175 184.665 ;
        RECT 75.465 184.495 75.635 184.665 ;
        RECT 75.925 184.495 76.095 184.665 ;
        RECT 76.385 184.495 76.555 184.665 ;
        RECT 76.845 184.495 77.015 184.665 ;
        RECT 77.305 184.495 77.475 184.665 ;
        RECT 77.765 184.495 77.935 184.665 ;
        RECT 78.225 184.495 78.395 184.665 ;
        RECT 78.685 184.495 78.855 184.665 ;
        RECT 79.145 184.495 79.315 184.665 ;
        RECT 79.605 184.495 79.775 184.665 ;
        RECT 80.065 184.495 80.235 184.665 ;
        RECT 80.525 184.495 80.695 184.665 ;
        RECT 80.985 184.495 81.155 184.665 ;
        RECT 81.445 184.495 81.615 184.665 ;
        RECT 81.905 184.495 82.075 184.665 ;
        RECT 82.365 184.495 82.535 184.665 ;
        RECT 82.825 184.495 82.995 184.665 ;
        RECT 83.285 184.495 83.455 184.665 ;
        RECT 83.745 184.495 83.915 184.665 ;
        RECT 84.205 184.495 84.375 184.665 ;
        RECT 84.665 184.495 84.835 184.665 ;
        RECT 85.125 184.495 85.295 184.665 ;
        RECT 85.585 184.495 85.755 184.665 ;
        RECT 86.045 184.495 86.215 184.665 ;
        RECT 86.505 184.495 86.675 184.665 ;
        RECT 86.965 184.495 87.135 184.665 ;
        RECT 87.425 184.495 87.595 184.665 ;
        RECT 87.885 184.495 88.055 184.665 ;
        RECT 88.345 184.495 88.515 184.665 ;
        RECT 88.805 184.495 88.975 184.665 ;
        RECT 89.265 184.495 89.435 184.665 ;
        RECT 89.725 184.495 89.895 184.665 ;
        RECT 90.185 184.495 90.355 184.665 ;
        RECT 90.645 184.495 90.815 184.665 ;
        RECT 91.105 184.495 91.275 184.665 ;
        RECT 91.565 184.495 91.735 184.665 ;
        RECT 92.025 184.495 92.195 184.665 ;
        RECT 27.165 183.985 27.335 184.155 ;
        RECT 27.165 182.625 27.335 182.795 ;
        RECT 28.545 182.965 28.715 183.135 ;
        RECT 29.005 182.965 29.175 183.135 ;
        RECT 34.065 183.985 34.235 184.155 ;
        RECT 29.925 182.965 30.095 183.135 ;
        RECT 40.965 183.985 41.135 184.155 ;
        RECT 28.085 182.285 28.255 182.455 ;
        RECT 29.465 182.285 29.635 182.455 ;
        RECT 40.505 182.965 40.675 183.135 ;
        RECT 41.885 182.965 42.055 183.135 ;
        RECT 42.345 182.965 42.515 183.135 ;
        RECT 44.185 182.625 44.355 182.795 ;
        RECT 47.405 183.985 47.575 184.155 ;
        RECT 46.025 182.965 46.195 183.135 ;
        RECT 46.485 182.965 46.655 183.135 ;
        RECT 45.105 182.625 45.275 182.795 ;
        RECT 47.865 182.965 48.035 183.135 ;
        RECT 48.785 182.965 48.955 183.135 ;
        RECT 50.295 182.965 50.465 183.135 ;
        RECT 51.085 182.965 51.255 183.135 ;
        RECT 56.145 183.985 56.315 184.155 ;
        RECT 64.885 183.985 65.055 184.155 ;
        RECT 56.605 182.965 56.775 183.135 ;
        RECT 57.525 182.965 57.695 183.135 ;
        RECT 68.105 183.645 68.275 183.815 ;
        RECT 73.625 183.645 73.795 183.815 ;
        RECT 69.485 182.965 69.655 183.135 ;
        RECT 69.945 182.965 70.115 183.135 ;
        RECT 70.405 182.965 70.575 183.135 ;
        RECT 71.325 182.965 71.495 183.135 ;
        RECT 72.245 182.625 72.415 182.795 ;
        RECT 80.065 183.985 80.235 184.155 ;
        RECT 83.285 183.985 83.455 184.155 ;
        RECT 86.965 183.985 87.135 184.155 ;
        RECT 87.885 183.985 88.055 184.155 ;
        RECT 80.985 182.965 81.155 183.135 ;
        RECT 81.905 182.965 82.075 183.135 ;
        RECT 82.365 182.965 82.535 183.135 ;
        RECT 84.665 182.965 84.835 183.135 ;
        RECT 85.125 182.965 85.295 183.135 ;
        RECT 85.585 182.965 85.755 183.135 ;
        RECT 86.505 182.965 86.675 183.135 ;
        RECT 87.755 182.285 87.925 182.455 ;
        RECT 88.805 182.625 88.975 182.795 ;
        RECT 18.425 181.775 18.595 181.945 ;
        RECT 18.885 181.775 19.055 181.945 ;
        RECT 19.345 181.775 19.515 181.945 ;
        RECT 19.805 181.775 19.975 181.945 ;
        RECT 20.265 181.775 20.435 181.945 ;
        RECT 20.725 181.775 20.895 181.945 ;
        RECT 21.185 181.775 21.355 181.945 ;
        RECT 21.645 181.775 21.815 181.945 ;
        RECT 22.105 181.775 22.275 181.945 ;
        RECT 22.565 181.775 22.735 181.945 ;
        RECT 23.025 181.775 23.195 181.945 ;
        RECT 23.485 181.775 23.655 181.945 ;
        RECT 23.945 181.775 24.115 181.945 ;
        RECT 24.405 181.775 24.575 181.945 ;
        RECT 24.865 181.775 25.035 181.945 ;
        RECT 25.325 181.775 25.495 181.945 ;
        RECT 25.785 181.775 25.955 181.945 ;
        RECT 26.245 181.775 26.415 181.945 ;
        RECT 26.705 181.775 26.875 181.945 ;
        RECT 27.165 181.775 27.335 181.945 ;
        RECT 27.625 181.775 27.795 181.945 ;
        RECT 28.085 181.775 28.255 181.945 ;
        RECT 28.545 181.775 28.715 181.945 ;
        RECT 29.005 181.775 29.175 181.945 ;
        RECT 29.465 181.775 29.635 181.945 ;
        RECT 29.925 181.775 30.095 181.945 ;
        RECT 30.385 181.775 30.555 181.945 ;
        RECT 30.845 181.775 31.015 181.945 ;
        RECT 31.305 181.775 31.475 181.945 ;
        RECT 31.765 181.775 31.935 181.945 ;
        RECT 32.225 181.775 32.395 181.945 ;
        RECT 32.685 181.775 32.855 181.945 ;
        RECT 33.145 181.775 33.315 181.945 ;
        RECT 33.605 181.775 33.775 181.945 ;
        RECT 34.065 181.775 34.235 181.945 ;
        RECT 34.525 181.775 34.695 181.945 ;
        RECT 34.985 181.775 35.155 181.945 ;
        RECT 35.445 181.775 35.615 181.945 ;
        RECT 35.905 181.775 36.075 181.945 ;
        RECT 36.365 181.775 36.535 181.945 ;
        RECT 36.825 181.775 36.995 181.945 ;
        RECT 37.285 181.775 37.455 181.945 ;
        RECT 37.745 181.775 37.915 181.945 ;
        RECT 38.205 181.775 38.375 181.945 ;
        RECT 38.665 181.775 38.835 181.945 ;
        RECT 39.125 181.775 39.295 181.945 ;
        RECT 39.585 181.775 39.755 181.945 ;
        RECT 40.045 181.775 40.215 181.945 ;
        RECT 40.505 181.775 40.675 181.945 ;
        RECT 40.965 181.775 41.135 181.945 ;
        RECT 41.425 181.775 41.595 181.945 ;
        RECT 41.885 181.775 42.055 181.945 ;
        RECT 42.345 181.775 42.515 181.945 ;
        RECT 42.805 181.775 42.975 181.945 ;
        RECT 43.265 181.775 43.435 181.945 ;
        RECT 43.725 181.775 43.895 181.945 ;
        RECT 44.185 181.775 44.355 181.945 ;
        RECT 44.645 181.775 44.815 181.945 ;
        RECT 45.105 181.775 45.275 181.945 ;
        RECT 45.565 181.775 45.735 181.945 ;
        RECT 46.025 181.775 46.195 181.945 ;
        RECT 46.485 181.775 46.655 181.945 ;
        RECT 46.945 181.775 47.115 181.945 ;
        RECT 47.405 181.775 47.575 181.945 ;
        RECT 47.865 181.775 48.035 181.945 ;
        RECT 48.325 181.775 48.495 181.945 ;
        RECT 48.785 181.775 48.955 181.945 ;
        RECT 49.245 181.775 49.415 181.945 ;
        RECT 49.705 181.775 49.875 181.945 ;
        RECT 50.165 181.775 50.335 181.945 ;
        RECT 50.625 181.775 50.795 181.945 ;
        RECT 51.085 181.775 51.255 181.945 ;
        RECT 51.545 181.775 51.715 181.945 ;
        RECT 52.005 181.775 52.175 181.945 ;
        RECT 52.465 181.775 52.635 181.945 ;
        RECT 52.925 181.775 53.095 181.945 ;
        RECT 53.385 181.775 53.555 181.945 ;
        RECT 53.845 181.775 54.015 181.945 ;
        RECT 54.305 181.775 54.475 181.945 ;
        RECT 54.765 181.775 54.935 181.945 ;
        RECT 55.225 181.775 55.395 181.945 ;
        RECT 55.685 181.775 55.855 181.945 ;
        RECT 56.145 181.775 56.315 181.945 ;
        RECT 56.605 181.775 56.775 181.945 ;
        RECT 57.065 181.775 57.235 181.945 ;
        RECT 57.525 181.775 57.695 181.945 ;
        RECT 57.985 181.775 58.155 181.945 ;
        RECT 58.445 181.775 58.615 181.945 ;
        RECT 58.905 181.775 59.075 181.945 ;
        RECT 59.365 181.775 59.535 181.945 ;
        RECT 59.825 181.775 59.995 181.945 ;
        RECT 60.285 181.775 60.455 181.945 ;
        RECT 60.745 181.775 60.915 181.945 ;
        RECT 61.205 181.775 61.375 181.945 ;
        RECT 61.665 181.775 61.835 181.945 ;
        RECT 62.125 181.775 62.295 181.945 ;
        RECT 62.585 181.775 62.755 181.945 ;
        RECT 63.045 181.775 63.215 181.945 ;
        RECT 63.505 181.775 63.675 181.945 ;
        RECT 63.965 181.775 64.135 181.945 ;
        RECT 64.425 181.775 64.595 181.945 ;
        RECT 64.885 181.775 65.055 181.945 ;
        RECT 65.345 181.775 65.515 181.945 ;
        RECT 65.805 181.775 65.975 181.945 ;
        RECT 66.265 181.775 66.435 181.945 ;
        RECT 66.725 181.775 66.895 181.945 ;
        RECT 67.185 181.775 67.355 181.945 ;
        RECT 67.645 181.775 67.815 181.945 ;
        RECT 68.105 181.775 68.275 181.945 ;
        RECT 68.565 181.775 68.735 181.945 ;
        RECT 69.025 181.775 69.195 181.945 ;
        RECT 69.485 181.775 69.655 181.945 ;
        RECT 69.945 181.775 70.115 181.945 ;
        RECT 70.405 181.775 70.575 181.945 ;
        RECT 70.865 181.775 71.035 181.945 ;
        RECT 71.325 181.775 71.495 181.945 ;
        RECT 71.785 181.775 71.955 181.945 ;
        RECT 72.245 181.775 72.415 181.945 ;
        RECT 72.705 181.775 72.875 181.945 ;
        RECT 73.165 181.775 73.335 181.945 ;
        RECT 73.625 181.775 73.795 181.945 ;
        RECT 74.085 181.775 74.255 181.945 ;
        RECT 74.545 181.775 74.715 181.945 ;
        RECT 75.005 181.775 75.175 181.945 ;
        RECT 75.465 181.775 75.635 181.945 ;
        RECT 75.925 181.775 76.095 181.945 ;
        RECT 76.385 181.775 76.555 181.945 ;
        RECT 76.845 181.775 77.015 181.945 ;
        RECT 77.305 181.775 77.475 181.945 ;
        RECT 77.765 181.775 77.935 181.945 ;
        RECT 78.225 181.775 78.395 181.945 ;
        RECT 78.685 181.775 78.855 181.945 ;
        RECT 79.145 181.775 79.315 181.945 ;
        RECT 79.605 181.775 79.775 181.945 ;
        RECT 80.065 181.775 80.235 181.945 ;
        RECT 80.525 181.775 80.695 181.945 ;
        RECT 80.985 181.775 81.155 181.945 ;
        RECT 81.445 181.775 81.615 181.945 ;
        RECT 81.905 181.775 82.075 181.945 ;
        RECT 82.365 181.775 82.535 181.945 ;
        RECT 82.825 181.775 82.995 181.945 ;
        RECT 83.285 181.775 83.455 181.945 ;
        RECT 83.745 181.775 83.915 181.945 ;
        RECT 84.205 181.775 84.375 181.945 ;
        RECT 84.665 181.775 84.835 181.945 ;
        RECT 85.125 181.775 85.295 181.945 ;
        RECT 85.585 181.775 85.755 181.945 ;
        RECT 86.045 181.775 86.215 181.945 ;
        RECT 86.505 181.775 86.675 181.945 ;
        RECT 86.965 181.775 87.135 181.945 ;
        RECT 87.425 181.775 87.595 181.945 ;
        RECT 87.885 181.775 88.055 181.945 ;
        RECT 88.345 181.775 88.515 181.945 ;
        RECT 88.805 181.775 88.975 181.945 ;
        RECT 89.265 181.775 89.435 181.945 ;
        RECT 89.725 181.775 89.895 181.945 ;
        RECT 90.185 181.775 90.355 181.945 ;
        RECT 90.645 181.775 90.815 181.945 ;
        RECT 91.105 181.775 91.275 181.945 ;
        RECT 91.565 181.775 91.735 181.945 ;
        RECT 92.025 181.775 92.195 181.945 ;
        RECT 37.285 181.265 37.455 181.435 ;
        RECT 38.125 180.925 38.295 181.095 ;
        RECT 39.125 180.925 39.295 181.095 ;
        RECT 42.345 181.265 42.515 181.435 ;
        RECT 41.885 180.585 42.055 180.755 ;
        RECT 42.805 180.585 42.975 180.755 ;
        RECT 38.205 179.565 38.375 179.735 ;
        RECT 59.365 180.585 59.535 180.755 ;
        RECT 60.285 180.585 60.455 180.755 ;
        RECT 60.745 180.585 60.915 180.755 ;
        RECT 61.665 180.585 61.835 180.755 ;
        RECT 58.445 179.905 58.615 180.075 ;
        RECT 62.585 180.585 62.755 180.755 ;
        RECT 61.205 179.565 61.375 179.735 ;
        RECT 63.965 179.565 64.135 179.735 ;
        RECT 71.785 180.585 71.955 180.755 ;
        RECT 72.245 180.245 72.415 180.415 ;
        RECT 72.705 180.245 72.875 180.415 ;
        RECT 73.165 180.245 73.335 180.415 ;
        RECT 74.085 179.565 74.255 179.735 ;
        RECT 18.425 179.055 18.595 179.225 ;
        RECT 18.885 179.055 19.055 179.225 ;
        RECT 19.345 179.055 19.515 179.225 ;
        RECT 19.805 179.055 19.975 179.225 ;
        RECT 20.265 179.055 20.435 179.225 ;
        RECT 20.725 179.055 20.895 179.225 ;
        RECT 21.185 179.055 21.355 179.225 ;
        RECT 21.645 179.055 21.815 179.225 ;
        RECT 22.105 179.055 22.275 179.225 ;
        RECT 22.565 179.055 22.735 179.225 ;
        RECT 23.025 179.055 23.195 179.225 ;
        RECT 23.485 179.055 23.655 179.225 ;
        RECT 23.945 179.055 24.115 179.225 ;
        RECT 24.405 179.055 24.575 179.225 ;
        RECT 24.865 179.055 25.035 179.225 ;
        RECT 25.325 179.055 25.495 179.225 ;
        RECT 25.785 179.055 25.955 179.225 ;
        RECT 26.245 179.055 26.415 179.225 ;
        RECT 26.705 179.055 26.875 179.225 ;
        RECT 27.165 179.055 27.335 179.225 ;
        RECT 27.625 179.055 27.795 179.225 ;
        RECT 28.085 179.055 28.255 179.225 ;
        RECT 28.545 179.055 28.715 179.225 ;
        RECT 29.005 179.055 29.175 179.225 ;
        RECT 29.465 179.055 29.635 179.225 ;
        RECT 29.925 179.055 30.095 179.225 ;
        RECT 30.385 179.055 30.555 179.225 ;
        RECT 30.845 179.055 31.015 179.225 ;
        RECT 31.305 179.055 31.475 179.225 ;
        RECT 31.765 179.055 31.935 179.225 ;
        RECT 32.225 179.055 32.395 179.225 ;
        RECT 32.685 179.055 32.855 179.225 ;
        RECT 33.145 179.055 33.315 179.225 ;
        RECT 33.605 179.055 33.775 179.225 ;
        RECT 34.065 179.055 34.235 179.225 ;
        RECT 34.525 179.055 34.695 179.225 ;
        RECT 34.985 179.055 35.155 179.225 ;
        RECT 35.445 179.055 35.615 179.225 ;
        RECT 35.905 179.055 36.075 179.225 ;
        RECT 36.365 179.055 36.535 179.225 ;
        RECT 36.825 179.055 36.995 179.225 ;
        RECT 37.285 179.055 37.455 179.225 ;
        RECT 37.745 179.055 37.915 179.225 ;
        RECT 38.205 179.055 38.375 179.225 ;
        RECT 38.665 179.055 38.835 179.225 ;
        RECT 39.125 179.055 39.295 179.225 ;
        RECT 39.585 179.055 39.755 179.225 ;
        RECT 40.045 179.055 40.215 179.225 ;
        RECT 40.505 179.055 40.675 179.225 ;
        RECT 40.965 179.055 41.135 179.225 ;
        RECT 41.425 179.055 41.595 179.225 ;
        RECT 41.885 179.055 42.055 179.225 ;
        RECT 42.345 179.055 42.515 179.225 ;
        RECT 42.805 179.055 42.975 179.225 ;
        RECT 43.265 179.055 43.435 179.225 ;
        RECT 43.725 179.055 43.895 179.225 ;
        RECT 44.185 179.055 44.355 179.225 ;
        RECT 44.645 179.055 44.815 179.225 ;
        RECT 45.105 179.055 45.275 179.225 ;
        RECT 45.565 179.055 45.735 179.225 ;
        RECT 46.025 179.055 46.195 179.225 ;
        RECT 46.485 179.055 46.655 179.225 ;
        RECT 46.945 179.055 47.115 179.225 ;
        RECT 47.405 179.055 47.575 179.225 ;
        RECT 47.865 179.055 48.035 179.225 ;
        RECT 48.325 179.055 48.495 179.225 ;
        RECT 48.785 179.055 48.955 179.225 ;
        RECT 49.245 179.055 49.415 179.225 ;
        RECT 49.705 179.055 49.875 179.225 ;
        RECT 50.165 179.055 50.335 179.225 ;
        RECT 50.625 179.055 50.795 179.225 ;
        RECT 51.085 179.055 51.255 179.225 ;
        RECT 51.545 179.055 51.715 179.225 ;
        RECT 52.005 179.055 52.175 179.225 ;
        RECT 52.465 179.055 52.635 179.225 ;
        RECT 52.925 179.055 53.095 179.225 ;
        RECT 53.385 179.055 53.555 179.225 ;
        RECT 53.845 179.055 54.015 179.225 ;
        RECT 54.305 179.055 54.475 179.225 ;
        RECT 54.765 179.055 54.935 179.225 ;
        RECT 55.225 179.055 55.395 179.225 ;
        RECT 55.685 179.055 55.855 179.225 ;
        RECT 56.145 179.055 56.315 179.225 ;
        RECT 56.605 179.055 56.775 179.225 ;
        RECT 57.065 179.055 57.235 179.225 ;
        RECT 57.525 179.055 57.695 179.225 ;
        RECT 57.985 179.055 58.155 179.225 ;
        RECT 58.445 179.055 58.615 179.225 ;
        RECT 58.905 179.055 59.075 179.225 ;
        RECT 59.365 179.055 59.535 179.225 ;
        RECT 59.825 179.055 59.995 179.225 ;
        RECT 60.285 179.055 60.455 179.225 ;
        RECT 60.745 179.055 60.915 179.225 ;
        RECT 61.205 179.055 61.375 179.225 ;
        RECT 61.665 179.055 61.835 179.225 ;
        RECT 62.125 179.055 62.295 179.225 ;
        RECT 62.585 179.055 62.755 179.225 ;
        RECT 63.045 179.055 63.215 179.225 ;
        RECT 63.505 179.055 63.675 179.225 ;
        RECT 63.965 179.055 64.135 179.225 ;
        RECT 64.425 179.055 64.595 179.225 ;
        RECT 64.885 179.055 65.055 179.225 ;
        RECT 65.345 179.055 65.515 179.225 ;
        RECT 65.805 179.055 65.975 179.225 ;
        RECT 66.265 179.055 66.435 179.225 ;
        RECT 66.725 179.055 66.895 179.225 ;
        RECT 67.185 179.055 67.355 179.225 ;
        RECT 67.645 179.055 67.815 179.225 ;
        RECT 68.105 179.055 68.275 179.225 ;
        RECT 68.565 179.055 68.735 179.225 ;
        RECT 69.025 179.055 69.195 179.225 ;
        RECT 69.485 179.055 69.655 179.225 ;
        RECT 69.945 179.055 70.115 179.225 ;
        RECT 70.405 179.055 70.575 179.225 ;
        RECT 70.865 179.055 71.035 179.225 ;
        RECT 71.325 179.055 71.495 179.225 ;
        RECT 71.785 179.055 71.955 179.225 ;
        RECT 72.245 179.055 72.415 179.225 ;
        RECT 72.705 179.055 72.875 179.225 ;
        RECT 73.165 179.055 73.335 179.225 ;
        RECT 73.625 179.055 73.795 179.225 ;
        RECT 74.085 179.055 74.255 179.225 ;
        RECT 74.545 179.055 74.715 179.225 ;
        RECT 75.005 179.055 75.175 179.225 ;
        RECT 75.465 179.055 75.635 179.225 ;
        RECT 75.925 179.055 76.095 179.225 ;
        RECT 76.385 179.055 76.555 179.225 ;
        RECT 76.845 179.055 77.015 179.225 ;
        RECT 77.305 179.055 77.475 179.225 ;
        RECT 77.765 179.055 77.935 179.225 ;
        RECT 78.225 179.055 78.395 179.225 ;
        RECT 78.685 179.055 78.855 179.225 ;
        RECT 79.145 179.055 79.315 179.225 ;
        RECT 79.605 179.055 79.775 179.225 ;
        RECT 80.065 179.055 80.235 179.225 ;
        RECT 80.525 179.055 80.695 179.225 ;
        RECT 80.985 179.055 81.155 179.225 ;
        RECT 81.445 179.055 81.615 179.225 ;
        RECT 81.905 179.055 82.075 179.225 ;
        RECT 82.365 179.055 82.535 179.225 ;
        RECT 82.825 179.055 82.995 179.225 ;
        RECT 83.285 179.055 83.455 179.225 ;
        RECT 83.745 179.055 83.915 179.225 ;
        RECT 84.205 179.055 84.375 179.225 ;
        RECT 84.665 179.055 84.835 179.225 ;
        RECT 85.125 179.055 85.295 179.225 ;
        RECT 85.585 179.055 85.755 179.225 ;
        RECT 86.045 179.055 86.215 179.225 ;
        RECT 86.505 179.055 86.675 179.225 ;
        RECT 86.965 179.055 87.135 179.225 ;
        RECT 87.425 179.055 87.595 179.225 ;
        RECT 87.885 179.055 88.055 179.225 ;
        RECT 88.345 179.055 88.515 179.225 ;
        RECT 88.805 179.055 88.975 179.225 ;
        RECT 89.265 179.055 89.435 179.225 ;
        RECT 89.725 179.055 89.895 179.225 ;
        RECT 90.185 179.055 90.355 179.225 ;
        RECT 90.645 179.055 90.815 179.225 ;
        RECT 91.105 179.055 91.275 179.225 ;
        RECT 91.565 179.055 91.735 179.225 ;
        RECT 92.025 179.055 92.195 179.225 ;
        RECT 24.430 178.205 24.600 178.375 ;
        RECT 23.945 177.525 24.115 177.695 ;
        RECT 24.825 177.865 24.995 178.035 ;
        RECT 25.280 177.185 25.450 177.355 ;
        RECT 26.530 178.205 26.700 178.375 ;
        RECT 26.015 177.865 26.185 178.035 ;
        RECT 28.100 178.205 28.270 178.375 ;
        RECT 28.535 177.865 28.705 178.035 ;
        RECT 30.845 178.205 31.015 178.375 ;
        RECT 33.145 178.205 33.315 178.375 ;
        RECT 32.685 177.525 32.855 177.695 ;
        RECT 33.605 177.525 33.775 177.695 ;
        RECT 34.065 177.865 34.235 178.035 ;
        RECT 34.985 177.525 35.155 177.695 ;
        RECT 35.905 177.525 36.075 177.695 ;
        RECT 31.765 176.845 31.935 177.015 ;
        RECT 40.045 178.545 40.215 178.715 ;
        RECT 40.965 178.545 41.135 178.715 ;
        RECT 39.125 177.185 39.295 177.355 ;
        RECT 38.665 176.845 38.835 177.015 ;
        RECT 43.725 178.205 43.895 178.375 ;
        RECT 41.885 177.525 42.055 177.695 ;
        RECT 42.805 177.525 42.975 177.695 ;
        RECT 40.125 176.845 40.295 177.015 ;
        RECT 44.185 177.525 44.355 177.695 ;
        RECT 45.105 176.845 45.275 177.015 ;
        RECT 47.865 177.525 48.035 177.695 ;
        RECT 46.945 176.845 47.115 177.015 ;
        RECT 50.165 177.525 50.335 177.695 ;
        RECT 51.085 177.525 51.255 177.695 ;
        RECT 52.465 177.525 52.635 177.695 ;
        RECT 51.775 177.185 51.945 177.355 ;
        RECT 49.245 176.845 49.415 177.015 ;
        RECT 53.845 177.185 54.015 177.355 ;
        RECT 58.445 178.545 58.615 178.715 ;
        RECT 60.745 178.545 60.915 178.715 ;
        RECT 54.765 177.525 54.935 177.695 ;
        RECT 55.225 177.525 55.395 177.695 ;
        RECT 59.365 178.205 59.535 178.375 ;
        RECT 56.145 177.525 56.315 177.695 ;
        RECT 52.925 176.845 53.095 177.015 ;
        RECT 57.525 177.185 57.695 177.355 ;
        RECT 58.525 176.845 58.695 177.015 ;
        RECT 59.825 177.185 59.995 177.355 ;
        RECT 60.825 177.185 60.995 177.355 ;
        RECT 61.665 176.845 61.835 177.015 ;
        RECT 62.585 177.525 62.755 177.695 ;
        RECT 71.350 178.205 71.520 178.375 ;
        RECT 63.965 176.845 64.135 177.015 ;
        RECT 70.405 177.525 70.575 177.695 ;
        RECT 70.865 177.525 71.035 177.695 ;
        RECT 69.945 176.845 70.115 177.015 ;
        RECT 71.745 177.865 71.915 178.035 ;
        RECT 72.200 177.185 72.370 177.355 ;
        RECT 73.450 178.205 73.620 178.375 ;
        RECT 72.935 177.865 73.105 178.035 ;
        RECT 75.020 178.205 75.190 178.375 ;
        RECT 75.455 177.865 75.625 178.035 ;
        RECT 77.765 178.205 77.935 178.375 ;
        RECT 78.225 178.545 78.395 178.715 ;
        RECT 80.985 177.865 81.155 178.035 ;
        RECT 83.285 176.845 83.455 177.015 ;
        RECT 86.045 177.865 86.215 178.035 ;
        RECT 87.425 177.525 87.595 177.695 ;
        RECT 85.585 176.845 85.755 177.015 ;
        RECT 88.345 177.525 88.515 177.695 ;
        RECT 87.885 176.845 88.055 177.015 ;
        RECT 18.425 176.335 18.595 176.505 ;
        RECT 18.885 176.335 19.055 176.505 ;
        RECT 19.345 176.335 19.515 176.505 ;
        RECT 19.805 176.335 19.975 176.505 ;
        RECT 20.265 176.335 20.435 176.505 ;
        RECT 20.725 176.335 20.895 176.505 ;
        RECT 21.185 176.335 21.355 176.505 ;
        RECT 21.645 176.335 21.815 176.505 ;
        RECT 22.105 176.335 22.275 176.505 ;
        RECT 22.565 176.335 22.735 176.505 ;
        RECT 23.025 176.335 23.195 176.505 ;
        RECT 23.485 176.335 23.655 176.505 ;
        RECT 23.945 176.335 24.115 176.505 ;
        RECT 24.405 176.335 24.575 176.505 ;
        RECT 24.865 176.335 25.035 176.505 ;
        RECT 25.325 176.335 25.495 176.505 ;
        RECT 25.785 176.335 25.955 176.505 ;
        RECT 26.245 176.335 26.415 176.505 ;
        RECT 26.705 176.335 26.875 176.505 ;
        RECT 27.165 176.335 27.335 176.505 ;
        RECT 27.625 176.335 27.795 176.505 ;
        RECT 28.085 176.335 28.255 176.505 ;
        RECT 28.545 176.335 28.715 176.505 ;
        RECT 29.005 176.335 29.175 176.505 ;
        RECT 29.465 176.335 29.635 176.505 ;
        RECT 29.925 176.335 30.095 176.505 ;
        RECT 30.385 176.335 30.555 176.505 ;
        RECT 30.845 176.335 31.015 176.505 ;
        RECT 31.305 176.335 31.475 176.505 ;
        RECT 31.765 176.335 31.935 176.505 ;
        RECT 32.225 176.335 32.395 176.505 ;
        RECT 32.685 176.335 32.855 176.505 ;
        RECT 33.145 176.335 33.315 176.505 ;
        RECT 33.605 176.335 33.775 176.505 ;
        RECT 34.065 176.335 34.235 176.505 ;
        RECT 34.525 176.335 34.695 176.505 ;
        RECT 34.985 176.335 35.155 176.505 ;
        RECT 35.445 176.335 35.615 176.505 ;
        RECT 35.905 176.335 36.075 176.505 ;
        RECT 36.365 176.335 36.535 176.505 ;
        RECT 36.825 176.335 36.995 176.505 ;
        RECT 37.285 176.335 37.455 176.505 ;
        RECT 37.745 176.335 37.915 176.505 ;
        RECT 38.205 176.335 38.375 176.505 ;
        RECT 38.665 176.335 38.835 176.505 ;
        RECT 39.125 176.335 39.295 176.505 ;
        RECT 39.585 176.335 39.755 176.505 ;
        RECT 40.045 176.335 40.215 176.505 ;
        RECT 40.505 176.335 40.675 176.505 ;
        RECT 40.965 176.335 41.135 176.505 ;
        RECT 41.425 176.335 41.595 176.505 ;
        RECT 41.885 176.335 42.055 176.505 ;
        RECT 42.345 176.335 42.515 176.505 ;
        RECT 42.805 176.335 42.975 176.505 ;
        RECT 43.265 176.335 43.435 176.505 ;
        RECT 43.725 176.335 43.895 176.505 ;
        RECT 44.185 176.335 44.355 176.505 ;
        RECT 44.645 176.335 44.815 176.505 ;
        RECT 45.105 176.335 45.275 176.505 ;
        RECT 45.565 176.335 45.735 176.505 ;
        RECT 46.025 176.335 46.195 176.505 ;
        RECT 46.485 176.335 46.655 176.505 ;
        RECT 46.945 176.335 47.115 176.505 ;
        RECT 47.405 176.335 47.575 176.505 ;
        RECT 47.865 176.335 48.035 176.505 ;
        RECT 48.325 176.335 48.495 176.505 ;
        RECT 48.785 176.335 48.955 176.505 ;
        RECT 49.245 176.335 49.415 176.505 ;
        RECT 49.705 176.335 49.875 176.505 ;
        RECT 50.165 176.335 50.335 176.505 ;
        RECT 50.625 176.335 50.795 176.505 ;
        RECT 51.085 176.335 51.255 176.505 ;
        RECT 51.545 176.335 51.715 176.505 ;
        RECT 52.005 176.335 52.175 176.505 ;
        RECT 52.465 176.335 52.635 176.505 ;
        RECT 52.925 176.335 53.095 176.505 ;
        RECT 53.385 176.335 53.555 176.505 ;
        RECT 53.845 176.335 54.015 176.505 ;
        RECT 54.305 176.335 54.475 176.505 ;
        RECT 54.765 176.335 54.935 176.505 ;
        RECT 55.225 176.335 55.395 176.505 ;
        RECT 55.685 176.335 55.855 176.505 ;
        RECT 56.145 176.335 56.315 176.505 ;
        RECT 56.605 176.335 56.775 176.505 ;
        RECT 57.065 176.335 57.235 176.505 ;
        RECT 57.525 176.335 57.695 176.505 ;
        RECT 57.985 176.335 58.155 176.505 ;
        RECT 58.445 176.335 58.615 176.505 ;
        RECT 58.905 176.335 59.075 176.505 ;
        RECT 59.365 176.335 59.535 176.505 ;
        RECT 59.825 176.335 59.995 176.505 ;
        RECT 60.285 176.335 60.455 176.505 ;
        RECT 60.745 176.335 60.915 176.505 ;
        RECT 61.205 176.335 61.375 176.505 ;
        RECT 61.665 176.335 61.835 176.505 ;
        RECT 62.125 176.335 62.295 176.505 ;
        RECT 62.585 176.335 62.755 176.505 ;
        RECT 63.045 176.335 63.215 176.505 ;
        RECT 63.505 176.335 63.675 176.505 ;
        RECT 63.965 176.335 64.135 176.505 ;
        RECT 64.425 176.335 64.595 176.505 ;
        RECT 64.885 176.335 65.055 176.505 ;
        RECT 65.345 176.335 65.515 176.505 ;
        RECT 65.805 176.335 65.975 176.505 ;
        RECT 66.265 176.335 66.435 176.505 ;
        RECT 66.725 176.335 66.895 176.505 ;
        RECT 67.185 176.335 67.355 176.505 ;
        RECT 67.645 176.335 67.815 176.505 ;
        RECT 68.105 176.335 68.275 176.505 ;
        RECT 68.565 176.335 68.735 176.505 ;
        RECT 69.025 176.335 69.195 176.505 ;
        RECT 69.485 176.335 69.655 176.505 ;
        RECT 69.945 176.335 70.115 176.505 ;
        RECT 70.405 176.335 70.575 176.505 ;
        RECT 70.865 176.335 71.035 176.505 ;
        RECT 71.325 176.335 71.495 176.505 ;
        RECT 71.785 176.335 71.955 176.505 ;
        RECT 72.245 176.335 72.415 176.505 ;
        RECT 72.705 176.335 72.875 176.505 ;
        RECT 73.165 176.335 73.335 176.505 ;
        RECT 73.625 176.335 73.795 176.505 ;
        RECT 74.085 176.335 74.255 176.505 ;
        RECT 74.545 176.335 74.715 176.505 ;
        RECT 75.005 176.335 75.175 176.505 ;
        RECT 75.465 176.335 75.635 176.505 ;
        RECT 75.925 176.335 76.095 176.505 ;
        RECT 76.385 176.335 76.555 176.505 ;
        RECT 76.845 176.335 77.015 176.505 ;
        RECT 77.305 176.335 77.475 176.505 ;
        RECT 77.765 176.335 77.935 176.505 ;
        RECT 78.225 176.335 78.395 176.505 ;
        RECT 78.685 176.335 78.855 176.505 ;
        RECT 79.145 176.335 79.315 176.505 ;
        RECT 79.605 176.335 79.775 176.505 ;
        RECT 80.065 176.335 80.235 176.505 ;
        RECT 80.525 176.335 80.695 176.505 ;
        RECT 80.985 176.335 81.155 176.505 ;
        RECT 81.445 176.335 81.615 176.505 ;
        RECT 81.905 176.335 82.075 176.505 ;
        RECT 82.365 176.335 82.535 176.505 ;
        RECT 82.825 176.335 82.995 176.505 ;
        RECT 83.285 176.335 83.455 176.505 ;
        RECT 83.745 176.335 83.915 176.505 ;
        RECT 84.205 176.335 84.375 176.505 ;
        RECT 84.665 176.335 84.835 176.505 ;
        RECT 85.125 176.335 85.295 176.505 ;
        RECT 85.585 176.335 85.755 176.505 ;
        RECT 86.045 176.335 86.215 176.505 ;
        RECT 86.505 176.335 86.675 176.505 ;
        RECT 86.965 176.335 87.135 176.505 ;
        RECT 87.425 176.335 87.595 176.505 ;
        RECT 87.885 176.335 88.055 176.505 ;
        RECT 88.345 176.335 88.515 176.505 ;
        RECT 88.805 176.335 88.975 176.505 ;
        RECT 89.265 176.335 89.435 176.505 ;
        RECT 89.725 176.335 89.895 176.505 ;
        RECT 90.185 176.335 90.355 176.505 ;
        RECT 90.645 176.335 90.815 176.505 ;
        RECT 91.105 176.335 91.275 176.505 ;
        RECT 91.565 176.335 91.735 176.505 ;
        RECT 92.025 176.335 92.195 176.505 ;
        RECT 25.325 174.125 25.495 174.295 ;
        RECT 32.225 175.825 32.395 175.995 ;
        RECT 28.545 174.805 28.715 174.975 ;
        RECT 31.765 175.145 31.935 175.315 ;
        RECT 32.685 175.145 32.855 175.315 ;
        RECT 35.445 175.825 35.615 175.995 ;
        RECT 34.985 175.145 35.155 175.315 ;
        RECT 35.905 175.145 36.075 175.315 ;
        RECT 40.045 175.825 40.215 175.995 ;
        RECT 39.585 175.145 39.755 175.315 ;
        RECT 44.645 174.805 44.815 174.975 ;
        RECT 45.130 174.465 45.300 174.635 ;
        RECT 45.525 174.805 45.695 174.975 ;
        RECT 45.980 175.485 46.150 175.655 ;
        RECT 46.715 174.805 46.885 174.975 ;
        RECT 47.230 174.465 47.400 174.635 ;
        RECT 48.800 174.465 48.970 174.635 ;
        RECT 49.235 174.805 49.405 174.975 ;
        RECT 51.545 175.825 51.715 175.995 ;
        RECT 52.005 175.485 52.175 175.655 ;
        RECT 58.445 175.825 58.615 175.995 ;
        RECT 61.205 175.145 61.375 175.315 ;
        RECT 61.665 175.145 61.835 175.315 ;
        RECT 62.585 175.145 62.755 175.315 ;
        RECT 63.505 175.485 63.675 175.655 ;
        RECT 63.965 175.145 64.135 175.315 ;
        RECT 64.885 175.145 65.055 175.315 ;
        RECT 65.345 175.145 65.515 175.315 ;
        RECT 65.805 175.145 65.975 175.315 ;
        RECT 67.645 175.145 67.815 175.315 ;
        RECT 68.565 175.825 68.735 175.995 ;
        RECT 69.025 175.145 69.195 175.315 ;
        RECT 67.185 174.125 67.355 174.295 ;
        RECT 67.645 174.125 67.815 174.295 ;
        RECT 70.405 174.805 70.575 174.975 ;
        RECT 74.085 175.825 74.255 175.995 ;
        RECT 75.005 175.145 75.175 175.315 ;
        RECT 75.465 174.465 75.635 174.635 ;
        RECT 76.385 175.145 76.555 175.315 ;
        RECT 77.305 175.145 77.475 175.315 ;
        RECT 78.225 175.145 78.395 175.315 ;
        RECT 79.145 175.145 79.315 175.315 ;
        RECT 80.985 175.145 81.155 175.315 ;
        RECT 81.905 175.145 82.075 175.315 ;
        RECT 75.925 174.465 76.095 174.635 ;
        RECT 79.605 174.805 79.775 174.975 ;
        RECT 82.365 174.805 82.535 174.975 ;
        RECT 82.830 174.465 83.000 174.635 ;
        RECT 83.290 175.485 83.460 175.655 ;
        RECT 83.745 175.145 83.915 175.315 ;
        RECT 84.690 175.485 84.860 175.655 ;
        RECT 86.530 175.485 86.700 175.655 ;
        RECT 85.150 174.465 85.320 174.635 ;
        RECT 86.530 174.465 86.700 174.635 ;
        RECT 90.185 174.125 90.355 174.295 ;
        RECT 18.425 173.615 18.595 173.785 ;
        RECT 18.885 173.615 19.055 173.785 ;
        RECT 19.345 173.615 19.515 173.785 ;
        RECT 19.805 173.615 19.975 173.785 ;
        RECT 20.265 173.615 20.435 173.785 ;
        RECT 20.725 173.615 20.895 173.785 ;
        RECT 21.185 173.615 21.355 173.785 ;
        RECT 21.645 173.615 21.815 173.785 ;
        RECT 22.105 173.615 22.275 173.785 ;
        RECT 22.565 173.615 22.735 173.785 ;
        RECT 23.025 173.615 23.195 173.785 ;
        RECT 23.485 173.615 23.655 173.785 ;
        RECT 23.945 173.615 24.115 173.785 ;
        RECT 24.405 173.615 24.575 173.785 ;
        RECT 24.865 173.615 25.035 173.785 ;
        RECT 25.325 173.615 25.495 173.785 ;
        RECT 25.785 173.615 25.955 173.785 ;
        RECT 26.245 173.615 26.415 173.785 ;
        RECT 26.705 173.615 26.875 173.785 ;
        RECT 27.165 173.615 27.335 173.785 ;
        RECT 27.625 173.615 27.795 173.785 ;
        RECT 28.085 173.615 28.255 173.785 ;
        RECT 28.545 173.615 28.715 173.785 ;
        RECT 29.005 173.615 29.175 173.785 ;
        RECT 29.465 173.615 29.635 173.785 ;
        RECT 29.925 173.615 30.095 173.785 ;
        RECT 30.385 173.615 30.555 173.785 ;
        RECT 30.845 173.615 31.015 173.785 ;
        RECT 31.305 173.615 31.475 173.785 ;
        RECT 31.765 173.615 31.935 173.785 ;
        RECT 32.225 173.615 32.395 173.785 ;
        RECT 32.685 173.615 32.855 173.785 ;
        RECT 33.145 173.615 33.315 173.785 ;
        RECT 33.605 173.615 33.775 173.785 ;
        RECT 34.065 173.615 34.235 173.785 ;
        RECT 34.525 173.615 34.695 173.785 ;
        RECT 34.985 173.615 35.155 173.785 ;
        RECT 35.445 173.615 35.615 173.785 ;
        RECT 35.905 173.615 36.075 173.785 ;
        RECT 36.365 173.615 36.535 173.785 ;
        RECT 36.825 173.615 36.995 173.785 ;
        RECT 37.285 173.615 37.455 173.785 ;
        RECT 37.745 173.615 37.915 173.785 ;
        RECT 38.205 173.615 38.375 173.785 ;
        RECT 38.665 173.615 38.835 173.785 ;
        RECT 39.125 173.615 39.295 173.785 ;
        RECT 39.585 173.615 39.755 173.785 ;
        RECT 40.045 173.615 40.215 173.785 ;
        RECT 40.505 173.615 40.675 173.785 ;
        RECT 40.965 173.615 41.135 173.785 ;
        RECT 41.425 173.615 41.595 173.785 ;
        RECT 41.885 173.615 42.055 173.785 ;
        RECT 42.345 173.615 42.515 173.785 ;
        RECT 42.805 173.615 42.975 173.785 ;
        RECT 43.265 173.615 43.435 173.785 ;
        RECT 43.725 173.615 43.895 173.785 ;
        RECT 44.185 173.615 44.355 173.785 ;
        RECT 44.645 173.615 44.815 173.785 ;
        RECT 45.105 173.615 45.275 173.785 ;
        RECT 45.565 173.615 45.735 173.785 ;
        RECT 46.025 173.615 46.195 173.785 ;
        RECT 46.485 173.615 46.655 173.785 ;
        RECT 46.945 173.615 47.115 173.785 ;
        RECT 47.405 173.615 47.575 173.785 ;
        RECT 47.865 173.615 48.035 173.785 ;
        RECT 48.325 173.615 48.495 173.785 ;
        RECT 48.785 173.615 48.955 173.785 ;
        RECT 49.245 173.615 49.415 173.785 ;
        RECT 49.705 173.615 49.875 173.785 ;
        RECT 50.165 173.615 50.335 173.785 ;
        RECT 50.625 173.615 50.795 173.785 ;
        RECT 51.085 173.615 51.255 173.785 ;
        RECT 51.545 173.615 51.715 173.785 ;
        RECT 52.005 173.615 52.175 173.785 ;
        RECT 52.465 173.615 52.635 173.785 ;
        RECT 52.925 173.615 53.095 173.785 ;
        RECT 53.385 173.615 53.555 173.785 ;
        RECT 53.845 173.615 54.015 173.785 ;
        RECT 54.305 173.615 54.475 173.785 ;
        RECT 54.765 173.615 54.935 173.785 ;
        RECT 55.225 173.615 55.395 173.785 ;
        RECT 55.685 173.615 55.855 173.785 ;
        RECT 56.145 173.615 56.315 173.785 ;
        RECT 56.605 173.615 56.775 173.785 ;
        RECT 57.065 173.615 57.235 173.785 ;
        RECT 57.525 173.615 57.695 173.785 ;
        RECT 57.985 173.615 58.155 173.785 ;
        RECT 58.445 173.615 58.615 173.785 ;
        RECT 58.905 173.615 59.075 173.785 ;
        RECT 59.365 173.615 59.535 173.785 ;
        RECT 59.825 173.615 59.995 173.785 ;
        RECT 60.285 173.615 60.455 173.785 ;
        RECT 60.745 173.615 60.915 173.785 ;
        RECT 61.205 173.615 61.375 173.785 ;
        RECT 61.665 173.615 61.835 173.785 ;
        RECT 62.125 173.615 62.295 173.785 ;
        RECT 62.585 173.615 62.755 173.785 ;
        RECT 63.045 173.615 63.215 173.785 ;
        RECT 63.505 173.615 63.675 173.785 ;
        RECT 63.965 173.615 64.135 173.785 ;
        RECT 64.425 173.615 64.595 173.785 ;
        RECT 64.885 173.615 65.055 173.785 ;
        RECT 65.345 173.615 65.515 173.785 ;
        RECT 65.805 173.615 65.975 173.785 ;
        RECT 66.265 173.615 66.435 173.785 ;
        RECT 66.725 173.615 66.895 173.785 ;
        RECT 67.185 173.615 67.355 173.785 ;
        RECT 67.645 173.615 67.815 173.785 ;
        RECT 68.105 173.615 68.275 173.785 ;
        RECT 68.565 173.615 68.735 173.785 ;
        RECT 69.025 173.615 69.195 173.785 ;
        RECT 69.485 173.615 69.655 173.785 ;
        RECT 69.945 173.615 70.115 173.785 ;
        RECT 70.405 173.615 70.575 173.785 ;
        RECT 70.865 173.615 71.035 173.785 ;
        RECT 71.325 173.615 71.495 173.785 ;
        RECT 71.785 173.615 71.955 173.785 ;
        RECT 72.245 173.615 72.415 173.785 ;
        RECT 72.705 173.615 72.875 173.785 ;
        RECT 73.165 173.615 73.335 173.785 ;
        RECT 73.625 173.615 73.795 173.785 ;
        RECT 74.085 173.615 74.255 173.785 ;
        RECT 74.545 173.615 74.715 173.785 ;
        RECT 75.005 173.615 75.175 173.785 ;
        RECT 75.465 173.615 75.635 173.785 ;
        RECT 75.925 173.615 76.095 173.785 ;
        RECT 76.385 173.615 76.555 173.785 ;
        RECT 76.845 173.615 77.015 173.785 ;
        RECT 77.305 173.615 77.475 173.785 ;
        RECT 77.765 173.615 77.935 173.785 ;
        RECT 78.225 173.615 78.395 173.785 ;
        RECT 78.685 173.615 78.855 173.785 ;
        RECT 79.145 173.615 79.315 173.785 ;
        RECT 79.605 173.615 79.775 173.785 ;
        RECT 80.065 173.615 80.235 173.785 ;
        RECT 80.525 173.615 80.695 173.785 ;
        RECT 80.985 173.615 81.155 173.785 ;
        RECT 81.445 173.615 81.615 173.785 ;
        RECT 81.905 173.615 82.075 173.785 ;
        RECT 82.365 173.615 82.535 173.785 ;
        RECT 82.825 173.615 82.995 173.785 ;
        RECT 83.285 173.615 83.455 173.785 ;
        RECT 83.745 173.615 83.915 173.785 ;
        RECT 84.205 173.615 84.375 173.785 ;
        RECT 84.665 173.615 84.835 173.785 ;
        RECT 85.125 173.615 85.295 173.785 ;
        RECT 85.585 173.615 85.755 173.785 ;
        RECT 86.045 173.615 86.215 173.785 ;
        RECT 86.505 173.615 86.675 173.785 ;
        RECT 86.965 173.615 87.135 173.785 ;
        RECT 87.425 173.615 87.595 173.785 ;
        RECT 87.885 173.615 88.055 173.785 ;
        RECT 88.345 173.615 88.515 173.785 ;
        RECT 88.805 173.615 88.975 173.785 ;
        RECT 89.265 173.615 89.435 173.785 ;
        RECT 89.725 173.615 89.895 173.785 ;
        RECT 90.185 173.615 90.355 173.785 ;
        RECT 90.645 173.615 90.815 173.785 ;
        RECT 91.105 173.615 91.275 173.785 ;
        RECT 91.565 173.615 91.735 173.785 ;
        RECT 92.025 173.615 92.195 173.785 ;
        RECT 23.510 172.765 23.680 172.935 ;
        RECT 23.025 172.085 23.195 172.255 ;
        RECT 23.905 172.425 24.075 172.595 ;
        RECT 24.360 171.745 24.530 171.915 ;
        RECT 25.610 172.765 25.780 172.935 ;
        RECT 25.095 172.425 25.265 172.595 ;
        RECT 27.180 172.765 27.350 172.935 ;
        RECT 27.615 172.425 27.785 172.595 ;
        RECT 29.925 173.105 30.095 173.275 ;
        RECT 31.765 172.765 31.935 172.935 ;
        RECT 31.765 171.745 31.935 171.915 ;
        RECT 33.145 172.085 33.315 172.255 ;
        RECT 35.445 172.765 35.615 172.935 ;
        RECT 37.745 173.105 37.915 173.275 ;
        RECT 32.685 171.405 32.855 171.575 ;
        RECT 36.825 172.425 36.995 172.595 ;
        RECT 38.665 172.765 38.835 172.935 ;
        RECT 38.205 172.085 38.375 172.255 ;
        RECT 41.425 173.105 41.595 173.275 ;
        RECT 39.585 171.405 39.755 171.575 ;
        RECT 40.045 171.405 40.215 171.575 ;
        RECT 40.505 172.085 40.675 172.255 ;
        RECT 42.805 172.085 42.975 172.255 ;
        RECT 43.725 171.405 43.895 171.575 ;
        RECT 46.945 173.105 47.115 173.275 ;
        RECT 48.785 172.425 48.955 172.595 ;
        RECT 47.865 172.085 48.035 172.255 ;
        RECT 58.905 172.765 59.075 172.935 ;
        RECT 58.445 172.085 58.615 172.255 ;
        RECT 59.365 172.085 59.535 172.255 ;
        RECT 59.825 172.085 59.995 172.255 ;
        RECT 62.585 172.765 62.755 172.935 ;
        RECT 60.745 172.085 60.915 172.255 ;
        RECT 61.205 172.085 61.375 172.255 ;
        RECT 57.525 171.405 57.695 171.575 ;
        RECT 65.370 172.765 65.540 172.935 ;
        RECT 61.665 171.405 61.835 171.575 ;
        RECT 62.585 171.745 62.755 171.915 ;
        RECT 64.885 172.425 65.055 172.595 ;
        RECT 63.505 172.085 63.675 172.255 ;
        RECT 63.965 172.085 64.135 172.255 ;
        RECT 65.765 172.425 65.935 172.595 ;
        RECT 66.220 172.085 66.390 172.255 ;
        RECT 67.470 172.765 67.640 172.935 ;
        RECT 66.955 172.425 67.125 172.595 ;
        RECT 69.040 172.765 69.210 172.935 ;
        RECT 69.475 172.425 69.645 172.595 ;
        RECT 71.785 173.105 71.955 173.275 ;
        RECT 81.445 173.105 81.615 173.275 ;
        RECT 81.445 172.085 81.615 172.255 ;
        RECT 83.745 172.425 83.915 172.595 ;
        RECT 82.365 172.085 82.535 172.255 ;
        RECT 83.285 172.085 83.455 172.255 ;
        RECT 84.205 172.085 84.375 172.255 ;
        RECT 18.425 170.895 18.595 171.065 ;
        RECT 18.885 170.895 19.055 171.065 ;
        RECT 19.345 170.895 19.515 171.065 ;
        RECT 19.805 170.895 19.975 171.065 ;
        RECT 20.265 170.895 20.435 171.065 ;
        RECT 20.725 170.895 20.895 171.065 ;
        RECT 21.185 170.895 21.355 171.065 ;
        RECT 21.645 170.895 21.815 171.065 ;
        RECT 22.105 170.895 22.275 171.065 ;
        RECT 22.565 170.895 22.735 171.065 ;
        RECT 23.025 170.895 23.195 171.065 ;
        RECT 23.485 170.895 23.655 171.065 ;
        RECT 23.945 170.895 24.115 171.065 ;
        RECT 24.405 170.895 24.575 171.065 ;
        RECT 24.865 170.895 25.035 171.065 ;
        RECT 25.325 170.895 25.495 171.065 ;
        RECT 25.785 170.895 25.955 171.065 ;
        RECT 26.245 170.895 26.415 171.065 ;
        RECT 26.705 170.895 26.875 171.065 ;
        RECT 27.165 170.895 27.335 171.065 ;
        RECT 27.625 170.895 27.795 171.065 ;
        RECT 28.085 170.895 28.255 171.065 ;
        RECT 28.545 170.895 28.715 171.065 ;
        RECT 29.005 170.895 29.175 171.065 ;
        RECT 29.465 170.895 29.635 171.065 ;
        RECT 29.925 170.895 30.095 171.065 ;
        RECT 30.385 170.895 30.555 171.065 ;
        RECT 30.845 170.895 31.015 171.065 ;
        RECT 31.305 170.895 31.475 171.065 ;
        RECT 31.765 170.895 31.935 171.065 ;
        RECT 32.225 170.895 32.395 171.065 ;
        RECT 32.685 170.895 32.855 171.065 ;
        RECT 33.145 170.895 33.315 171.065 ;
        RECT 33.605 170.895 33.775 171.065 ;
        RECT 34.065 170.895 34.235 171.065 ;
        RECT 34.525 170.895 34.695 171.065 ;
        RECT 34.985 170.895 35.155 171.065 ;
        RECT 35.445 170.895 35.615 171.065 ;
        RECT 35.905 170.895 36.075 171.065 ;
        RECT 36.365 170.895 36.535 171.065 ;
        RECT 36.825 170.895 36.995 171.065 ;
        RECT 37.285 170.895 37.455 171.065 ;
        RECT 37.745 170.895 37.915 171.065 ;
        RECT 38.205 170.895 38.375 171.065 ;
        RECT 38.665 170.895 38.835 171.065 ;
        RECT 39.125 170.895 39.295 171.065 ;
        RECT 39.585 170.895 39.755 171.065 ;
        RECT 40.045 170.895 40.215 171.065 ;
        RECT 40.505 170.895 40.675 171.065 ;
        RECT 40.965 170.895 41.135 171.065 ;
        RECT 41.425 170.895 41.595 171.065 ;
        RECT 41.885 170.895 42.055 171.065 ;
        RECT 42.345 170.895 42.515 171.065 ;
        RECT 42.805 170.895 42.975 171.065 ;
        RECT 43.265 170.895 43.435 171.065 ;
        RECT 43.725 170.895 43.895 171.065 ;
        RECT 44.185 170.895 44.355 171.065 ;
        RECT 44.645 170.895 44.815 171.065 ;
        RECT 45.105 170.895 45.275 171.065 ;
        RECT 45.565 170.895 45.735 171.065 ;
        RECT 46.025 170.895 46.195 171.065 ;
        RECT 46.485 170.895 46.655 171.065 ;
        RECT 46.945 170.895 47.115 171.065 ;
        RECT 47.405 170.895 47.575 171.065 ;
        RECT 47.865 170.895 48.035 171.065 ;
        RECT 48.325 170.895 48.495 171.065 ;
        RECT 48.785 170.895 48.955 171.065 ;
        RECT 49.245 170.895 49.415 171.065 ;
        RECT 49.705 170.895 49.875 171.065 ;
        RECT 50.165 170.895 50.335 171.065 ;
        RECT 50.625 170.895 50.795 171.065 ;
        RECT 51.085 170.895 51.255 171.065 ;
        RECT 51.545 170.895 51.715 171.065 ;
        RECT 52.005 170.895 52.175 171.065 ;
        RECT 52.465 170.895 52.635 171.065 ;
        RECT 52.925 170.895 53.095 171.065 ;
        RECT 53.385 170.895 53.555 171.065 ;
        RECT 53.845 170.895 54.015 171.065 ;
        RECT 54.305 170.895 54.475 171.065 ;
        RECT 54.765 170.895 54.935 171.065 ;
        RECT 55.225 170.895 55.395 171.065 ;
        RECT 55.685 170.895 55.855 171.065 ;
        RECT 56.145 170.895 56.315 171.065 ;
        RECT 56.605 170.895 56.775 171.065 ;
        RECT 57.065 170.895 57.235 171.065 ;
        RECT 57.525 170.895 57.695 171.065 ;
        RECT 57.985 170.895 58.155 171.065 ;
        RECT 58.445 170.895 58.615 171.065 ;
        RECT 58.905 170.895 59.075 171.065 ;
        RECT 59.365 170.895 59.535 171.065 ;
        RECT 59.825 170.895 59.995 171.065 ;
        RECT 60.285 170.895 60.455 171.065 ;
        RECT 60.745 170.895 60.915 171.065 ;
        RECT 61.205 170.895 61.375 171.065 ;
        RECT 61.665 170.895 61.835 171.065 ;
        RECT 62.125 170.895 62.295 171.065 ;
        RECT 62.585 170.895 62.755 171.065 ;
        RECT 63.045 170.895 63.215 171.065 ;
        RECT 63.505 170.895 63.675 171.065 ;
        RECT 63.965 170.895 64.135 171.065 ;
        RECT 64.425 170.895 64.595 171.065 ;
        RECT 64.885 170.895 65.055 171.065 ;
        RECT 65.345 170.895 65.515 171.065 ;
        RECT 65.805 170.895 65.975 171.065 ;
        RECT 66.265 170.895 66.435 171.065 ;
        RECT 66.725 170.895 66.895 171.065 ;
        RECT 67.185 170.895 67.355 171.065 ;
        RECT 67.645 170.895 67.815 171.065 ;
        RECT 68.105 170.895 68.275 171.065 ;
        RECT 68.565 170.895 68.735 171.065 ;
        RECT 69.025 170.895 69.195 171.065 ;
        RECT 69.485 170.895 69.655 171.065 ;
        RECT 69.945 170.895 70.115 171.065 ;
        RECT 70.405 170.895 70.575 171.065 ;
        RECT 70.865 170.895 71.035 171.065 ;
        RECT 71.325 170.895 71.495 171.065 ;
        RECT 71.785 170.895 71.955 171.065 ;
        RECT 72.245 170.895 72.415 171.065 ;
        RECT 72.705 170.895 72.875 171.065 ;
        RECT 73.165 170.895 73.335 171.065 ;
        RECT 73.625 170.895 73.795 171.065 ;
        RECT 74.085 170.895 74.255 171.065 ;
        RECT 74.545 170.895 74.715 171.065 ;
        RECT 75.005 170.895 75.175 171.065 ;
        RECT 75.465 170.895 75.635 171.065 ;
        RECT 75.925 170.895 76.095 171.065 ;
        RECT 76.385 170.895 76.555 171.065 ;
        RECT 76.845 170.895 77.015 171.065 ;
        RECT 77.305 170.895 77.475 171.065 ;
        RECT 77.765 170.895 77.935 171.065 ;
        RECT 78.225 170.895 78.395 171.065 ;
        RECT 78.685 170.895 78.855 171.065 ;
        RECT 79.145 170.895 79.315 171.065 ;
        RECT 79.605 170.895 79.775 171.065 ;
        RECT 80.065 170.895 80.235 171.065 ;
        RECT 80.525 170.895 80.695 171.065 ;
        RECT 80.985 170.895 81.155 171.065 ;
        RECT 81.445 170.895 81.615 171.065 ;
        RECT 81.905 170.895 82.075 171.065 ;
        RECT 82.365 170.895 82.535 171.065 ;
        RECT 82.825 170.895 82.995 171.065 ;
        RECT 83.285 170.895 83.455 171.065 ;
        RECT 83.745 170.895 83.915 171.065 ;
        RECT 84.205 170.895 84.375 171.065 ;
        RECT 84.665 170.895 84.835 171.065 ;
        RECT 85.125 170.895 85.295 171.065 ;
        RECT 85.585 170.895 85.755 171.065 ;
        RECT 86.045 170.895 86.215 171.065 ;
        RECT 86.505 170.895 86.675 171.065 ;
        RECT 86.965 170.895 87.135 171.065 ;
        RECT 87.425 170.895 87.595 171.065 ;
        RECT 87.885 170.895 88.055 171.065 ;
        RECT 88.345 170.895 88.515 171.065 ;
        RECT 88.805 170.895 88.975 171.065 ;
        RECT 89.265 170.895 89.435 171.065 ;
        RECT 89.725 170.895 89.895 171.065 ;
        RECT 90.185 170.895 90.355 171.065 ;
        RECT 90.645 170.895 90.815 171.065 ;
        RECT 91.105 170.895 91.275 171.065 ;
        RECT 91.565 170.895 91.735 171.065 ;
        RECT 92.025 170.895 92.195 171.065 ;
        RECT 28.085 170.385 28.255 170.555 ;
        RECT 27.165 169.705 27.335 169.875 ;
        RECT 28.085 169.705 28.255 169.875 ;
        RECT 37.285 170.045 37.455 170.215 ;
        RECT 30.845 169.025 31.015 169.195 ;
        RECT 38.205 169.365 38.375 169.535 ;
        RECT 38.665 169.365 38.835 169.535 ;
        RECT 39.125 169.705 39.295 169.875 ;
        RECT 39.585 169.365 39.755 169.535 ;
        RECT 40.505 168.685 40.675 168.855 ;
        RECT 52.465 169.705 52.635 169.875 ;
        RECT 52.950 169.025 53.120 169.195 ;
        RECT 53.345 169.365 53.515 169.535 ;
        RECT 53.800 169.705 53.970 169.875 ;
        RECT 54.535 169.365 54.705 169.535 ;
        RECT 55.050 169.025 55.220 169.195 ;
        RECT 56.620 169.025 56.790 169.195 ;
        RECT 57.055 169.365 57.225 169.535 ;
        RECT 59.365 170.385 59.535 170.555 ;
        RECT 59.825 169.705 59.995 169.875 ;
        RECT 60.745 169.705 60.915 169.875 ;
        RECT 60.285 169.025 60.455 169.195 ;
        RECT 75.005 169.365 75.175 169.535 ;
        RECT 75.465 169.705 75.635 169.875 ;
        RECT 75.925 169.365 76.095 169.535 ;
        RECT 76.385 169.365 76.555 169.535 ;
        RECT 77.305 168.685 77.475 168.855 ;
        RECT 81.445 170.045 81.615 170.215 ;
        RECT 79.605 169.705 79.775 169.875 ;
        RECT 80.065 169.705 80.235 169.875 ;
        RECT 80.805 169.705 80.975 169.875 ;
        RECT 81.905 169.705 82.075 169.875 ;
        RECT 79.145 169.365 79.315 169.535 ;
        RECT 77.765 169.025 77.935 169.195 ;
        RECT 78.685 168.685 78.855 168.855 ;
        RECT 83.285 168.685 83.455 168.855 ;
        RECT 18.425 168.175 18.595 168.345 ;
        RECT 18.885 168.175 19.055 168.345 ;
        RECT 19.345 168.175 19.515 168.345 ;
        RECT 19.805 168.175 19.975 168.345 ;
        RECT 20.265 168.175 20.435 168.345 ;
        RECT 20.725 168.175 20.895 168.345 ;
        RECT 21.185 168.175 21.355 168.345 ;
        RECT 21.645 168.175 21.815 168.345 ;
        RECT 22.105 168.175 22.275 168.345 ;
        RECT 22.565 168.175 22.735 168.345 ;
        RECT 23.025 168.175 23.195 168.345 ;
        RECT 23.485 168.175 23.655 168.345 ;
        RECT 23.945 168.175 24.115 168.345 ;
        RECT 24.405 168.175 24.575 168.345 ;
        RECT 24.865 168.175 25.035 168.345 ;
        RECT 25.325 168.175 25.495 168.345 ;
        RECT 25.785 168.175 25.955 168.345 ;
        RECT 26.245 168.175 26.415 168.345 ;
        RECT 26.705 168.175 26.875 168.345 ;
        RECT 27.165 168.175 27.335 168.345 ;
        RECT 27.625 168.175 27.795 168.345 ;
        RECT 28.085 168.175 28.255 168.345 ;
        RECT 28.545 168.175 28.715 168.345 ;
        RECT 29.005 168.175 29.175 168.345 ;
        RECT 29.465 168.175 29.635 168.345 ;
        RECT 29.925 168.175 30.095 168.345 ;
        RECT 30.385 168.175 30.555 168.345 ;
        RECT 30.845 168.175 31.015 168.345 ;
        RECT 31.305 168.175 31.475 168.345 ;
        RECT 31.765 168.175 31.935 168.345 ;
        RECT 32.225 168.175 32.395 168.345 ;
        RECT 32.685 168.175 32.855 168.345 ;
        RECT 33.145 168.175 33.315 168.345 ;
        RECT 33.605 168.175 33.775 168.345 ;
        RECT 34.065 168.175 34.235 168.345 ;
        RECT 34.525 168.175 34.695 168.345 ;
        RECT 34.985 168.175 35.155 168.345 ;
        RECT 35.445 168.175 35.615 168.345 ;
        RECT 35.905 168.175 36.075 168.345 ;
        RECT 36.365 168.175 36.535 168.345 ;
        RECT 36.825 168.175 36.995 168.345 ;
        RECT 37.285 168.175 37.455 168.345 ;
        RECT 37.745 168.175 37.915 168.345 ;
        RECT 38.205 168.175 38.375 168.345 ;
        RECT 38.665 168.175 38.835 168.345 ;
        RECT 39.125 168.175 39.295 168.345 ;
        RECT 39.585 168.175 39.755 168.345 ;
        RECT 40.045 168.175 40.215 168.345 ;
        RECT 40.505 168.175 40.675 168.345 ;
        RECT 40.965 168.175 41.135 168.345 ;
        RECT 41.425 168.175 41.595 168.345 ;
        RECT 41.885 168.175 42.055 168.345 ;
        RECT 42.345 168.175 42.515 168.345 ;
        RECT 42.805 168.175 42.975 168.345 ;
        RECT 43.265 168.175 43.435 168.345 ;
        RECT 43.725 168.175 43.895 168.345 ;
        RECT 44.185 168.175 44.355 168.345 ;
        RECT 44.645 168.175 44.815 168.345 ;
        RECT 45.105 168.175 45.275 168.345 ;
        RECT 45.565 168.175 45.735 168.345 ;
        RECT 46.025 168.175 46.195 168.345 ;
        RECT 46.485 168.175 46.655 168.345 ;
        RECT 46.945 168.175 47.115 168.345 ;
        RECT 47.405 168.175 47.575 168.345 ;
        RECT 47.865 168.175 48.035 168.345 ;
        RECT 48.325 168.175 48.495 168.345 ;
        RECT 48.785 168.175 48.955 168.345 ;
        RECT 49.245 168.175 49.415 168.345 ;
        RECT 49.705 168.175 49.875 168.345 ;
        RECT 50.165 168.175 50.335 168.345 ;
        RECT 50.625 168.175 50.795 168.345 ;
        RECT 51.085 168.175 51.255 168.345 ;
        RECT 51.545 168.175 51.715 168.345 ;
        RECT 52.005 168.175 52.175 168.345 ;
        RECT 52.465 168.175 52.635 168.345 ;
        RECT 52.925 168.175 53.095 168.345 ;
        RECT 53.385 168.175 53.555 168.345 ;
        RECT 53.845 168.175 54.015 168.345 ;
        RECT 54.305 168.175 54.475 168.345 ;
        RECT 54.765 168.175 54.935 168.345 ;
        RECT 55.225 168.175 55.395 168.345 ;
        RECT 55.685 168.175 55.855 168.345 ;
        RECT 56.145 168.175 56.315 168.345 ;
        RECT 56.605 168.175 56.775 168.345 ;
        RECT 57.065 168.175 57.235 168.345 ;
        RECT 57.525 168.175 57.695 168.345 ;
        RECT 57.985 168.175 58.155 168.345 ;
        RECT 58.445 168.175 58.615 168.345 ;
        RECT 58.905 168.175 59.075 168.345 ;
        RECT 59.365 168.175 59.535 168.345 ;
        RECT 59.825 168.175 59.995 168.345 ;
        RECT 60.285 168.175 60.455 168.345 ;
        RECT 60.745 168.175 60.915 168.345 ;
        RECT 61.205 168.175 61.375 168.345 ;
        RECT 61.665 168.175 61.835 168.345 ;
        RECT 62.125 168.175 62.295 168.345 ;
        RECT 62.585 168.175 62.755 168.345 ;
        RECT 63.045 168.175 63.215 168.345 ;
        RECT 63.505 168.175 63.675 168.345 ;
        RECT 63.965 168.175 64.135 168.345 ;
        RECT 64.425 168.175 64.595 168.345 ;
        RECT 64.885 168.175 65.055 168.345 ;
        RECT 65.345 168.175 65.515 168.345 ;
        RECT 65.805 168.175 65.975 168.345 ;
        RECT 66.265 168.175 66.435 168.345 ;
        RECT 66.725 168.175 66.895 168.345 ;
        RECT 67.185 168.175 67.355 168.345 ;
        RECT 67.645 168.175 67.815 168.345 ;
        RECT 68.105 168.175 68.275 168.345 ;
        RECT 68.565 168.175 68.735 168.345 ;
        RECT 69.025 168.175 69.195 168.345 ;
        RECT 69.485 168.175 69.655 168.345 ;
        RECT 69.945 168.175 70.115 168.345 ;
        RECT 70.405 168.175 70.575 168.345 ;
        RECT 70.865 168.175 71.035 168.345 ;
        RECT 71.325 168.175 71.495 168.345 ;
        RECT 71.785 168.175 71.955 168.345 ;
        RECT 72.245 168.175 72.415 168.345 ;
        RECT 72.705 168.175 72.875 168.345 ;
        RECT 73.165 168.175 73.335 168.345 ;
        RECT 73.625 168.175 73.795 168.345 ;
        RECT 74.085 168.175 74.255 168.345 ;
        RECT 74.545 168.175 74.715 168.345 ;
        RECT 75.005 168.175 75.175 168.345 ;
        RECT 75.465 168.175 75.635 168.345 ;
        RECT 75.925 168.175 76.095 168.345 ;
        RECT 76.385 168.175 76.555 168.345 ;
        RECT 76.845 168.175 77.015 168.345 ;
        RECT 77.305 168.175 77.475 168.345 ;
        RECT 77.765 168.175 77.935 168.345 ;
        RECT 78.225 168.175 78.395 168.345 ;
        RECT 78.685 168.175 78.855 168.345 ;
        RECT 79.145 168.175 79.315 168.345 ;
        RECT 79.605 168.175 79.775 168.345 ;
        RECT 80.065 168.175 80.235 168.345 ;
        RECT 80.525 168.175 80.695 168.345 ;
        RECT 80.985 168.175 81.155 168.345 ;
        RECT 81.445 168.175 81.615 168.345 ;
        RECT 81.905 168.175 82.075 168.345 ;
        RECT 82.365 168.175 82.535 168.345 ;
        RECT 82.825 168.175 82.995 168.345 ;
        RECT 83.285 168.175 83.455 168.345 ;
        RECT 83.745 168.175 83.915 168.345 ;
        RECT 84.205 168.175 84.375 168.345 ;
        RECT 84.665 168.175 84.835 168.345 ;
        RECT 85.125 168.175 85.295 168.345 ;
        RECT 85.585 168.175 85.755 168.345 ;
        RECT 86.045 168.175 86.215 168.345 ;
        RECT 86.505 168.175 86.675 168.345 ;
        RECT 86.965 168.175 87.135 168.345 ;
        RECT 87.425 168.175 87.595 168.345 ;
        RECT 87.885 168.175 88.055 168.345 ;
        RECT 88.345 168.175 88.515 168.345 ;
        RECT 88.805 168.175 88.975 168.345 ;
        RECT 89.265 168.175 89.435 168.345 ;
        RECT 89.725 168.175 89.895 168.345 ;
        RECT 90.185 168.175 90.355 168.345 ;
        RECT 90.645 168.175 90.815 168.345 ;
        RECT 91.105 168.175 91.275 168.345 ;
        RECT 91.565 168.175 91.735 168.345 ;
        RECT 92.025 168.175 92.195 168.345 ;
        RECT 34.525 167.325 34.695 167.495 ;
        RECT 37.285 167.665 37.455 167.835 ;
        RECT 35.445 165.965 35.615 166.135 ;
        RECT 35.905 166.305 36.075 166.475 ;
        RECT 36.365 165.965 36.535 166.135 ;
        RECT 39.585 167.665 39.755 167.835 ;
        RECT 37.745 166.985 37.915 167.155 ;
        RECT 38.665 166.645 38.835 166.815 ;
        RECT 40.990 167.325 41.160 167.495 ;
        RECT 40.505 166.645 40.675 166.815 ;
        RECT 41.385 166.985 41.555 167.155 ;
        RECT 41.840 166.305 42.010 166.475 ;
        RECT 43.090 167.325 43.260 167.495 ;
        RECT 42.575 166.985 42.745 167.155 ;
        RECT 44.660 167.325 44.830 167.495 ;
        RECT 45.095 166.985 45.265 167.155 ;
        RECT 47.405 167.325 47.575 167.495 ;
        RECT 49.705 166.985 49.875 167.155 ;
        RECT 52.925 166.985 53.095 167.155 ;
        RECT 54.765 167.665 54.935 167.835 ;
        RECT 53.845 166.645 54.015 166.815 ;
        RECT 54.765 166.645 54.935 166.815 ;
        RECT 55.225 166.645 55.395 166.815 ;
        RECT 55.685 165.965 55.855 166.135 ;
        RECT 63.965 167.325 64.135 167.495 ;
        RECT 64.885 167.325 65.055 167.495 ;
        RECT 62.585 166.645 62.755 166.815 ;
        RECT 66.265 167.325 66.435 167.495 ;
        RECT 63.045 165.965 63.215 166.135 ;
        RECT 63.965 166.645 64.135 166.815 ;
        RECT 64.425 166.645 64.595 166.815 ;
        RECT 65.805 166.985 65.975 167.155 ;
        RECT 65.805 166.305 65.975 166.475 ;
        RECT 66.265 166.305 66.435 166.475 ;
        RECT 67.645 166.645 67.815 166.815 ;
        RECT 67.185 166.305 67.355 166.475 ;
        RECT 72.705 167.665 72.875 167.835 ;
        RECT 76.385 167.665 76.555 167.835 ;
        RECT 70.405 166.645 70.575 166.815 ;
        RECT 70.865 166.305 71.035 166.475 ;
        RECT 71.325 166.645 71.495 166.815 ;
        RECT 72.245 166.645 72.415 166.815 ;
        RECT 72.705 166.645 72.875 166.815 ;
        RECT 73.625 166.645 73.795 166.815 ;
        RECT 76.845 166.645 77.015 166.815 ;
        RECT 69.485 165.965 69.655 166.135 ;
        RECT 78.225 166.985 78.395 167.155 ;
        RECT 81.905 167.665 82.075 167.835 ;
        RECT 77.765 166.645 77.935 166.815 ;
        RECT 78.685 166.645 78.855 166.815 ;
        RECT 80.985 166.645 81.155 166.815 ;
        RECT 84.665 166.645 84.835 166.815 ;
        RECT 85.125 166.645 85.295 166.815 ;
        RECT 85.585 166.645 85.755 166.815 ;
        RECT 83.285 165.965 83.455 166.135 ;
        RECT 86.505 166.645 86.675 166.815 ;
        RECT 18.425 165.455 18.595 165.625 ;
        RECT 18.885 165.455 19.055 165.625 ;
        RECT 19.345 165.455 19.515 165.625 ;
        RECT 19.805 165.455 19.975 165.625 ;
        RECT 20.265 165.455 20.435 165.625 ;
        RECT 20.725 165.455 20.895 165.625 ;
        RECT 21.185 165.455 21.355 165.625 ;
        RECT 21.645 165.455 21.815 165.625 ;
        RECT 22.105 165.455 22.275 165.625 ;
        RECT 22.565 165.455 22.735 165.625 ;
        RECT 23.025 165.455 23.195 165.625 ;
        RECT 23.485 165.455 23.655 165.625 ;
        RECT 23.945 165.455 24.115 165.625 ;
        RECT 24.405 165.455 24.575 165.625 ;
        RECT 24.865 165.455 25.035 165.625 ;
        RECT 25.325 165.455 25.495 165.625 ;
        RECT 25.785 165.455 25.955 165.625 ;
        RECT 26.245 165.455 26.415 165.625 ;
        RECT 26.705 165.455 26.875 165.625 ;
        RECT 27.165 165.455 27.335 165.625 ;
        RECT 27.625 165.455 27.795 165.625 ;
        RECT 28.085 165.455 28.255 165.625 ;
        RECT 28.545 165.455 28.715 165.625 ;
        RECT 29.005 165.455 29.175 165.625 ;
        RECT 29.465 165.455 29.635 165.625 ;
        RECT 29.925 165.455 30.095 165.625 ;
        RECT 30.385 165.455 30.555 165.625 ;
        RECT 30.845 165.455 31.015 165.625 ;
        RECT 31.305 165.455 31.475 165.625 ;
        RECT 31.765 165.455 31.935 165.625 ;
        RECT 32.225 165.455 32.395 165.625 ;
        RECT 32.685 165.455 32.855 165.625 ;
        RECT 33.145 165.455 33.315 165.625 ;
        RECT 33.605 165.455 33.775 165.625 ;
        RECT 34.065 165.455 34.235 165.625 ;
        RECT 34.525 165.455 34.695 165.625 ;
        RECT 34.985 165.455 35.155 165.625 ;
        RECT 35.445 165.455 35.615 165.625 ;
        RECT 35.905 165.455 36.075 165.625 ;
        RECT 36.365 165.455 36.535 165.625 ;
        RECT 36.825 165.455 36.995 165.625 ;
        RECT 37.285 165.455 37.455 165.625 ;
        RECT 37.745 165.455 37.915 165.625 ;
        RECT 38.205 165.455 38.375 165.625 ;
        RECT 38.665 165.455 38.835 165.625 ;
        RECT 39.125 165.455 39.295 165.625 ;
        RECT 39.585 165.455 39.755 165.625 ;
        RECT 40.045 165.455 40.215 165.625 ;
        RECT 40.505 165.455 40.675 165.625 ;
        RECT 40.965 165.455 41.135 165.625 ;
        RECT 41.425 165.455 41.595 165.625 ;
        RECT 41.885 165.455 42.055 165.625 ;
        RECT 42.345 165.455 42.515 165.625 ;
        RECT 42.805 165.455 42.975 165.625 ;
        RECT 43.265 165.455 43.435 165.625 ;
        RECT 43.725 165.455 43.895 165.625 ;
        RECT 44.185 165.455 44.355 165.625 ;
        RECT 44.645 165.455 44.815 165.625 ;
        RECT 45.105 165.455 45.275 165.625 ;
        RECT 45.565 165.455 45.735 165.625 ;
        RECT 46.025 165.455 46.195 165.625 ;
        RECT 46.485 165.455 46.655 165.625 ;
        RECT 46.945 165.455 47.115 165.625 ;
        RECT 47.405 165.455 47.575 165.625 ;
        RECT 47.865 165.455 48.035 165.625 ;
        RECT 48.325 165.455 48.495 165.625 ;
        RECT 48.785 165.455 48.955 165.625 ;
        RECT 49.245 165.455 49.415 165.625 ;
        RECT 49.705 165.455 49.875 165.625 ;
        RECT 50.165 165.455 50.335 165.625 ;
        RECT 50.625 165.455 50.795 165.625 ;
        RECT 51.085 165.455 51.255 165.625 ;
        RECT 51.545 165.455 51.715 165.625 ;
        RECT 52.005 165.455 52.175 165.625 ;
        RECT 52.465 165.455 52.635 165.625 ;
        RECT 52.925 165.455 53.095 165.625 ;
        RECT 53.385 165.455 53.555 165.625 ;
        RECT 53.845 165.455 54.015 165.625 ;
        RECT 54.305 165.455 54.475 165.625 ;
        RECT 54.765 165.455 54.935 165.625 ;
        RECT 55.225 165.455 55.395 165.625 ;
        RECT 55.685 165.455 55.855 165.625 ;
        RECT 56.145 165.455 56.315 165.625 ;
        RECT 56.605 165.455 56.775 165.625 ;
        RECT 57.065 165.455 57.235 165.625 ;
        RECT 57.525 165.455 57.695 165.625 ;
        RECT 57.985 165.455 58.155 165.625 ;
        RECT 58.445 165.455 58.615 165.625 ;
        RECT 58.905 165.455 59.075 165.625 ;
        RECT 59.365 165.455 59.535 165.625 ;
        RECT 59.825 165.455 59.995 165.625 ;
        RECT 60.285 165.455 60.455 165.625 ;
        RECT 60.745 165.455 60.915 165.625 ;
        RECT 61.205 165.455 61.375 165.625 ;
        RECT 61.665 165.455 61.835 165.625 ;
        RECT 62.125 165.455 62.295 165.625 ;
        RECT 62.585 165.455 62.755 165.625 ;
        RECT 63.045 165.455 63.215 165.625 ;
        RECT 63.505 165.455 63.675 165.625 ;
        RECT 63.965 165.455 64.135 165.625 ;
        RECT 64.425 165.455 64.595 165.625 ;
        RECT 64.885 165.455 65.055 165.625 ;
        RECT 65.345 165.455 65.515 165.625 ;
        RECT 65.805 165.455 65.975 165.625 ;
        RECT 66.265 165.455 66.435 165.625 ;
        RECT 66.725 165.455 66.895 165.625 ;
        RECT 67.185 165.455 67.355 165.625 ;
        RECT 67.645 165.455 67.815 165.625 ;
        RECT 68.105 165.455 68.275 165.625 ;
        RECT 68.565 165.455 68.735 165.625 ;
        RECT 69.025 165.455 69.195 165.625 ;
        RECT 69.485 165.455 69.655 165.625 ;
        RECT 69.945 165.455 70.115 165.625 ;
        RECT 70.405 165.455 70.575 165.625 ;
        RECT 70.865 165.455 71.035 165.625 ;
        RECT 71.325 165.455 71.495 165.625 ;
        RECT 71.785 165.455 71.955 165.625 ;
        RECT 72.245 165.455 72.415 165.625 ;
        RECT 72.705 165.455 72.875 165.625 ;
        RECT 73.165 165.455 73.335 165.625 ;
        RECT 73.625 165.455 73.795 165.625 ;
        RECT 74.085 165.455 74.255 165.625 ;
        RECT 74.545 165.455 74.715 165.625 ;
        RECT 75.005 165.455 75.175 165.625 ;
        RECT 75.465 165.455 75.635 165.625 ;
        RECT 75.925 165.455 76.095 165.625 ;
        RECT 76.385 165.455 76.555 165.625 ;
        RECT 76.845 165.455 77.015 165.625 ;
        RECT 77.305 165.455 77.475 165.625 ;
        RECT 77.765 165.455 77.935 165.625 ;
        RECT 78.225 165.455 78.395 165.625 ;
        RECT 78.685 165.455 78.855 165.625 ;
        RECT 79.145 165.455 79.315 165.625 ;
        RECT 79.605 165.455 79.775 165.625 ;
        RECT 80.065 165.455 80.235 165.625 ;
        RECT 80.525 165.455 80.695 165.625 ;
        RECT 80.985 165.455 81.155 165.625 ;
        RECT 81.445 165.455 81.615 165.625 ;
        RECT 81.905 165.455 82.075 165.625 ;
        RECT 82.365 165.455 82.535 165.625 ;
        RECT 82.825 165.455 82.995 165.625 ;
        RECT 83.285 165.455 83.455 165.625 ;
        RECT 83.745 165.455 83.915 165.625 ;
        RECT 84.205 165.455 84.375 165.625 ;
        RECT 84.665 165.455 84.835 165.625 ;
        RECT 85.125 165.455 85.295 165.625 ;
        RECT 85.585 165.455 85.755 165.625 ;
        RECT 86.045 165.455 86.215 165.625 ;
        RECT 86.505 165.455 86.675 165.625 ;
        RECT 86.965 165.455 87.135 165.625 ;
        RECT 87.425 165.455 87.595 165.625 ;
        RECT 87.885 165.455 88.055 165.625 ;
        RECT 88.345 165.455 88.515 165.625 ;
        RECT 88.805 165.455 88.975 165.625 ;
        RECT 89.265 165.455 89.435 165.625 ;
        RECT 89.725 165.455 89.895 165.625 ;
        RECT 90.185 165.455 90.355 165.625 ;
        RECT 90.645 165.455 90.815 165.625 ;
        RECT 91.105 165.455 91.275 165.625 ;
        RECT 91.565 165.455 91.735 165.625 ;
        RECT 92.025 165.455 92.195 165.625 ;
        RECT 30.370 164.265 30.540 164.435 ;
        RECT 29.465 163.245 29.635 163.415 ;
        RECT 32.685 163.925 32.855 164.095 ;
        RECT 35.020 164.265 35.190 164.435 ;
        RECT 32.225 163.245 32.395 163.415 ;
        RECT 35.445 163.925 35.615 164.095 ;
        RECT 36.365 164.265 36.535 164.435 ;
        RECT 37.285 164.265 37.455 164.435 ;
        RECT 42.345 164.945 42.515 165.115 ;
        RECT 33.145 163.245 33.315 163.415 ;
        RECT 36.825 163.245 36.995 163.415 ;
        RECT 41.885 164.265 42.055 164.435 ;
        RECT 42.805 164.265 42.975 164.435 ;
        RECT 46.485 164.265 46.655 164.435 ;
        RECT 47.405 164.265 47.575 164.435 ;
        RECT 46.945 163.925 47.115 164.095 ;
        RECT 48.785 164.265 48.955 164.435 ;
        RECT 47.865 163.585 48.035 163.755 ;
        RECT 49.705 163.925 49.875 164.095 ;
        RECT 50.165 163.925 50.335 164.095 ;
        RECT 49.245 163.585 49.415 163.755 ;
        RECT 51.085 164.265 51.255 164.435 ;
        RECT 75.925 164.945 76.095 165.115 ;
        RECT 78.225 164.945 78.395 165.115 ;
        RECT 75.465 164.265 75.635 164.435 ;
        RECT 76.845 164.265 77.015 164.435 ;
        RECT 76.845 163.585 77.015 163.755 ;
        RECT 78.985 164.605 79.155 164.775 ;
        RECT 80.065 164.605 80.235 164.775 ;
        RECT 79.145 163.245 79.315 163.415 ;
        RECT 82.365 164.265 82.535 164.435 ;
        RECT 82.830 163.585 83.000 163.755 ;
        RECT 83.290 164.605 83.460 164.775 ;
        RECT 83.745 164.265 83.915 164.435 ;
        RECT 84.690 164.605 84.860 164.775 ;
        RECT 86.530 164.605 86.700 164.775 ;
        RECT 85.150 163.585 85.320 163.755 ;
        RECT 86.530 163.585 86.700 163.755 ;
        RECT 90.645 164.265 90.815 164.435 ;
        RECT 18.425 162.735 18.595 162.905 ;
        RECT 18.885 162.735 19.055 162.905 ;
        RECT 19.345 162.735 19.515 162.905 ;
        RECT 19.805 162.735 19.975 162.905 ;
        RECT 20.265 162.735 20.435 162.905 ;
        RECT 20.725 162.735 20.895 162.905 ;
        RECT 21.185 162.735 21.355 162.905 ;
        RECT 21.645 162.735 21.815 162.905 ;
        RECT 22.105 162.735 22.275 162.905 ;
        RECT 22.565 162.735 22.735 162.905 ;
        RECT 23.025 162.735 23.195 162.905 ;
        RECT 23.485 162.735 23.655 162.905 ;
        RECT 23.945 162.735 24.115 162.905 ;
        RECT 24.405 162.735 24.575 162.905 ;
        RECT 24.865 162.735 25.035 162.905 ;
        RECT 25.325 162.735 25.495 162.905 ;
        RECT 25.785 162.735 25.955 162.905 ;
        RECT 26.245 162.735 26.415 162.905 ;
        RECT 26.705 162.735 26.875 162.905 ;
        RECT 27.165 162.735 27.335 162.905 ;
        RECT 27.625 162.735 27.795 162.905 ;
        RECT 28.085 162.735 28.255 162.905 ;
        RECT 28.545 162.735 28.715 162.905 ;
        RECT 29.005 162.735 29.175 162.905 ;
        RECT 29.465 162.735 29.635 162.905 ;
        RECT 29.925 162.735 30.095 162.905 ;
        RECT 30.385 162.735 30.555 162.905 ;
        RECT 30.845 162.735 31.015 162.905 ;
        RECT 31.305 162.735 31.475 162.905 ;
        RECT 31.765 162.735 31.935 162.905 ;
        RECT 32.225 162.735 32.395 162.905 ;
        RECT 32.685 162.735 32.855 162.905 ;
        RECT 33.145 162.735 33.315 162.905 ;
        RECT 33.605 162.735 33.775 162.905 ;
        RECT 34.065 162.735 34.235 162.905 ;
        RECT 34.525 162.735 34.695 162.905 ;
        RECT 34.985 162.735 35.155 162.905 ;
        RECT 35.445 162.735 35.615 162.905 ;
        RECT 35.905 162.735 36.075 162.905 ;
        RECT 36.365 162.735 36.535 162.905 ;
        RECT 36.825 162.735 36.995 162.905 ;
        RECT 37.285 162.735 37.455 162.905 ;
        RECT 37.745 162.735 37.915 162.905 ;
        RECT 38.205 162.735 38.375 162.905 ;
        RECT 38.665 162.735 38.835 162.905 ;
        RECT 39.125 162.735 39.295 162.905 ;
        RECT 39.585 162.735 39.755 162.905 ;
        RECT 40.045 162.735 40.215 162.905 ;
        RECT 40.505 162.735 40.675 162.905 ;
        RECT 40.965 162.735 41.135 162.905 ;
        RECT 41.425 162.735 41.595 162.905 ;
        RECT 41.885 162.735 42.055 162.905 ;
        RECT 42.345 162.735 42.515 162.905 ;
        RECT 42.805 162.735 42.975 162.905 ;
        RECT 43.265 162.735 43.435 162.905 ;
        RECT 43.725 162.735 43.895 162.905 ;
        RECT 44.185 162.735 44.355 162.905 ;
        RECT 44.645 162.735 44.815 162.905 ;
        RECT 45.105 162.735 45.275 162.905 ;
        RECT 45.565 162.735 45.735 162.905 ;
        RECT 46.025 162.735 46.195 162.905 ;
        RECT 46.485 162.735 46.655 162.905 ;
        RECT 46.945 162.735 47.115 162.905 ;
        RECT 47.405 162.735 47.575 162.905 ;
        RECT 47.865 162.735 48.035 162.905 ;
        RECT 48.325 162.735 48.495 162.905 ;
        RECT 48.785 162.735 48.955 162.905 ;
        RECT 49.245 162.735 49.415 162.905 ;
        RECT 49.705 162.735 49.875 162.905 ;
        RECT 50.165 162.735 50.335 162.905 ;
        RECT 50.625 162.735 50.795 162.905 ;
        RECT 51.085 162.735 51.255 162.905 ;
        RECT 51.545 162.735 51.715 162.905 ;
        RECT 52.005 162.735 52.175 162.905 ;
        RECT 52.465 162.735 52.635 162.905 ;
        RECT 52.925 162.735 53.095 162.905 ;
        RECT 53.385 162.735 53.555 162.905 ;
        RECT 53.845 162.735 54.015 162.905 ;
        RECT 54.305 162.735 54.475 162.905 ;
        RECT 54.765 162.735 54.935 162.905 ;
        RECT 55.225 162.735 55.395 162.905 ;
        RECT 55.685 162.735 55.855 162.905 ;
        RECT 56.145 162.735 56.315 162.905 ;
        RECT 56.605 162.735 56.775 162.905 ;
        RECT 57.065 162.735 57.235 162.905 ;
        RECT 57.525 162.735 57.695 162.905 ;
        RECT 57.985 162.735 58.155 162.905 ;
        RECT 58.445 162.735 58.615 162.905 ;
        RECT 58.905 162.735 59.075 162.905 ;
        RECT 59.365 162.735 59.535 162.905 ;
        RECT 59.825 162.735 59.995 162.905 ;
        RECT 60.285 162.735 60.455 162.905 ;
        RECT 60.745 162.735 60.915 162.905 ;
        RECT 61.205 162.735 61.375 162.905 ;
        RECT 61.665 162.735 61.835 162.905 ;
        RECT 62.125 162.735 62.295 162.905 ;
        RECT 62.585 162.735 62.755 162.905 ;
        RECT 63.045 162.735 63.215 162.905 ;
        RECT 63.505 162.735 63.675 162.905 ;
        RECT 63.965 162.735 64.135 162.905 ;
        RECT 64.425 162.735 64.595 162.905 ;
        RECT 64.885 162.735 65.055 162.905 ;
        RECT 65.345 162.735 65.515 162.905 ;
        RECT 65.805 162.735 65.975 162.905 ;
        RECT 66.265 162.735 66.435 162.905 ;
        RECT 66.725 162.735 66.895 162.905 ;
        RECT 67.185 162.735 67.355 162.905 ;
        RECT 67.645 162.735 67.815 162.905 ;
        RECT 68.105 162.735 68.275 162.905 ;
        RECT 68.565 162.735 68.735 162.905 ;
        RECT 69.025 162.735 69.195 162.905 ;
        RECT 69.485 162.735 69.655 162.905 ;
        RECT 69.945 162.735 70.115 162.905 ;
        RECT 70.405 162.735 70.575 162.905 ;
        RECT 70.865 162.735 71.035 162.905 ;
        RECT 71.325 162.735 71.495 162.905 ;
        RECT 71.785 162.735 71.955 162.905 ;
        RECT 72.245 162.735 72.415 162.905 ;
        RECT 72.705 162.735 72.875 162.905 ;
        RECT 73.165 162.735 73.335 162.905 ;
        RECT 73.625 162.735 73.795 162.905 ;
        RECT 74.085 162.735 74.255 162.905 ;
        RECT 74.545 162.735 74.715 162.905 ;
        RECT 75.005 162.735 75.175 162.905 ;
        RECT 75.465 162.735 75.635 162.905 ;
        RECT 75.925 162.735 76.095 162.905 ;
        RECT 76.385 162.735 76.555 162.905 ;
        RECT 76.845 162.735 77.015 162.905 ;
        RECT 77.305 162.735 77.475 162.905 ;
        RECT 77.765 162.735 77.935 162.905 ;
        RECT 78.225 162.735 78.395 162.905 ;
        RECT 78.685 162.735 78.855 162.905 ;
        RECT 79.145 162.735 79.315 162.905 ;
        RECT 79.605 162.735 79.775 162.905 ;
        RECT 80.065 162.735 80.235 162.905 ;
        RECT 80.525 162.735 80.695 162.905 ;
        RECT 80.985 162.735 81.155 162.905 ;
        RECT 81.445 162.735 81.615 162.905 ;
        RECT 81.905 162.735 82.075 162.905 ;
        RECT 82.365 162.735 82.535 162.905 ;
        RECT 82.825 162.735 82.995 162.905 ;
        RECT 83.285 162.735 83.455 162.905 ;
        RECT 83.745 162.735 83.915 162.905 ;
        RECT 84.205 162.735 84.375 162.905 ;
        RECT 84.665 162.735 84.835 162.905 ;
        RECT 85.125 162.735 85.295 162.905 ;
        RECT 85.585 162.735 85.755 162.905 ;
        RECT 86.045 162.735 86.215 162.905 ;
        RECT 86.505 162.735 86.675 162.905 ;
        RECT 86.965 162.735 87.135 162.905 ;
        RECT 87.425 162.735 87.595 162.905 ;
        RECT 87.885 162.735 88.055 162.905 ;
        RECT 88.345 162.735 88.515 162.905 ;
        RECT 88.805 162.735 88.975 162.905 ;
        RECT 89.265 162.735 89.435 162.905 ;
        RECT 89.725 162.735 89.895 162.905 ;
        RECT 90.185 162.735 90.355 162.905 ;
        RECT 90.645 162.735 90.815 162.905 ;
        RECT 91.105 162.735 91.275 162.905 ;
        RECT 91.565 162.735 91.735 162.905 ;
        RECT 92.025 162.735 92.195 162.905 ;
        RECT 23.050 161.885 23.220 162.055 ;
        RECT 22.565 161.545 22.735 161.715 ;
        RECT 23.445 161.545 23.615 161.715 ;
        RECT 23.900 160.865 24.070 161.035 ;
        RECT 25.150 161.885 25.320 162.055 ;
        RECT 24.635 161.545 24.805 161.715 ;
        RECT 26.720 161.885 26.890 162.055 ;
        RECT 27.155 161.545 27.325 161.715 ;
        RECT 29.925 161.205 30.095 161.375 ;
        RECT 30.845 161.205 31.015 161.375 ;
        RECT 29.465 160.525 29.635 160.695 ;
        RECT 30.385 160.865 30.555 161.035 ;
        RECT 37.285 162.225 37.455 162.395 ;
        RECT 36.365 161.545 36.535 161.715 ;
        RECT 38.665 161.545 38.835 161.715 ;
        RECT 37.745 161.205 37.915 161.375 ;
        RECT 38.205 161.205 38.375 161.375 ;
        RECT 34.985 160.525 35.155 160.695 ;
        RECT 39.125 161.205 39.295 161.375 ;
        RECT 45.105 161.205 45.275 161.375 ;
        RECT 45.565 161.205 45.735 161.375 ;
        RECT 46.025 161.205 46.195 161.375 ;
        RECT 46.485 161.205 46.655 161.375 ;
        RECT 47.865 161.885 48.035 162.055 ;
        RECT 47.405 161.205 47.575 161.375 ;
        RECT 44.185 160.525 44.355 160.695 ;
        RECT 50.625 162.225 50.795 162.395 ;
        RECT 48.785 160.525 48.955 160.695 ;
        RECT 49.245 160.865 49.415 161.035 ;
        RECT 49.705 160.525 49.875 160.695 ;
        RECT 52.005 161.205 52.175 161.375 ;
        RECT 52.465 161.205 52.635 161.375 ;
        RECT 54.765 161.545 54.935 161.715 ;
        RECT 54.305 161.205 54.475 161.375 ;
        RECT 56.145 161.885 56.315 162.055 ;
        RECT 57.985 161.885 58.155 162.055 ;
        RECT 57.525 161.205 57.695 161.375 ;
        RECT 60.120 161.205 60.290 161.375 ;
        RECT 59.825 160.525 59.995 160.695 ;
        RECT 60.745 160.525 60.915 160.695 ;
        RECT 63.965 162.225 64.135 162.395 ;
        RECT 64.885 161.885 65.055 162.055 ;
        RECT 63.045 161.205 63.215 161.375 ;
        RECT 64.425 161.205 64.595 161.375 ;
        RECT 62.125 160.525 62.295 160.695 ;
        RECT 64.885 160.865 65.055 161.035 ;
        RECT 65.805 161.205 65.975 161.375 ;
        RECT 66.265 161.205 66.435 161.375 ;
        RECT 70.405 162.225 70.575 162.395 ;
        RECT 69.945 161.205 70.115 161.375 ;
        RECT 71.325 161.545 71.495 161.715 ;
        RECT 71.785 161.205 71.955 161.375 ;
        RECT 72.705 161.205 72.875 161.375 ;
        RECT 71.325 160.525 71.495 160.695 ;
        RECT 72.245 160.525 72.415 160.695 ;
        RECT 79.145 161.205 79.315 161.375 ;
        RECT 80.525 161.205 80.695 161.375 ;
        RECT 81.445 161.205 81.615 161.375 ;
        RECT 83.285 161.205 83.455 161.375 ;
        RECT 86.965 162.225 87.135 162.395 ;
        RECT 86.505 161.205 86.675 161.375 ;
        RECT 89.725 161.885 89.895 162.055 ;
        RECT 87.885 160.525 88.055 160.695 ;
        RECT 88.345 160.525 88.515 160.695 ;
        RECT 88.805 161.205 88.975 161.375 ;
        RECT 18.425 160.015 18.595 160.185 ;
        RECT 18.885 160.015 19.055 160.185 ;
        RECT 19.345 160.015 19.515 160.185 ;
        RECT 19.805 160.015 19.975 160.185 ;
        RECT 20.265 160.015 20.435 160.185 ;
        RECT 20.725 160.015 20.895 160.185 ;
        RECT 21.185 160.015 21.355 160.185 ;
        RECT 21.645 160.015 21.815 160.185 ;
        RECT 22.105 160.015 22.275 160.185 ;
        RECT 22.565 160.015 22.735 160.185 ;
        RECT 23.025 160.015 23.195 160.185 ;
        RECT 23.485 160.015 23.655 160.185 ;
        RECT 23.945 160.015 24.115 160.185 ;
        RECT 24.405 160.015 24.575 160.185 ;
        RECT 24.865 160.015 25.035 160.185 ;
        RECT 25.325 160.015 25.495 160.185 ;
        RECT 25.785 160.015 25.955 160.185 ;
        RECT 26.245 160.015 26.415 160.185 ;
        RECT 26.705 160.015 26.875 160.185 ;
        RECT 27.165 160.015 27.335 160.185 ;
        RECT 27.625 160.015 27.795 160.185 ;
        RECT 28.085 160.015 28.255 160.185 ;
        RECT 28.545 160.015 28.715 160.185 ;
        RECT 29.005 160.015 29.175 160.185 ;
        RECT 29.465 160.015 29.635 160.185 ;
        RECT 29.925 160.015 30.095 160.185 ;
        RECT 30.385 160.015 30.555 160.185 ;
        RECT 30.845 160.015 31.015 160.185 ;
        RECT 31.305 160.015 31.475 160.185 ;
        RECT 31.765 160.015 31.935 160.185 ;
        RECT 32.225 160.015 32.395 160.185 ;
        RECT 32.685 160.015 32.855 160.185 ;
        RECT 33.145 160.015 33.315 160.185 ;
        RECT 33.605 160.015 33.775 160.185 ;
        RECT 34.065 160.015 34.235 160.185 ;
        RECT 34.525 160.015 34.695 160.185 ;
        RECT 34.985 160.015 35.155 160.185 ;
        RECT 35.445 160.015 35.615 160.185 ;
        RECT 35.905 160.015 36.075 160.185 ;
        RECT 36.365 160.015 36.535 160.185 ;
        RECT 36.825 160.015 36.995 160.185 ;
        RECT 37.285 160.015 37.455 160.185 ;
        RECT 37.745 160.015 37.915 160.185 ;
        RECT 38.205 160.015 38.375 160.185 ;
        RECT 38.665 160.015 38.835 160.185 ;
        RECT 39.125 160.015 39.295 160.185 ;
        RECT 39.585 160.015 39.755 160.185 ;
        RECT 40.045 160.015 40.215 160.185 ;
        RECT 40.505 160.015 40.675 160.185 ;
        RECT 40.965 160.015 41.135 160.185 ;
        RECT 41.425 160.015 41.595 160.185 ;
        RECT 41.885 160.015 42.055 160.185 ;
        RECT 42.345 160.015 42.515 160.185 ;
        RECT 42.805 160.015 42.975 160.185 ;
        RECT 43.265 160.015 43.435 160.185 ;
        RECT 43.725 160.015 43.895 160.185 ;
        RECT 44.185 160.015 44.355 160.185 ;
        RECT 44.645 160.015 44.815 160.185 ;
        RECT 45.105 160.015 45.275 160.185 ;
        RECT 45.565 160.015 45.735 160.185 ;
        RECT 46.025 160.015 46.195 160.185 ;
        RECT 46.485 160.015 46.655 160.185 ;
        RECT 46.945 160.015 47.115 160.185 ;
        RECT 47.405 160.015 47.575 160.185 ;
        RECT 47.865 160.015 48.035 160.185 ;
        RECT 48.325 160.015 48.495 160.185 ;
        RECT 48.785 160.015 48.955 160.185 ;
        RECT 49.245 160.015 49.415 160.185 ;
        RECT 49.705 160.015 49.875 160.185 ;
        RECT 50.165 160.015 50.335 160.185 ;
        RECT 50.625 160.015 50.795 160.185 ;
        RECT 51.085 160.015 51.255 160.185 ;
        RECT 51.545 160.015 51.715 160.185 ;
        RECT 52.005 160.015 52.175 160.185 ;
        RECT 52.465 160.015 52.635 160.185 ;
        RECT 52.925 160.015 53.095 160.185 ;
        RECT 53.385 160.015 53.555 160.185 ;
        RECT 53.845 160.015 54.015 160.185 ;
        RECT 54.305 160.015 54.475 160.185 ;
        RECT 54.765 160.015 54.935 160.185 ;
        RECT 55.225 160.015 55.395 160.185 ;
        RECT 55.685 160.015 55.855 160.185 ;
        RECT 56.145 160.015 56.315 160.185 ;
        RECT 56.605 160.015 56.775 160.185 ;
        RECT 57.065 160.015 57.235 160.185 ;
        RECT 57.525 160.015 57.695 160.185 ;
        RECT 57.985 160.015 58.155 160.185 ;
        RECT 58.445 160.015 58.615 160.185 ;
        RECT 58.905 160.015 59.075 160.185 ;
        RECT 59.365 160.015 59.535 160.185 ;
        RECT 59.825 160.015 59.995 160.185 ;
        RECT 60.285 160.015 60.455 160.185 ;
        RECT 60.745 160.015 60.915 160.185 ;
        RECT 61.205 160.015 61.375 160.185 ;
        RECT 61.665 160.015 61.835 160.185 ;
        RECT 62.125 160.015 62.295 160.185 ;
        RECT 62.585 160.015 62.755 160.185 ;
        RECT 63.045 160.015 63.215 160.185 ;
        RECT 63.505 160.015 63.675 160.185 ;
        RECT 63.965 160.015 64.135 160.185 ;
        RECT 64.425 160.015 64.595 160.185 ;
        RECT 64.885 160.015 65.055 160.185 ;
        RECT 65.345 160.015 65.515 160.185 ;
        RECT 65.805 160.015 65.975 160.185 ;
        RECT 66.265 160.015 66.435 160.185 ;
        RECT 66.725 160.015 66.895 160.185 ;
        RECT 67.185 160.015 67.355 160.185 ;
        RECT 67.645 160.015 67.815 160.185 ;
        RECT 68.105 160.015 68.275 160.185 ;
        RECT 68.565 160.015 68.735 160.185 ;
        RECT 69.025 160.015 69.195 160.185 ;
        RECT 69.485 160.015 69.655 160.185 ;
        RECT 69.945 160.015 70.115 160.185 ;
        RECT 70.405 160.015 70.575 160.185 ;
        RECT 70.865 160.015 71.035 160.185 ;
        RECT 71.325 160.015 71.495 160.185 ;
        RECT 71.785 160.015 71.955 160.185 ;
        RECT 72.245 160.015 72.415 160.185 ;
        RECT 72.705 160.015 72.875 160.185 ;
        RECT 73.165 160.015 73.335 160.185 ;
        RECT 73.625 160.015 73.795 160.185 ;
        RECT 74.085 160.015 74.255 160.185 ;
        RECT 74.545 160.015 74.715 160.185 ;
        RECT 75.005 160.015 75.175 160.185 ;
        RECT 75.465 160.015 75.635 160.185 ;
        RECT 75.925 160.015 76.095 160.185 ;
        RECT 76.385 160.015 76.555 160.185 ;
        RECT 76.845 160.015 77.015 160.185 ;
        RECT 77.305 160.015 77.475 160.185 ;
        RECT 77.765 160.015 77.935 160.185 ;
        RECT 78.225 160.015 78.395 160.185 ;
        RECT 78.685 160.015 78.855 160.185 ;
        RECT 79.145 160.015 79.315 160.185 ;
        RECT 79.605 160.015 79.775 160.185 ;
        RECT 80.065 160.015 80.235 160.185 ;
        RECT 80.525 160.015 80.695 160.185 ;
        RECT 80.985 160.015 81.155 160.185 ;
        RECT 81.445 160.015 81.615 160.185 ;
        RECT 81.905 160.015 82.075 160.185 ;
        RECT 82.365 160.015 82.535 160.185 ;
        RECT 82.825 160.015 82.995 160.185 ;
        RECT 83.285 160.015 83.455 160.185 ;
        RECT 83.745 160.015 83.915 160.185 ;
        RECT 84.205 160.015 84.375 160.185 ;
        RECT 84.665 160.015 84.835 160.185 ;
        RECT 85.125 160.015 85.295 160.185 ;
        RECT 85.585 160.015 85.755 160.185 ;
        RECT 86.045 160.015 86.215 160.185 ;
        RECT 86.505 160.015 86.675 160.185 ;
        RECT 86.965 160.015 87.135 160.185 ;
        RECT 87.425 160.015 87.595 160.185 ;
        RECT 87.885 160.015 88.055 160.185 ;
        RECT 88.345 160.015 88.515 160.185 ;
        RECT 88.805 160.015 88.975 160.185 ;
        RECT 89.265 160.015 89.435 160.185 ;
        RECT 89.725 160.015 89.895 160.185 ;
        RECT 90.185 160.015 90.355 160.185 ;
        RECT 90.645 160.015 90.815 160.185 ;
        RECT 91.105 160.015 91.275 160.185 ;
        RECT 91.565 160.015 91.735 160.185 ;
        RECT 92.025 160.015 92.195 160.185 ;
        RECT 34.065 159.165 34.235 159.335 ;
        RECT 34.985 158.825 35.155 158.995 ;
        RECT 35.445 158.825 35.615 158.995 ;
        RECT 35.905 158.825 36.075 158.995 ;
        RECT 36.825 158.825 36.995 158.995 ;
        RECT 38.205 158.825 38.375 158.995 ;
        RECT 34.065 157.805 34.235 157.975 ;
        RECT 36.365 158.485 36.535 158.655 ;
        RECT 40.965 158.825 41.135 158.995 ;
        RECT 41.885 158.825 42.055 158.995 ;
        RECT 42.805 158.825 42.975 158.995 ;
        RECT 45.565 158.825 45.735 158.995 ;
        RECT 42.805 157.805 42.975 157.975 ;
        RECT 47.405 159.505 47.575 159.675 ;
        RECT 48.220 159.505 48.390 159.675 ;
        RECT 46.485 158.825 46.655 158.995 ;
        RECT 46.945 158.825 47.115 158.995 ;
        RECT 45.565 158.145 45.735 158.315 ;
        RECT 49.245 159.165 49.415 159.335 ;
        RECT 49.705 158.825 49.875 158.995 ;
        RECT 48.325 157.805 48.495 157.975 ;
        RECT 52.925 159.505 53.095 159.675 ;
        RECT 53.385 158.825 53.555 158.995 ;
        RECT 54.765 159.165 54.935 159.335 ;
        RECT 54.305 158.825 54.475 158.995 ;
        RECT 61.205 159.505 61.375 159.675 ;
        RECT 54.305 157.805 54.475 157.975 ;
        RECT 65.805 159.505 65.975 159.675 ;
        RECT 71.785 158.825 71.955 158.995 ;
        RECT 72.245 158.825 72.415 158.995 ;
        RECT 73.165 159.165 73.335 159.335 ;
        RECT 73.165 157.805 73.335 157.975 ;
        RECT 76.385 159.505 76.555 159.675 ;
        RECT 75.925 158.825 76.095 158.995 ;
        RECT 79.605 158.485 79.775 158.655 ;
        RECT 80.070 158.145 80.240 158.315 ;
        RECT 80.530 159.165 80.700 159.335 ;
        RECT 80.985 158.825 81.155 158.995 ;
        RECT 81.930 159.165 82.100 159.335 ;
        RECT 83.770 159.165 83.940 159.335 ;
        RECT 82.390 158.145 82.560 158.315 ;
        RECT 83.770 158.145 83.940 158.315 ;
        RECT 87.425 157.805 87.595 157.975 ;
        RECT 18.425 157.295 18.595 157.465 ;
        RECT 18.885 157.295 19.055 157.465 ;
        RECT 19.345 157.295 19.515 157.465 ;
        RECT 19.805 157.295 19.975 157.465 ;
        RECT 20.265 157.295 20.435 157.465 ;
        RECT 20.725 157.295 20.895 157.465 ;
        RECT 21.185 157.295 21.355 157.465 ;
        RECT 21.645 157.295 21.815 157.465 ;
        RECT 22.105 157.295 22.275 157.465 ;
        RECT 22.565 157.295 22.735 157.465 ;
        RECT 23.025 157.295 23.195 157.465 ;
        RECT 23.485 157.295 23.655 157.465 ;
        RECT 23.945 157.295 24.115 157.465 ;
        RECT 24.405 157.295 24.575 157.465 ;
        RECT 24.865 157.295 25.035 157.465 ;
        RECT 25.325 157.295 25.495 157.465 ;
        RECT 25.785 157.295 25.955 157.465 ;
        RECT 26.245 157.295 26.415 157.465 ;
        RECT 26.705 157.295 26.875 157.465 ;
        RECT 27.165 157.295 27.335 157.465 ;
        RECT 27.625 157.295 27.795 157.465 ;
        RECT 28.085 157.295 28.255 157.465 ;
        RECT 28.545 157.295 28.715 157.465 ;
        RECT 29.005 157.295 29.175 157.465 ;
        RECT 29.465 157.295 29.635 157.465 ;
        RECT 29.925 157.295 30.095 157.465 ;
        RECT 30.385 157.295 30.555 157.465 ;
        RECT 30.845 157.295 31.015 157.465 ;
        RECT 31.305 157.295 31.475 157.465 ;
        RECT 31.765 157.295 31.935 157.465 ;
        RECT 32.225 157.295 32.395 157.465 ;
        RECT 32.685 157.295 32.855 157.465 ;
        RECT 33.145 157.295 33.315 157.465 ;
        RECT 33.605 157.295 33.775 157.465 ;
        RECT 34.065 157.295 34.235 157.465 ;
        RECT 34.525 157.295 34.695 157.465 ;
        RECT 34.985 157.295 35.155 157.465 ;
        RECT 35.445 157.295 35.615 157.465 ;
        RECT 35.905 157.295 36.075 157.465 ;
        RECT 36.365 157.295 36.535 157.465 ;
        RECT 36.825 157.295 36.995 157.465 ;
        RECT 37.285 157.295 37.455 157.465 ;
        RECT 37.745 157.295 37.915 157.465 ;
        RECT 38.205 157.295 38.375 157.465 ;
        RECT 38.665 157.295 38.835 157.465 ;
        RECT 39.125 157.295 39.295 157.465 ;
        RECT 39.585 157.295 39.755 157.465 ;
        RECT 40.045 157.295 40.215 157.465 ;
        RECT 40.505 157.295 40.675 157.465 ;
        RECT 40.965 157.295 41.135 157.465 ;
        RECT 41.425 157.295 41.595 157.465 ;
        RECT 41.885 157.295 42.055 157.465 ;
        RECT 42.345 157.295 42.515 157.465 ;
        RECT 42.805 157.295 42.975 157.465 ;
        RECT 43.265 157.295 43.435 157.465 ;
        RECT 43.725 157.295 43.895 157.465 ;
        RECT 44.185 157.295 44.355 157.465 ;
        RECT 44.645 157.295 44.815 157.465 ;
        RECT 45.105 157.295 45.275 157.465 ;
        RECT 45.565 157.295 45.735 157.465 ;
        RECT 46.025 157.295 46.195 157.465 ;
        RECT 46.485 157.295 46.655 157.465 ;
        RECT 46.945 157.295 47.115 157.465 ;
        RECT 47.405 157.295 47.575 157.465 ;
        RECT 47.865 157.295 48.035 157.465 ;
        RECT 48.325 157.295 48.495 157.465 ;
        RECT 48.785 157.295 48.955 157.465 ;
        RECT 49.245 157.295 49.415 157.465 ;
        RECT 49.705 157.295 49.875 157.465 ;
        RECT 50.165 157.295 50.335 157.465 ;
        RECT 50.625 157.295 50.795 157.465 ;
        RECT 51.085 157.295 51.255 157.465 ;
        RECT 51.545 157.295 51.715 157.465 ;
        RECT 52.005 157.295 52.175 157.465 ;
        RECT 52.465 157.295 52.635 157.465 ;
        RECT 52.925 157.295 53.095 157.465 ;
        RECT 53.385 157.295 53.555 157.465 ;
        RECT 53.845 157.295 54.015 157.465 ;
        RECT 54.305 157.295 54.475 157.465 ;
        RECT 54.765 157.295 54.935 157.465 ;
        RECT 55.225 157.295 55.395 157.465 ;
        RECT 55.685 157.295 55.855 157.465 ;
        RECT 56.145 157.295 56.315 157.465 ;
        RECT 56.605 157.295 56.775 157.465 ;
        RECT 57.065 157.295 57.235 157.465 ;
        RECT 57.525 157.295 57.695 157.465 ;
        RECT 57.985 157.295 58.155 157.465 ;
        RECT 58.445 157.295 58.615 157.465 ;
        RECT 58.905 157.295 59.075 157.465 ;
        RECT 59.365 157.295 59.535 157.465 ;
        RECT 59.825 157.295 59.995 157.465 ;
        RECT 60.285 157.295 60.455 157.465 ;
        RECT 60.745 157.295 60.915 157.465 ;
        RECT 61.205 157.295 61.375 157.465 ;
        RECT 61.665 157.295 61.835 157.465 ;
        RECT 62.125 157.295 62.295 157.465 ;
        RECT 62.585 157.295 62.755 157.465 ;
        RECT 63.045 157.295 63.215 157.465 ;
        RECT 63.505 157.295 63.675 157.465 ;
        RECT 63.965 157.295 64.135 157.465 ;
        RECT 64.425 157.295 64.595 157.465 ;
        RECT 64.885 157.295 65.055 157.465 ;
        RECT 65.345 157.295 65.515 157.465 ;
        RECT 65.805 157.295 65.975 157.465 ;
        RECT 66.265 157.295 66.435 157.465 ;
        RECT 66.725 157.295 66.895 157.465 ;
        RECT 67.185 157.295 67.355 157.465 ;
        RECT 67.645 157.295 67.815 157.465 ;
        RECT 68.105 157.295 68.275 157.465 ;
        RECT 68.565 157.295 68.735 157.465 ;
        RECT 69.025 157.295 69.195 157.465 ;
        RECT 69.485 157.295 69.655 157.465 ;
        RECT 69.945 157.295 70.115 157.465 ;
        RECT 70.405 157.295 70.575 157.465 ;
        RECT 70.865 157.295 71.035 157.465 ;
        RECT 71.325 157.295 71.495 157.465 ;
        RECT 71.785 157.295 71.955 157.465 ;
        RECT 72.245 157.295 72.415 157.465 ;
        RECT 72.705 157.295 72.875 157.465 ;
        RECT 73.165 157.295 73.335 157.465 ;
        RECT 73.625 157.295 73.795 157.465 ;
        RECT 74.085 157.295 74.255 157.465 ;
        RECT 74.545 157.295 74.715 157.465 ;
        RECT 75.005 157.295 75.175 157.465 ;
        RECT 75.465 157.295 75.635 157.465 ;
        RECT 75.925 157.295 76.095 157.465 ;
        RECT 76.385 157.295 76.555 157.465 ;
        RECT 76.845 157.295 77.015 157.465 ;
        RECT 77.305 157.295 77.475 157.465 ;
        RECT 77.765 157.295 77.935 157.465 ;
        RECT 78.225 157.295 78.395 157.465 ;
        RECT 78.685 157.295 78.855 157.465 ;
        RECT 79.145 157.295 79.315 157.465 ;
        RECT 79.605 157.295 79.775 157.465 ;
        RECT 80.065 157.295 80.235 157.465 ;
        RECT 80.525 157.295 80.695 157.465 ;
        RECT 80.985 157.295 81.155 157.465 ;
        RECT 81.445 157.295 81.615 157.465 ;
        RECT 81.905 157.295 82.075 157.465 ;
        RECT 82.365 157.295 82.535 157.465 ;
        RECT 82.825 157.295 82.995 157.465 ;
        RECT 83.285 157.295 83.455 157.465 ;
        RECT 83.745 157.295 83.915 157.465 ;
        RECT 84.205 157.295 84.375 157.465 ;
        RECT 84.665 157.295 84.835 157.465 ;
        RECT 85.125 157.295 85.295 157.465 ;
        RECT 85.585 157.295 85.755 157.465 ;
        RECT 86.045 157.295 86.215 157.465 ;
        RECT 86.505 157.295 86.675 157.465 ;
        RECT 86.965 157.295 87.135 157.465 ;
        RECT 87.425 157.295 87.595 157.465 ;
        RECT 87.885 157.295 88.055 157.465 ;
        RECT 88.345 157.295 88.515 157.465 ;
        RECT 88.805 157.295 88.975 157.465 ;
        RECT 89.265 157.295 89.435 157.465 ;
        RECT 89.725 157.295 89.895 157.465 ;
        RECT 90.185 157.295 90.355 157.465 ;
        RECT 90.645 157.295 90.815 157.465 ;
        RECT 91.105 157.295 91.275 157.465 ;
        RECT 91.565 157.295 91.735 157.465 ;
        RECT 92.025 157.295 92.195 157.465 ;
        RECT 32.710 156.445 32.880 156.615 ;
        RECT 32.225 156.105 32.395 156.275 ;
        RECT 33.105 156.105 33.275 156.275 ;
        RECT 33.560 155.425 33.730 155.595 ;
        RECT 34.810 156.445 34.980 156.615 ;
        RECT 34.295 156.105 34.465 156.275 ;
        RECT 36.380 156.445 36.550 156.615 ;
        RECT 36.815 156.105 36.985 156.275 ;
        RECT 39.125 156.785 39.295 156.955 ;
        RECT 40.990 156.445 41.160 156.615 ;
        RECT 40.505 155.765 40.675 155.935 ;
        RECT 41.385 156.105 41.555 156.275 ;
        RECT 41.840 155.765 42.010 155.935 ;
        RECT 43.090 156.445 43.260 156.615 ;
        RECT 42.575 156.105 42.745 156.275 ;
        RECT 44.660 156.445 44.830 156.615 ;
        RECT 45.095 156.105 45.265 156.275 ;
        RECT 47.405 156.785 47.575 156.955 ;
        RECT 49.705 156.785 49.875 156.955 ;
        RECT 52.015 156.105 52.185 156.275 ;
        RECT 52.450 156.445 52.620 156.615 ;
        RECT 54.020 156.445 54.190 156.615 ;
        RECT 54.535 156.105 54.705 156.275 ;
        RECT 55.270 155.765 55.440 155.935 ;
        RECT 55.725 156.105 55.895 156.275 ;
        RECT 56.120 156.445 56.290 156.615 ;
        RECT 60.770 156.445 60.940 156.615 ;
        RECT 56.605 155.765 56.775 155.935 ;
        RECT 60.285 155.765 60.455 155.935 ;
        RECT 61.165 156.105 61.335 156.275 ;
        RECT 61.620 155.425 61.790 155.595 ;
        RECT 62.870 156.445 63.040 156.615 ;
        RECT 62.355 156.105 62.525 156.275 ;
        RECT 64.440 156.445 64.610 156.615 ;
        RECT 64.875 156.105 65.045 156.275 ;
        RECT 67.185 156.785 67.355 156.955 ;
        RECT 72.710 156.445 72.880 156.615 ;
        RECT 72.245 156.105 72.415 156.275 ;
        RECT 73.625 155.765 73.795 155.935 ;
        RECT 73.170 155.425 73.340 155.595 ;
        RECT 75.030 156.445 75.200 156.615 ;
        RECT 74.570 155.425 74.740 155.595 ;
        RECT 76.410 156.445 76.580 156.615 ;
        RECT 76.410 155.425 76.580 155.595 ;
        RECT 80.065 156.785 80.235 156.955 ;
        RECT 18.425 154.575 18.595 154.745 ;
        RECT 18.885 154.575 19.055 154.745 ;
        RECT 19.345 154.575 19.515 154.745 ;
        RECT 19.805 154.575 19.975 154.745 ;
        RECT 20.265 154.575 20.435 154.745 ;
        RECT 20.725 154.575 20.895 154.745 ;
        RECT 21.185 154.575 21.355 154.745 ;
        RECT 21.645 154.575 21.815 154.745 ;
        RECT 22.105 154.575 22.275 154.745 ;
        RECT 22.565 154.575 22.735 154.745 ;
        RECT 23.025 154.575 23.195 154.745 ;
        RECT 23.485 154.575 23.655 154.745 ;
        RECT 23.945 154.575 24.115 154.745 ;
        RECT 24.405 154.575 24.575 154.745 ;
        RECT 24.865 154.575 25.035 154.745 ;
        RECT 25.325 154.575 25.495 154.745 ;
        RECT 25.785 154.575 25.955 154.745 ;
        RECT 26.245 154.575 26.415 154.745 ;
        RECT 26.705 154.575 26.875 154.745 ;
        RECT 27.165 154.575 27.335 154.745 ;
        RECT 27.625 154.575 27.795 154.745 ;
        RECT 28.085 154.575 28.255 154.745 ;
        RECT 28.545 154.575 28.715 154.745 ;
        RECT 29.005 154.575 29.175 154.745 ;
        RECT 29.465 154.575 29.635 154.745 ;
        RECT 29.925 154.575 30.095 154.745 ;
        RECT 30.385 154.575 30.555 154.745 ;
        RECT 30.845 154.575 31.015 154.745 ;
        RECT 31.305 154.575 31.475 154.745 ;
        RECT 31.765 154.575 31.935 154.745 ;
        RECT 32.225 154.575 32.395 154.745 ;
        RECT 32.685 154.575 32.855 154.745 ;
        RECT 33.145 154.575 33.315 154.745 ;
        RECT 33.605 154.575 33.775 154.745 ;
        RECT 34.065 154.575 34.235 154.745 ;
        RECT 34.525 154.575 34.695 154.745 ;
        RECT 34.985 154.575 35.155 154.745 ;
        RECT 35.445 154.575 35.615 154.745 ;
        RECT 35.905 154.575 36.075 154.745 ;
        RECT 36.365 154.575 36.535 154.745 ;
        RECT 36.825 154.575 36.995 154.745 ;
        RECT 37.285 154.575 37.455 154.745 ;
        RECT 37.745 154.575 37.915 154.745 ;
        RECT 38.205 154.575 38.375 154.745 ;
        RECT 38.665 154.575 38.835 154.745 ;
        RECT 39.125 154.575 39.295 154.745 ;
        RECT 39.585 154.575 39.755 154.745 ;
        RECT 40.045 154.575 40.215 154.745 ;
        RECT 40.505 154.575 40.675 154.745 ;
        RECT 40.965 154.575 41.135 154.745 ;
        RECT 41.425 154.575 41.595 154.745 ;
        RECT 41.885 154.575 42.055 154.745 ;
        RECT 42.345 154.575 42.515 154.745 ;
        RECT 42.805 154.575 42.975 154.745 ;
        RECT 43.265 154.575 43.435 154.745 ;
        RECT 43.725 154.575 43.895 154.745 ;
        RECT 44.185 154.575 44.355 154.745 ;
        RECT 44.645 154.575 44.815 154.745 ;
        RECT 45.105 154.575 45.275 154.745 ;
        RECT 45.565 154.575 45.735 154.745 ;
        RECT 46.025 154.575 46.195 154.745 ;
        RECT 46.485 154.575 46.655 154.745 ;
        RECT 46.945 154.575 47.115 154.745 ;
        RECT 47.405 154.575 47.575 154.745 ;
        RECT 47.865 154.575 48.035 154.745 ;
        RECT 48.325 154.575 48.495 154.745 ;
        RECT 48.785 154.575 48.955 154.745 ;
        RECT 49.245 154.575 49.415 154.745 ;
        RECT 49.705 154.575 49.875 154.745 ;
        RECT 50.165 154.575 50.335 154.745 ;
        RECT 50.625 154.575 50.795 154.745 ;
        RECT 51.085 154.575 51.255 154.745 ;
        RECT 51.545 154.575 51.715 154.745 ;
        RECT 52.005 154.575 52.175 154.745 ;
        RECT 52.465 154.575 52.635 154.745 ;
        RECT 52.925 154.575 53.095 154.745 ;
        RECT 53.385 154.575 53.555 154.745 ;
        RECT 53.845 154.575 54.015 154.745 ;
        RECT 54.305 154.575 54.475 154.745 ;
        RECT 54.765 154.575 54.935 154.745 ;
        RECT 55.225 154.575 55.395 154.745 ;
        RECT 55.685 154.575 55.855 154.745 ;
        RECT 56.145 154.575 56.315 154.745 ;
        RECT 56.605 154.575 56.775 154.745 ;
        RECT 57.065 154.575 57.235 154.745 ;
        RECT 57.525 154.575 57.695 154.745 ;
        RECT 57.985 154.575 58.155 154.745 ;
        RECT 58.445 154.575 58.615 154.745 ;
        RECT 58.905 154.575 59.075 154.745 ;
        RECT 59.365 154.575 59.535 154.745 ;
        RECT 59.825 154.575 59.995 154.745 ;
        RECT 60.285 154.575 60.455 154.745 ;
        RECT 60.745 154.575 60.915 154.745 ;
        RECT 61.205 154.575 61.375 154.745 ;
        RECT 61.665 154.575 61.835 154.745 ;
        RECT 62.125 154.575 62.295 154.745 ;
        RECT 62.585 154.575 62.755 154.745 ;
        RECT 63.045 154.575 63.215 154.745 ;
        RECT 63.505 154.575 63.675 154.745 ;
        RECT 63.965 154.575 64.135 154.745 ;
        RECT 64.425 154.575 64.595 154.745 ;
        RECT 64.885 154.575 65.055 154.745 ;
        RECT 65.345 154.575 65.515 154.745 ;
        RECT 65.805 154.575 65.975 154.745 ;
        RECT 66.265 154.575 66.435 154.745 ;
        RECT 66.725 154.575 66.895 154.745 ;
        RECT 67.185 154.575 67.355 154.745 ;
        RECT 67.645 154.575 67.815 154.745 ;
        RECT 68.105 154.575 68.275 154.745 ;
        RECT 68.565 154.575 68.735 154.745 ;
        RECT 69.025 154.575 69.195 154.745 ;
        RECT 69.485 154.575 69.655 154.745 ;
        RECT 69.945 154.575 70.115 154.745 ;
        RECT 70.405 154.575 70.575 154.745 ;
        RECT 70.865 154.575 71.035 154.745 ;
        RECT 71.325 154.575 71.495 154.745 ;
        RECT 71.785 154.575 71.955 154.745 ;
        RECT 72.245 154.575 72.415 154.745 ;
        RECT 72.705 154.575 72.875 154.745 ;
        RECT 73.165 154.575 73.335 154.745 ;
        RECT 73.625 154.575 73.795 154.745 ;
        RECT 74.085 154.575 74.255 154.745 ;
        RECT 74.545 154.575 74.715 154.745 ;
        RECT 75.005 154.575 75.175 154.745 ;
        RECT 75.465 154.575 75.635 154.745 ;
        RECT 75.925 154.575 76.095 154.745 ;
        RECT 76.385 154.575 76.555 154.745 ;
        RECT 76.845 154.575 77.015 154.745 ;
        RECT 77.305 154.575 77.475 154.745 ;
        RECT 77.765 154.575 77.935 154.745 ;
        RECT 78.225 154.575 78.395 154.745 ;
        RECT 78.685 154.575 78.855 154.745 ;
        RECT 79.145 154.575 79.315 154.745 ;
        RECT 79.605 154.575 79.775 154.745 ;
        RECT 80.065 154.575 80.235 154.745 ;
        RECT 80.525 154.575 80.695 154.745 ;
        RECT 80.985 154.575 81.155 154.745 ;
        RECT 81.445 154.575 81.615 154.745 ;
        RECT 81.905 154.575 82.075 154.745 ;
        RECT 82.365 154.575 82.535 154.745 ;
        RECT 82.825 154.575 82.995 154.745 ;
        RECT 83.285 154.575 83.455 154.745 ;
        RECT 83.745 154.575 83.915 154.745 ;
        RECT 84.205 154.575 84.375 154.745 ;
        RECT 84.665 154.575 84.835 154.745 ;
        RECT 85.125 154.575 85.295 154.745 ;
        RECT 85.585 154.575 85.755 154.745 ;
        RECT 86.045 154.575 86.215 154.745 ;
        RECT 86.505 154.575 86.675 154.745 ;
        RECT 86.965 154.575 87.135 154.745 ;
        RECT 87.425 154.575 87.595 154.745 ;
        RECT 87.885 154.575 88.055 154.745 ;
        RECT 88.345 154.575 88.515 154.745 ;
        RECT 88.805 154.575 88.975 154.745 ;
        RECT 89.265 154.575 89.435 154.745 ;
        RECT 89.725 154.575 89.895 154.745 ;
        RECT 90.185 154.575 90.355 154.745 ;
        RECT 90.645 154.575 90.815 154.745 ;
        RECT 91.105 154.575 91.275 154.745 ;
        RECT 91.565 154.575 91.735 154.745 ;
        RECT 92.025 154.575 92.195 154.745 ;
        RECT 18.425 151.855 18.595 152.025 ;
        RECT 18.885 151.855 19.055 152.025 ;
        RECT 19.345 151.855 19.515 152.025 ;
        RECT 19.805 151.855 19.975 152.025 ;
        RECT 20.265 151.855 20.435 152.025 ;
        RECT 20.725 151.855 20.895 152.025 ;
        RECT 21.185 151.855 21.355 152.025 ;
        RECT 21.645 151.855 21.815 152.025 ;
        RECT 22.105 151.855 22.275 152.025 ;
        RECT 22.565 151.855 22.735 152.025 ;
        RECT 23.025 151.855 23.195 152.025 ;
        RECT 23.485 151.855 23.655 152.025 ;
        RECT 23.945 151.855 24.115 152.025 ;
        RECT 24.405 151.855 24.575 152.025 ;
        RECT 24.865 151.855 25.035 152.025 ;
        RECT 25.325 151.855 25.495 152.025 ;
        RECT 25.785 151.855 25.955 152.025 ;
        RECT 26.245 151.855 26.415 152.025 ;
        RECT 26.705 151.855 26.875 152.025 ;
        RECT 27.165 151.855 27.335 152.025 ;
        RECT 27.625 151.855 27.795 152.025 ;
        RECT 28.085 151.855 28.255 152.025 ;
        RECT 28.545 151.855 28.715 152.025 ;
        RECT 29.005 151.855 29.175 152.025 ;
        RECT 29.465 151.855 29.635 152.025 ;
        RECT 29.925 151.855 30.095 152.025 ;
        RECT 30.385 151.855 30.555 152.025 ;
        RECT 30.845 151.855 31.015 152.025 ;
        RECT 31.305 151.855 31.475 152.025 ;
        RECT 31.765 151.855 31.935 152.025 ;
        RECT 32.225 151.855 32.395 152.025 ;
        RECT 32.685 151.855 32.855 152.025 ;
        RECT 33.145 151.855 33.315 152.025 ;
        RECT 33.605 151.855 33.775 152.025 ;
        RECT 34.065 151.855 34.235 152.025 ;
        RECT 34.525 151.855 34.695 152.025 ;
        RECT 34.985 151.855 35.155 152.025 ;
        RECT 35.445 151.855 35.615 152.025 ;
        RECT 35.905 151.855 36.075 152.025 ;
        RECT 36.365 151.855 36.535 152.025 ;
        RECT 36.825 151.855 36.995 152.025 ;
        RECT 37.285 151.855 37.455 152.025 ;
        RECT 37.745 151.855 37.915 152.025 ;
        RECT 38.205 151.855 38.375 152.025 ;
        RECT 38.665 151.855 38.835 152.025 ;
        RECT 39.125 151.855 39.295 152.025 ;
        RECT 39.585 151.855 39.755 152.025 ;
        RECT 40.045 151.855 40.215 152.025 ;
        RECT 40.505 151.855 40.675 152.025 ;
        RECT 40.965 151.855 41.135 152.025 ;
        RECT 41.425 151.855 41.595 152.025 ;
        RECT 41.885 151.855 42.055 152.025 ;
        RECT 42.345 151.855 42.515 152.025 ;
        RECT 42.805 151.855 42.975 152.025 ;
        RECT 43.265 151.855 43.435 152.025 ;
        RECT 43.725 151.855 43.895 152.025 ;
        RECT 44.185 151.855 44.355 152.025 ;
        RECT 44.645 151.855 44.815 152.025 ;
        RECT 45.105 151.855 45.275 152.025 ;
        RECT 45.565 151.855 45.735 152.025 ;
        RECT 46.025 151.855 46.195 152.025 ;
        RECT 46.485 151.855 46.655 152.025 ;
        RECT 46.945 151.855 47.115 152.025 ;
        RECT 47.405 151.855 47.575 152.025 ;
        RECT 47.865 151.855 48.035 152.025 ;
        RECT 48.325 151.855 48.495 152.025 ;
        RECT 48.785 151.855 48.955 152.025 ;
        RECT 49.245 151.855 49.415 152.025 ;
        RECT 49.705 151.855 49.875 152.025 ;
        RECT 50.165 151.855 50.335 152.025 ;
        RECT 50.625 151.855 50.795 152.025 ;
        RECT 51.085 151.855 51.255 152.025 ;
        RECT 51.545 151.855 51.715 152.025 ;
        RECT 52.005 151.855 52.175 152.025 ;
        RECT 52.465 151.855 52.635 152.025 ;
        RECT 52.925 151.855 53.095 152.025 ;
        RECT 53.385 151.855 53.555 152.025 ;
        RECT 53.845 151.855 54.015 152.025 ;
        RECT 54.305 151.855 54.475 152.025 ;
        RECT 54.765 151.855 54.935 152.025 ;
        RECT 55.225 151.855 55.395 152.025 ;
        RECT 55.685 151.855 55.855 152.025 ;
        RECT 56.145 151.855 56.315 152.025 ;
        RECT 56.605 151.855 56.775 152.025 ;
        RECT 57.065 151.855 57.235 152.025 ;
        RECT 57.525 151.855 57.695 152.025 ;
        RECT 57.985 151.855 58.155 152.025 ;
        RECT 58.445 151.855 58.615 152.025 ;
        RECT 58.905 151.855 59.075 152.025 ;
        RECT 59.365 151.855 59.535 152.025 ;
        RECT 59.825 151.855 59.995 152.025 ;
        RECT 60.285 151.855 60.455 152.025 ;
        RECT 60.745 151.855 60.915 152.025 ;
        RECT 61.205 151.855 61.375 152.025 ;
        RECT 61.665 151.855 61.835 152.025 ;
        RECT 62.125 151.855 62.295 152.025 ;
        RECT 62.585 151.855 62.755 152.025 ;
        RECT 63.045 151.855 63.215 152.025 ;
        RECT 63.505 151.855 63.675 152.025 ;
        RECT 63.965 151.855 64.135 152.025 ;
        RECT 64.425 151.855 64.595 152.025 ;
        RECT 64.885 151.855 65.055 152.025 ;
        RECT 65.345 151.855 65.515 152.025 ;
        RECT 65.805 151.855 65.975 152.025 ;
        RECT 66.265 151.855 66.435 152.025 ;
        RECT 66.725 151.855 66.895 152.025 ;
        RECT 67.185 151.855 67.355 152.025 ;
        RECT 67.645 151.855 67.815 152.025 ;
        RECT 68.105 151.855 68.275 152.025 ;
        RECT 68.565 151.855 68.735 152.025 ;
        RECT 69.025 151.855 69.195 152.025 ;
        RECT 69.485 151.855 69.655 152.025 ;
        RECT 69.945 151.855 70.115 152.025 ;
        RECT 70.405 151.855 70.575 152.025 ;
        RECT 70.865 151.855 71.035 152.025 ;
        RECT 71.325 151.855 71.495 152.025 ;
        RECT 71.785 151.855 71.955 152.025 ;
        RECT 72.245 151.855 72.415 152.025 ;
        RECT 72.705 151.855 72.875 152.025 ;
        RECT 73.165 151.855 73.335 152.025 ;
        RECT 73.625 151.855 73.795 152.025 ;
        RECT 74.085 151.855 74.255 152.025 ;
        RECT 74.545 151.855 74.715 152.025 ;
        RECT 75.005 151.855 75.175 152.025 ;
        RECT 75.465 151.855 75.635 152.025 ;
        RECT 75.925 151.855 76.095 152.025 ;
        RECT 76.385 151.855 76.555 152.025 ;
        RECT 76.845 151.855 77.015 152.025 ;
        RECT 77.305 151.855 77.475 152.025 ;
        RECT 77.765 151.855 77.935 152.025 ;
        RECT 78.225 151.855 78.395 152.025 ;
        RECT 78.685 151.855 78.855 152.025 ;
        RECT 79.145 151.855 79.315 152.025 ;
        RECT 79.605 151.855 79.775 152.025 ;
        RECT 80.065 151.855 80.235 152.025 ;
        RECT 80.525 151.855 80.695 152.025 ;
        RECT 80.985 151.855 81.155 152.025 ;
        RECT 81.445 151.855 81.615 152.025 ;
        RECT 81.905 151.855 82.075 152.025 ;
        RECT 82.365 151.855 82.535 152.025 ;
        RECT 82.825 151.855 82.995 152.025 ;
        RECT 83.285 151.855 83.455 152.025 ;
        RECT 83.745 151.855 83.915 152.025 ;
        RECT 84.205 151.855 84.375 152.025 ;
        RECT 84.665 151.855 84.835 152.025 ;
        RECT 85.125 151.855 85.295 152.025 ;
        RECT 85.585 151.855 85.755 152.025 ;
        RECT 86.045 151.855 86.215 152.025 ;
        RECT 86.505 151.855 86.675 152.025 ;
        RECT 86.965 151.855 87.135 152.025 ;
        RECT 87.425 151.855 87.595 152.025 ;
        RECT 87.885 151.855 88.055 152.025 ;
        RECT 88.345 151.855 88.515 152.025 ;
        RECT 88.805 151.855 88.975 152.025 ;
        RECT 89.265 151.855 89.435 152.025 ;
        RECT 89.725 151.855 89.895 152.025 ;
        RECT 90.185 151.855 90.355 152.025 ;
        RECT 90.645 151.855 90.815 152.025 ;
        RECT 91.105 151.855 91.275 152.025 ;
        RECT 91.565 151.855 91.735 152.025 ;
        RECT 92.025 151.855 92.195 152.025 ;
        RECT 64.430 151.005 64.600 151.175 ;
        RECT 63.965 150.665 64.135 150.835 ;
        RECT 65.345 150.665 65.515 150.835 ;
        RECT 64.890 149.985 65.060 150.155 ;
        RECT 66.750 151.005 66.920 151.175 ;
        RECT 66.290 149.985 66.460 150.155 ;
        RECT 68.130 151.005 68.300 151.175 ;
        RECT 68.130 149.985 68.300 150.155 ;
        RECT 71.785 151.345 71.955 151.515 ;
        RECT 18.425 149.135 18.595 149.305 ;
        RECT 18.885 149.135 19.055 149.305 ;
        RECT 19.345 149.135 19.515 149.305 ;
        RECT 19.805 149.135 19.975 149.305 ;
        RECT 20.265 149.135 20.435 149.305 ;
        RECT 20.725 149.135 20.895 149.305 ;
        RECT 21.185 149.135 21.355 149.305 ;
        RECT 21.645 149.135 21.815 149.305 ;
        RECT 22.105 149.135 22.275 149.305 ;
        RECT 22.565 149.135 22.735 149.305 ;
        RECT 23.025 149.135 23.195 149.305 ;
        RECT 23.485 149.135 23.655 149.305 ;
        RECT 23.945 149.135 24.115 149.305 ;
        RECT 24.405 149.135 24.575 149.305 ;
        RECT 24.865 149.135 25.035 149.305 ;
        RECT 25.325 149.135 25.495 149.305 ;
        RECT 25.785 149.135 25.955 149.305 ;
        RECT 26.245 149.135 26.415 149.305 ;
        RECT 26.705 149.135 26.875 149.305 ;
        RECT 27.165 149.135 27.335 149.305 ;
        RECT 27.625 149.135 27.795 149.305 ;
        RECT 28.085 149.135 28.255 149.305 ;
        RECT 28.545 149.135 28.715 149.305 ;
        RECT 29.005 149.135 29.175 149.305 ;
        RECT 29.465 149.135 29.635 149.305 ;
        RECT 29.925 149.135 30.095 149.305 ;
        RECT 30.385 149.135 30.555 149.305 ;
        RECT 30.845 149.135 31.015 149.305 ;
        RECT 31.305 149.135 31.475 149.305 ;
        RECT 31.765 149.135 31.935 149.305 ;
        RECT 32.225 149.135 32.395 149.305 ;
        RECT 32.685 149.135 32.855 149.305 ;
        RECT 33.145 149.135 33.315 149.305 ;
        RECT 33.605 149.135 33.775 149.305 ;
        RECT 34.065 149.135 34.235 149.305 ;
        RECT 34.525 149.135 34.695 149.305 ;
        RECT 34.985 149.135 35.155 149.305 ;
        RECT 35.445 149.135 35.615 149.305 ;
        RECT 35.905 149.135 36.075 149.305 ;
        RECT 36.365 149.135 36.535 149.305 ;
        RECT 36.825 149.135 36.995 149.305 ;
        RECT 37.285 149.135 37.455 149.305 ;
        RECT 37.745 149.135 37.915 149.305 ;
        RECT 38.205 149.135 38.375 149.305 ;
        RECT 38.665 149.135 38.835 149.305 ;
        RECT 39.125 149.135 39.295 149.305 ;
        RECT 39.585 149.135 39.755 149.305 ;
        RECT 40.045 149.135 40.215 149.305 ;
        RECT 40.505 149.135 40.675 149.305 ;
        RECT 40.965 149.135 41.135 149.305 ;
        RECT 41.425 149.135 41.595 149.305 ;
        RECT 41.885 149.135 42.055 149.305 ;
        RECT 42.345 149.135 42.515 149.305 ;
        RECT 42.805 149.135 42.975 149.305 ;
        RECT 43.265 149.135 43.435 149.305 ;
        RECT 43.725 149.135 43.895 149.305 ;
        RECT 44.185 149.135 44.355 149.305 ;
        RECT 44.645 149.135 44.815 149.305 ;
        RECT 45.105 149.135 45.275 149.305 ;
        RECT 45.565 149.135 45.735 149.305 ;
        RECT 46.025 149.135 46.195 149.305 ;
        RECT 46.485 149.135 46.655 149.305 ;
        RECT 46.945 149.135 47.115 149.305 ;
        RECT 47.405 149.135 47.575 149.305 ;
        RECT 47.865 149.135 48.035 149.305 ;
        RECT 48.325 149.135 48.495 149.305 ;
        RECT 48.785 149.135 48.955 149.305 ;
        RECT 49.245 149.135 49.415 149.305 ;
        RECT 49.705 149.135 49.875 149.305 ;
        RECT 50.165 149.135 50.335 149.305 ;
        RECT 50.625 149.135 50.795 149.305 ;
        RECT 51.085 149.135 51.255 149.305 ;
        RECT 51.545 149.135 51.715 149.305 ;
        RECT 52.005 149.135 52.175 149.305 ;
        RECT 52.465 149.135 52.635 149.305 ;
        RECT 52.925 149.135 53.095 149.305 ;
        RECT 53.385 149.135 53.555 149.305 ;
        RECT 53.845 149.135 54.015 149.305 ;
        RECT 54.305 149.135 54.475 149.305 ;
        RECT 54.765 149.135 54.935 149.305 ;
        RECT 55.225 149.135 55.395 149.305 ;
        RECT 55.685 149.135 55.855 149.305 ;
        RECT 56.145 149.135 56.315 149.305 ;
        RECT 56.605 149.135 56.775 149.305 ;
        RECT 57.065 149.135 57.235 149.305 ;
        RECT 57.525 149.135 57.695 149.305 ;
        RECT 57.985 149.135 58.155 149.305 ;
        RECT 58.445 149.135 58.615 149.305 ;
        RECT 58.905 149.135 59.075 149.305 ;
        RECT 59.365 149.135 59.535 149.305 ;
        RECT 59.825 149.135 59.995 149.305 ;
        RECT 60.285 149.135 60.455 149.305 ;
        RECT 60.745 149.135 60.915 149.305 ;
        RECT 61.205 149.135 61.375 149.305 ;
        RECT 61.665 149.135 61.835 149.305 ;
        RECT 62.125 149.135 62.295 149.305 ;
        RECT 62.585 149.135 62.755 149.305 ;
        RECT 63.045 149.135 63.215 149.305 ;
        RECT 63.505 149.135 63.675 149.305 ;
        RECT 63.965 149.135 64.135 149.305 ;
        RECT 64.425 149.135 64.595 149.305 ;
        RECT 64.885 149.135 65.055 149.305 ;
        RECT 65.345 149.135 65.515 149.305 ;
        RECT 65.805 149.135 65.975 149.305 ;
        RECT 66.265 149.135 66.435 149.305 ;
        RECT 66.725 149.135 66.895 149.305 ;
        RECT 67.185 149.135 67.355 149.305 ;
        RECT 67.645 149.135 67.815 149.305 ;
        RECT 68.105 149.135 68.275 149.305 ;
        RECT 68.565 149.135 68.735 149.305 ;
        RECT 69.025 149.135 69.195 149.305 ;
        RECT 69.485 149.135 69.655 149.305 ;
        RECT 69.945 149.135 70.115 149.305 ;
        RECT 70.405 149.135 70.575 149.305 ;
        RECT 70.865 149.135 71.035 149.305 ;
        RECT 71.325 149.135 71.495 149.305 ;
        RECT 71.785 149.135 71.955 149.305 ;
        RECT 72.245 149.135 72.415 149.305 ;
        RECT 72.705 149.135 72.875 149.305 ;
        RECT 73.165 149.135 73.335 149.305 ;
        RECT 73.625 149.135 73.795 149.305 ;
        RECT 74.085 149.135 74.255 149.305 ;
        RECT 74.545 149.135 74.715 149.305 ;
        RECT 75.005 149.135 75.175 149.305 ;
        RECT 75.465 149.135 75.635 149.305 ;
        RECT 75.925 149.135 76.095 149.305 ;
        RECT 76.385 149.135 76.555 149.305 ;
        RECT 76.845 149.135 77.015 149.305 ;
        RECT 77.305 149.135 77.475 149.305 ;
        RECT 77.765 149.135 77.935 149.305 ;
        RECT 78.225 149.135 78.395 149.305 ;
        RECT 78.685 149.135 78.855 149.305 ;
        RECT 79.145 149.135 79.315 149.305 ;
        RECT 79.605 149.135 79.775 149.305 ;
        RECT 80.065 149.135 80.235 149.305 ;
        RECT 80.525 149.135 80.695 149.305 ;
        RECT 80.985 149.135 81.155 149.305 ;
        RECT 81.445 149.135 81.615 149.305 ;
        RECT 81.905 149.135 82.075 149.305 ;
        RECT 82.365 149.135 82.535 149.305 ;
        RECT 82.825 149.135 82.995 149.305 ;
        RECT 83.285 149.135 83.455 149.305 ;
        RECT 83.745 149.135 83.915 149.305 ;
        RECT 84.205 149.135 84.375 149.305 ;
        RECT 84.665 149.135 84.835 149.305 ;
        RECT 85.125 149.135 85.295 149.305 ;
        RECT 85.585 149.135 85.755 149.305 ;
        RECT 86.045 149.135 86.215 149.305 ;
        RECT 86.505 149.135 86.675 149.305 ;
        RECT 86.965 149.135 87.135 149.305 ;
        RECT 87.425 149.135 87.595 149.305 ;
        RECT 87.885 149.135 88.055 149.305 ;
        RECT 88.345 149.135 88.515 149.305 ;
        RECT 88.805 149.135 88.975 149.305 ;
        RECT 89.265 149.135 89.435 149.305 ;
        RECT 89.725 149.135 89.895 149.305 ;
        RECT 90.185 149.135 90.355 149.305 ;
        RECT 90.645 149.135 90.815 149.305 ;
        RECT 91.105 149.135 91.275 149.305 ;
        RECT 91.565 149.135 91.735 149.305 ;
        RECT 92.025 149.135 92.195 149.305 ;
        RECT 18.425 146.415 18.595 146.585 ;
        RECT 18.885 146.415 19.055 146.585 ;
        RECT 19.345 146.415 19.515 146.585 ;
        RECT 19.805 146.415 19.975 146.585 ;
        RECT 20.265 146.415 20.435 146.585 ;
        RECT 20.725 146.415 20.895 146.585 ;
        RECT 21.185 146.415 21.355 146.585 ;
        RECT 21.645 146.415 21.815 146.585 ;
        RECT 22.105 146.415 22.275 146.585 ;
        RECT 22.565 146.415 22.735 146.585 ;
        RECT 23.025 146.415 23.195 146.585 ;
        RECT 23.485 146.415 23.655 146.585 ;
        RECT 23.945 146.415 24.115 146.585 ;
        RECT 24.405 146.415 24.575 146.585 ;
        RECT 24.865 146.415 25.035 146.585 ;
        RECT 25.325 146.415 25.495 146.585 ;
        RECT 25.785 146.415 25.955 146.585 ;
        RECT 26.245 146.415 26.415 146.585 ;
        RECT 26.705 146.415 26.875 146.585 ;
        RECT 27.165 146.415 27.335 146.585 ;
        RECT 27.625 146.415 27.795 146.585 ;
        RECT 28.085 146.415 28.255 146.585 ;
        RECT 28.545 146.415 28.715 146.585 ;
        RECT 29.005 146.415 29.175 146.585 ;
        RECT 29.465 146.415 29.635 146.585 ;
        RECT 29.925 146.415 30.095 146.585 ;
        RECT 30.385 146.415 30.555 146.585 ;
        RECT 30.845 146.415 31.015 146.585 ;
        RECT 31.305 146.415 31.475 146.585 ;
        RECT 31.765 146.415 31.935 146.585 ;
        RECT 32.225 146.415 32.395 146.585 ;
        RECT 32.685 146.415 32.855 146.585 ;
        RECT 33.145 146.415 33.315 146.585 ;
        RECT 33.605 146.415 33.775 146.585 ;
        RECT 34.065 146.415 34.235 146.585 ;
        RECT 34.525 146.415 34.695 146.585 ;
        RECT 34.985 146.415 35.155 146.585 ;
        RECT 35.445 146.415 35.615 146.585 ;
        RECT 35.905 146.415 36.075 146.585 ;
        RECT 36.365 146.415 36.535 146.585 ;
        RECT 36.825 146.415 36.995 146.585 ;
        RECT 37.285 146.415 37.455 146.585 ;
        RECT 37.745 146.415 37.915 146.585 ;
        RECT 38.205 146.415 38.375 146.585 ;
        RECT 38.665 146.415 38.835 146.585 ;
        RECT 39.125 146.415 39.295 146.585 ;
        RECT 39.585 146.415 39.755 146.585 ;
        RECT 40.045 146.415 40.215 146.585 ;
        RECT 40.505 146.415 40.675 146.585 ;
        RECT 40.965 146.415 41.135 146.585 ;
        RECT 41.425 146.415 41.595 146.585 ;
        RECT 41.885 146.415 42.055 146.585 ;
        RECT 42.345 146.415 42.515 146.585 ;
        RECT 42.805 146.415 42.975 146.585 ;
        RECT 43.265 146.415 43.435 146.585 ;
        RECT 43.725 146.415 43.895 146.585 ;
        RECT 44.185 146.415 44.355 146.585 ;
        RECT 44.645 146.415 44.815 146.585 ;
        RECT 45.105 146.415 45.275 146.585 ;
        RECT 45.565 146.415 45.735 146.585 ;
        RECT 46.025 146.415 46.195 146.585 ;
        RECT 46.485 146.415 46.655 146.585 ;
        RECT 46.945 146.415 47.115 146.585 ;
        RECT 47.405 146.415 47.575 146.585 ;
        RECT 47.865 146.415 48.035 146.585 ;
        RECT 48.325 146.415 48.495 146.585 ;
        RECT 48.785 146.415 48.955 146.585 ;
        RECT 49.245 146.415 49.415 146.585 ;
        RECT 49.705 146.415 49.875 146.585 ;
        RECT 50.165 146.415 50.335 146.585 ;
        RECT 50.625 146.415 50.795 146.585 ;
        RECT 51.085 146.415 51.255 146.585 ;
        RECT 51.545 146.415 51.715 146.585 ;
        RECT 52.005 146.415 52.175 146.585 ;
        RECT 52.465 146.415 52.635 146.585 ;
        RECT 52.925 146.415 53.095 146.585 ;
        RECT 53.385 146.415 53.555 146.585 ;
        RECT 53.845 146.415 54.015 146.585 ;
        RECT 54.305 146.415 54.475 146.585 ;
        RECT 54.765 146.415 54.935 146.585 ;
        RECT 55.225 146.415 55.395 146.585 ;
        RECT 55.685 146.415 55.855 146.585 ;
        RECT 56.145 146.415 56.315 146.585 ;
        RECT 56.605 146.415 56.775 146.585 ;
        RECT 57.065 146.415 57.235 146.585 ;
        RECT 57.525 146.415 57.695 146.585 ;
        RECT 57.985 146.415 58.155 146.585 ;
        RECT 58.445 146.415 58.615 146.585 ;
        RECT 58.905 146.415 59.075 146.585 ;
        RECT 59.365 146.415 59.535 146.585 ;
        RECT 59.825 146.415 59.995 146.585 ;
        RECT 60.285 146.415 60.455 146.585 ;
        RECT 60.745 146.415 60.915 146.585 ;
        RECT 61.205 146.415 61.375 146.585 ;
        RECT 61.665 146.415 61.835 146.585 ;
        RECT 62.125 146.415 62.295 146.585 ;
        RECT 62.585 146.415 62.755 146.585 ;
        RECT 63.045 146.415 63.215 146.585 ;
        RECT 63.505 146.415 63.675 146.585 ;
        RECT 63.965 146.415 64.135 146.585 ;
        RECT 64.425 146.415 64.595 146.585 ;
        RECT 64.885 146.415 65.055 146.585 ;
        RECT 65.345 146.415 65.515 146.585 ;
        RECT 65.805 146.415 65.975 146.585 ;
        RECT 66.265 146.415 66.435 146.585 ;
        RECT 66.725 146.415 66.895 146.585 ;
        RECT 67.185 146.415 67.355 146.585 ;
        RECT 67.645 146.415 67.815 146.585 ;
        RECT 68.105 146.415 68.275 146.585 ;
        RECT 68.565 146.415 68.735 146.585 ;
        RECT 69.025 146.415 69.195 146.585 ;
        RECT 69.485 146.415 69.655 146.585 ;
        RECT 69.945 146.415 70.115 146.585 ;
        RECT 70.405 146.415 70.575 146.585 ;
        RECT 70.865 146.415 71.035 146.585 ;
        RECT 71.325 146.415 71.495 146.585 ;
        RECT 71.785 146.415 71.955 146.585 ;
        RECT 72.245 146.415 72.415 146.585 ;
        RECT 72.705 146.415 72.875 146.585 ;
        RECT 73.165 146.415 73.335 146.585 ;
        RECT 73.625 146.415 73.795 146.585 ;
        RECT 74.085 146.415 74.255 146.585 ;
        RECT 74.545 146.415 74.715 146.585 ;
        RECT 75.005 146.415 75.175 146.585 ;
        RECT 75.465 146.415 75.635 146.585 ;
        RECT 75.925 146.415 76.095 146.585 ;
        RECT 76.385 146.415 76.555 146.585 ;
        RECT 76.845 146.415 77.015 146.585 ;
        RECT 77.305 146.415 77.475 146.585 ;
        RECT 77.765 146.415 77.935 146.585 ;
        RECT 78.225 146.415 78.395 146.585 ;
        RECT 78.685 146.415 78.855 146.585 ;
        RECT 79.145 146.415 79.315 146.585 ;
        RECT 79.605 146.415 79.775 146.585 ;
        RECT 80.065 146.415 80.235 146.585 ;
        RECT 80.525 146.415 80.695 146.585 ;
        RECT 80.985 146.415 81.155 146.585 ;
        RECT 81.445 146.415 81.615 146.585 ;
        RECT 81.905 146.415 82.075 146.585 ;
        RECT 82.365 146.415 82.535 146.585 ;
        RECT 82.825 146.415 82.995 146.585 ;
        RECT 83.285 146.415 83.455 146.585 ;
        RECT 83.745 146.415 83.915 146.585 ;
        RECT 84.205 146.415 84.375 146.585 ;
        RECT 84.665 146.415 84.835 146.585 ;
        RECT 85.125 146.415 85.295 146.585 ;
        RECT 85.585 146.415 85.755 146.585 ;
        RECT 86.045 146.415 86.215 146.585 ;
        RECT 86.505 146.415 86.675 146.585 ;
        RECT 86.965 146.415 87.135 146.585 ;
        RECT 87.425 146.415 87.595 146.585 ;
        RECT 87.885 146.415 88.055 146.585 ;
        RECT 88.345 146.415 88.515 146.585 ;
        RECT 88.805 146.415 88.975 146.585 ;
        RECT 89.265 146.415 89.435 146.585 ;
        RECT 89.725 146.415 89.895 146.585 ;
        RECT 90.185 146.415 90.355 146.585 ;
        RECT 90.645 146.415 90.815 146.585 ;
        RECT 91.105 146.415 91.275 146.585 ;
        RECT 91.565 146.415 91.735 146.585 ;
        RECT 92.025 146.415 92.195 146.585 ;
        RECT 18.425 143.695 18.595 143.865 ;
        RECT 18.885 143.695 19.055 143.865 ;
        RECT 19.345 143.695 19.515 143.865 ;
        RECT 19.805 143.695 19.975 143.865 ;
        RECT 20.265 143.695 20.435 143.865 ;
        RECT 20.725 143.695 20.895 143.865 ;
        RECT 21.185 143.695 21.355 143.865 ;
        RECT 21.645 143.695 21.815 143.865 ;
        RECT 22.105 143.695 22.275 143.865 ;
        RECT 22.565 143.695 22.735 143.865 ;
        RECT 23.025 143.695 23.195 143.865 ;
        RECT 23.485 143.695 23.655 143.865 ;
        RECT 23.945 143.695 24.115 143.865 ;
        RECT 24.405 143.695 24.575 143.865 ;
        RECT 24.865 143.695 25.035 143.865 ;
        RECT 25.325 143.695 25.495 143.865 ;
        RECT 25.785 143.695 25.955 143.865 ;
        RECT 26.245 143.695 26.415 143.865 ;
        RECT 26.705 143.695 26.875 143.865 ;
        RECT 27.165 143.695 27.335 143.865 ;
        RECT 27.625 143.695 27.795 143.865 ;
        RECT 28.085 143.695 28.255 143.865 ;
        RECT 28.545 143.695 28.715 143.865 ;
        RECT 29.005 143.695 29.175 143.865 ;
        RECT 29.465 143.695 29.635 143.865 ;
        RECT 29.925 143.695 30.095 143.865 ;
        RECT 30.385 143.695 30.555 143.865 ;
        RECT 30.845 143.695 31.015 143.865 ;
        RECT 31.305 143.695 31.475 143.865 ;
        RECT 31.765 143.695 31.935 143.865 ;
        RECT 32.225 143.695 32.395 143.865 ;
        RECT 32.685 143.695 32.855 143.865 ;
        RECT 33.145 143.695 33.315 143.865 ;
        RECT 33.605 143.695 33.775 143.865 ;
        RECT 34.065 143.695 34.235 143.865 ;
        RECT 34.525 143.695 34.695 143.865 ;
        RECT 34.985 143.695 35.155 143.865 ;
        RECT 35.445 143.695 35.615 143.865 ;
        RECT 35.905 143.695 36.075 143.865 ;
        RECT 36.365 143.695 36.535 143.865 ;
        RECT 36.825 143.695 36.995 143.865 ;
        RECT 37.285 143.695 37.455 143.865 ;
        RECT 37.745 143.695 37.915 143.865 ;
        RECT 38.205 143.695 38.375 143.865 ;
        RECT 38.665 143.695 38.835 143.865 ;
        RECT 39.125 143.695 39.295 143.865 ;
        RECT 39.585 143.695 39.755 143.865 ;
        RECT 40.045 143.695 40.215 143.865 ;
        RECT 40.505 143.695 40.675 143.865 ;
        RECT 40.965 143.695 41.135 143.865 ;
        RECT 41.425 143.695 41.595 143.865 ;
        RECT 41.885 143.695 42.055 143.865 ;
        RECT 42.345 143.695 42.515 143.865 ;
        RECT 42.805 143.695 42.975 143.865 ;
        RECT 43.265 143.695 43.435 143.865 ;
        RECT 43.725 143.695 43.895 143.865 ;
        RECT 44.185 143.695 44.355 143.865 ;
        RECT 44.645 143.695 44.815 143.865 ;
        RECT 45.105 143.695 45.275 143.865 ;
        RECT 45.565 143.695 45.735 143.865 ;
        RECT 46.025 143.695 46.195 143.865 ;
        RECT 46.485 143.695 46.655 143.865 ;
        RECT 46.945 143.695 47.115 143.865 ;
        RECT 47.405 143.695 47.575 143.865 ;
        RECT 47.865 143.695 48.035 143.865 ;
        RECT 48.325 143.695 48.495 143.865 ;
        RECT 48.785 143.695 48.955 143.865 ;
        RECT 49.245 143.695 49.415 143.865 ;
        RECT 49.705 143.695 49.875 143.865 ;
        RECT 50.165 143.695 50.335 143.865 ;
        RECT 50.625 143.695 50.795 143.865 ;
        RECT 51.085 143.695 51.255 143.865 ;
        RECT 51.545 143.695 51.715 143.865 ;
        RECT 52.005 143.695 52.175 143.865 ;
        RECT 52.465 143.695 52.635 143.865 ;
        RECT 52.925 143.695 53.095 143.865 ;
        RECT 53.385 143.695 53.555 143.865 ;
        RECT 53.845 143.695 54.015 143.865 ;
        RECT 54.305 143.695 54.475 143.865 ;
        RECT 54.765 143.695 54.935 143.865 ;
        RECT 55.225 143.695 55.395 143.865 ;
        RECT 55.685 143.695 55.855 143.865 ;
        RECT 56.145 143.695 56.315 143.865 ;
        RECT 56.605 143.695 56.775 143.865 ;
        RECT 57.065 143.695 57.235 143.865 ;
        RECT 57.525 143.695 57.695 143.865 ;
        RECT 57.985 143.695 58.155 143.865 ;
        RECT 58.445 143.695 58.615 143.865 ;
        RECT 58.905 143.695 59.075 143.865 ;
        RECT 59.365 143.695 59.535 143.865 ;
        RECT 59.825 143.695 59.995 143.865 ;
        RECT 60.285 143.695 60.455 143.865 ;
        RECT 60.745 143.695 60.915 143.865 ;
        RECT 61.205 143.695 61.375 143.865 ;
        RECT 61.665 143.695 61.835 143.865 ;
        RECT 62.125 143.695 62.295 143.865 ;
        RECT 62.585 143.695 62.755 143.865 ;
        RECT 63.045 143.695 63.215 143.865 ;
        RECT 63.505 143.695 63.675 143.865 ;
        RECT 63.965 143.695 64.135 143.865 ;
        RECT 64.425 143.695 64.595 143.865 ;
        RECT 64.885 143.695 65.055 143.865 ;
        RECT 65.345 143.695 65.515 143.865 ;
        RECT 65.805 143.695 65.975 143.865 ;
        RECT 66.265 143.695 66.435 143.865 ;
        RECT 66.725 143.695 66.895 143.865 ;
        RECT 67.185 143.695 67.355 143.865 ;
        RECT 67.645 143.695 67.815 143.865 ;
        RECT 68.105 143.695 68.275 143.865 ;
        RECT 68.565 143.695 68.735 143.865 ;
        RECT 69.025 143.695 69.195 143.865 ;
        RECT 69.485 143.695 69.655 143.865 ;
        RECT 69.945 143.695 70.115 143.865 ;
        RECT 70.405 143.695 70.575 143.865 ;
        RECT 70.865 143.695 71.035 143.865 ;
        RECT 71.325 143.695 71.495 143.865 ;
        RECT 71.785 143.695 71.955 143.865 ;
        RECT 72.245 143.695 72.415 143.865 ;
        RECT 72.705 143.695 72.875 143.865 ;
        RECT 73.165 143.695 73.335 143.865 ;
        RECT 73.625 143.695 73.795 143.865 ;
        RECT 74.085 143.695 74.255 143.865 ;
        RECT 74.545 143.695 74.715 143.865 ;
        RECT 75.005 143.695 75.175 143.865 ;
        RECT 75.465 143.695 75.635 143.865 ;
        RECT 75.925 143.695 76.095 143.865 ;
        RECT 76.385 143.695 76.555 143.865 ;
        RECT 76.845 143.695 77.015 143.865 ;
        RECT 77.305 143.695 77.475 143.865 ;
        RECT 77.765 143.695 77.935 143.865 ;
        RECT 78.225 143.695 78.395 143.865 ;
        RECT 78.685 143.695 78.855 143.865 ;
        RECT 79.145 143.695 79.315 143.865 ;
        RECT 79.605 143.695 79.775 143.865 ;
        RECT 80.065 143.695 80.235 143.865 ;
        RECT 80.525 143.695 80.695 143.865 ;
        RECT 80.985 143.695 81.155 143.865 ;
        RECT 81.445 143.695 81.615 143.865 ;
        RECT 81.905 143.695 82.075 143.865 ;
        RECT 82.365 143.695 82.535 143.865 ;
        RECT 82.825 143.695 82.995 143.865 ;
        RECT 83.285 143.695 83.455 143.865 ;
        RECT 83.745 143.695 83.915 143.865 ;
        RECT 84.205 143.695 84.375 143.865 ;
        RECT 84.665 143.695 84.835 143.865 ;
        RECT 85.125 143.695 85.295 143.865 ;
        RECT 85.585 143.695 85.755 143.865 ;
        RECT 86.045 143.695 86.215 143.865 ;
        RECT 86.505 143.695 86.675 143.865 ;
        RECT 86.965 143.695 87.135 143.865 ;
        RECT 87.425 143.695 87.595 143.865 ;
        RECT 87.885 143.695 88.055 143.865 ;
        RECT 88.345 143.695 88.515 143.865 ;
        RECT 88.805 143.695 88.975 143.865 ;
        RECT 89.265 143.695 89.435 143.865 ;
        RECT 89.725 143.695 89.895 143.865 ;
        RECT 90.185 143.695 90.355 143.865 ;
        RECT 90.645 143.695 90.815 143.865 ;
        RECT 91.105 143.695 91.275 143.865 ;
        RECT 91.565 143.695 91.735 143.865 ;
        RECT 92.025 143.695 92.195 143.865 ;
        RECT 113.070 142.775 113.260 144.760 ;
        RECT 114.070 142.775 114.260 144.760 ;
        RECT 115.070 142.775 115.260 144.760 ;
        RECT 116.070 142.775 116.260 144.760 ;
        RECT 117.070 142.775 117.260 144.760 ;
        RECT 118.070 142.775 118.260 144.760 ;
        RECT 119.070 142.775 119.260 144.760 ;
        RECT 120.070 142.775 120.260 144.760 ;
        RECT 18.425 140.975 18.595 141.145 ;
        RECT 18.885 140.975 19.055 141.145 ;
        RECT 19.345 140.975 19.515 141.145 ;
        RECT 19.805 140.975 19.975 141.145 ;
        RECT 20.265 140.975 20.435 141.145 ;
        RECT 20.725 140.975 20.895 141.145 ;
        RECT 21.185 140.975 21.355 141.145 ;
        RECT 21.645 140.975 21.815 141.145 ;
        RECT 22.105 140.975 22.275 141.145 ;
        RECT 22.565 140.975 22.735 141.145 ;
        RECT 23.025 140.975 23.195 141.145 ;
        RECT 23.485 140.975 23.655 141.145 ;
        RECT 23.945 140.975 24.115 141.145 ;
        RECT 24.405 140.975 24.575 141.145 ;
        RECT 24.865 140.975 25.035 141.145 ;
        RECT 25.325 140.975 25.495 141.145 ;
        RECT 25.785 140.975 25.955 141.145 ;
        RECT 26.245 140.975 26.415 141.145 ;
        RECT 26.705 140.975 26.875 141.145 ;
        RECT 27.165 140.975 27.335 141.145 ;
        RECT 27.625 140.975 27.795 141.145 ;
        RECT 28.085 140.975 28.255 141.145 ;
        RECT 28.545 140.975 28.715 141.145 ;
        RECT 29.005 140.975 29.175 141.145 ;
        RECT 29.465 140.975 29.635 141.145 ;
        RECT 29.925 140.975 30.095 141.145 ;
        RECT 30.385 140.975 30.555 141.145 ;
        RECT 30.845 140.975 31.015 141.145 ;
        RECT 31.305 140.975 31.475 141.145 ;
        RECT 31.765 140.975 31.935 141.145 ;
        RECT 32.225 140.975 32.395 141.145 ;
        RECT 32.685 140.975 32.855 141.145 ;
        RECT 33.145 140.975 33.315 141.145 ;
        RECT 33.605 140.975 33.775 141.145 ;
        RECT 34.065 140.975 34.235 141.145 ;
        RECT 34.525 140.975 34.695 141.145 ;
        RECT 34.985 140.975 35.155 141.145 ;
        RECT 35.445 140.975 35.615 141.145 ;
        RECT 35.905 140.975 36.075 141.145 ;
        RECT 36.365 140.975 36.535 141.145 ;
        RECT 36.825 140.975 36.995 141.145 ;
        RECT 37.285 140.975 37.455 141.145 ;
        RECT 37.745 140.975 37.915 141.145 ;
        RECT 38.205 140.975 38.375 141.145 ;
        RECT 38.665 140.975 38.835 141.145 ;
        RECT 39.125 140.975 39.295 141.145 ;
        RECT 39.585 140.975 39.755 141.145 ;
        RECT 40.045 140.975 40.215 141.145 ;
        RECT 40.505 140.975 40.675 141.145 ;
        RECT 40.965 140.975 41.135 141.145 ;
        RECT 41.425 140.975 41.595 141.145 ;
        RECT 41.885 140.975 42.055 141.145 ;
        RECT 42.345 140.975 42.515 141.145 ;
        RECT 42.805 140.975 42.975 141.145 ;
        RECT 43.265 140.975 43.435 141.145 ;
        RECT 43.725 140.975 43.895 141.145 ;
        RECT 44.185 140.975 44.355 141.145 ;
        RECT 44.645 140.975 44.815 141.145 ;
        RECT 45.105 140.975 45.275 141.145 ;
        RECT 45.565 140.975 45.735 141.145 ;
        RECT 46.025 140.975 46.195 141.145 ;
        RECT 46.485 140.975 46.655 141.145 ;
        RECT 46.945 140.975 47.115 141.145 ;
        RECT 47.405 140.975 47.575 141.145 ;
        RECT 47.865 140.975 48.035 141.145 ;
        RECT 48.325 140.975 48.495 141.145 ;
        RECT 48.785 140.975 48.955 141.145 ;
        RECT 49.245 140.975 49.415 141.145 ;
        RECT 49.705 140.975 49.875 141.145 ;
        RECT 50.165 140.975 50.335 141.145 ;
        RECT 50.625 140.975 50.795 141.145 ;
        RECT 51.085 140.975 51.255 141.145 ;
        RECT 51.545 140.975 51.715 141.145 ;
        RECT 52.005 140.975 52.175 141.145 ;
        RECT 52.465 140.975 52.635 141.145 ;
        RECT 52.925 140.975 53.095 141.145 ;
        RECT 53.385 140.975 53.555 141.145 ;
        RECT 53.845 140.975 54.015 141.145 ;
        RECT 54.305 140.975 54.475 141.145 ;
        RECT 54.765 140.975 54.935 141.145 ;
        RECT 55.225 140.975 55.395 141.145 ;
        RECT 55.685 140.975 55.855 141.145 ;
        RECT 56.145 140.975 56.315 141.145 ;
        RECT 56.605 140.975 56.775 141.145 ;
        RECT 57.065 140.975 57.235 141.145 ;
        RECT 57.525 140.975 57.695 141.145 ;
        RECT 57.985 140.975 58.155 141.145 ;
        RECT 58.445 140.975 58.615 141.145 ;
        RECT 58.905 140.975 59.075 141.145 ;
        RECT 59.365 140.975 59.535 141.145 ;
        RECT 59.825 140.975 59.995 141.145 ;
        RECT 60.285 140.975 60.455 141.145 ;
        RECT 60.745 140.975 60.915 141.145 ;
        RECT 61.205 140.975 61.375 141.145 ;
        RECT 61.665 140.975 61.835 141.145 ;
        RECT 62.125 140.975 62.295 141.145 ;
        RECT 62.585 140.975 62.755 141.145 ;
        RECT 63.045 140.975 63.215 141.145 ;
        RECT 63.505 140.975 63.675 141.145 ;
        RECT 63.965 140.975 64.135 141.145 ;
        RECT 64.425 140.975 64.595 141.145 ;
        RECT 64.885 140.975 65.055 141.145 ;
        RECT 65.345 140.975 65.515 141.145 ;
        RECT 65.805 140.975 65.975 141.145 ;
        RECT 66.265 140.975 66.435 141.145 ;
        RECT 66.725 140.975 66.895 141.145 ;
        RECT 67.185 140.975 67.355 141.145 ;
        RECT 67.645 140.975 67.815 141.145 ;
        RECT 68.105 140.975 68.275 141.145 ;
        RECT 68.565 140.975 68.735 141.145 ;
        RECT 69.025 140.975 69.195 141.145 ;
        RECT 69.485 140.975 69.655 141.145 ;
        RECT 69.945 140.975 70.115 141.145 ;
        RECT 70.405 140.975 70.575 141.145 ;
        RECT 70.865 140.975 71.035 141.145 ;
        RECT 71.325 140.975 71.495 141.145 ;
        RECT 71.785 140.975 71.955 141.145 ;
        RECT 72.245 140.975 72.415 141.145 ;
        RECT 72.705 140.975 72.875 141.145 ;
        RECT 73.165 140.975 73.335 141.145 ;
        RECT 73.625 140.975 73.795 141.145 ;
        RECT 74.085 140.975 74.255 141.145 ;
        RECT 74.545 140.975 74.715 141.145 ;
        RECT 75.005 140.975 75.175 141.145 ;
        RECT 75.465 140.975 75.635 141.145 ;
        RECT 75.925 140.975 76.095 141.145 ;
        RECT 76.385 140.975 76.555 141.145 ;
        RECT 76.845 140.975 77.015 141.145 ;
        RECT 77.305 140.975 77.475 141.145 ;
        RECT 77.765 140.975 77.935 141.145 ;
        RECT 78.225 140.975 78.395 141.145 ;
        RECT 78.685 140.975 78.855 141.145 ;
        RECT 79.145 140.975 79.315 141.145 ;
        RECT 79.605 140.975 79.775 141.145 ;
        RECT 80.065 140.975 80.235 141.145 ;
        RECT 80.525 140.975 80.695 141.145 ;
        RECT 80.985 140.975 81.155 141.145 ;
        RECT 81.445 140.975 81.615 141.145 ;
        RECT 81.905 140.975 82.075 141.145 ;
        RECT 82.365 140.975 82.535 141.145 ;
        RECT 82.825 140.975 82.995 141.145 ;
        RECT 83.285 140.975 83.455 141.145 ;
        RECT 83.745 140.975 83.915 141.145 ;
        RECT 84.205 140.975 84.375 141.145 ;
        RECT 84.665 140.975 84.835 141.145 ;
        RECT 85.125 140.975 85.295 141.145 ;
        RECT 85.585 140.975 85.755 141.145 ;
        RECT 86.045 140.975 86.215 141.145 ;
        RECT 86.505 140.975 86.675 141.145 ;
        RECT 86.965 140.975 87.135 141.145 ;
        RECT 87.425 140.975 87.595 141.145 ;
        RECT 87.885 140.975 88.055 141.145 ;
        RECT 88.345 140.975 88.515 141.145 ;
        RECT 88.805 140.975 88.975 141.145 ;
        RECT 89.265 140.975 89.435 141.145 ;
        RECT 89.725 140.975 89.895 141.145 ;
        RECT 90.185 140.975 90.355 141.145 ;
        RECT 90.645 140.975 90.815 141.145 ;
        RECT 91.105 140.975 91.275 141.145 ;
        RECT 91.565 140.975 91.735 141.145 ;
        RECT 92.025 140.975 92.195 141.145 ;
        RECT 113.070 139.620 113.260 141.605 ;
        RECT 114.070 139.620 114.260 141.605 ;
        RECT 115.070 139.620 115.260 141.605 ;
        RECT 116.070 139.620 116.260 141.605 ;
        RECT 117.070 139.620 117.260 141.605 ;
        RECT 118.070 139.620 118.260 141.605 ;
        RECT 119.070 139.620 119.260 141.605 ;
        RECT 120.070 139.620 120.260 141.605 ;
        RECT 18.425 138.255 18.595 138.425 ;
        RECT 18.885 138.255 19.055 138.425 ;
        RECT 19.345 138.255 19.515 138.425 ;
        RECT 19.805 138.255 19.975 138.425 ;
        RECT 20.265 138.255 20.435 138.425 ;
        RECT 20.725 138.255 20.895 138.425 ;
        RECT 21.185 138.255 21.355 138.425 ;
        RECT 21.645 138.255 21.815 138.425 ;
        RECT 22.105 138.255 22.275 138.425 ;
        RECT 22.565 138.255 22.735 138.425 ;
        RECT 23.025 138.255 23.195 138.425 ;
        RECT 23.485 138.255 23.655 138.425 ;
        RECT 23.945 138.255 24.115 138.425 ;
        RECT 24.405 138.255 24.575 138.425 ;
        RECT 24.865 138.255 25.035 138.425 ;
        RECT 25.325 138.255 25.495 138.425 ;
        RECT 25.785 138.255 25.955 138.425 ;
        RECT 26.245 138.255 26.415 138.425 ;
        RECT 26.705 138.255 26.875 138.425 ;
        RECT 27.165 138.255 27.335 138.425 ;
        RECT 27.625 138.255 27.795 138.425 ;
        RECT 28.085 138.255 28.255 138.425 ;
        RECT 28.545 138.255 28.715 138.425 ;
        RECT 29.005 138.255 29.175 138.425 ;
        RECT 29.465 138.255 29.635 138.425 ;
        RECT 29.925 138.255 30.095 138.425 ;
        RECT 30.385 138.255 30.555 138.425 ;
        RECT 30.845 138.255 31.015 138.425 ;
        RECT 31.305 138.255 31.475 138.425 ;
        RECT 31.765 138.255 31.935 138.425 ;
        RECT 32.225 138.255 32.395 138.425 ;
        RECT 32.685 138.255 32.855 138.425 ;
        RECT 33.145 138.255 33.315 138.425 ;
        RECT 33.605 138.255 33.775 138.425 ;
        RECT 34.065 138.255 34.235 138.425 ;
        RECT 34.525 138.255 34.695 138.425 ;
        RECT 34.985 138.255 35.155 138.425 ;
        RECT 35.445 138.255 35.615 138.425 ;
        RECT 35.905 138.255 36.075 138.425 ;
        RECT 36.365 138.255 36.535 138.425 ;
        RECT 36.825 138.255 36.995 138.425 ;
        RECT 37.285 138.255 37.455 138.425 ;
        RECT 37.745 138.255 37.915 138.425 ;
        RECT 38.205 138.255 38.375 138.425 ;
        RECT 38.665 138.255 38.835 138.425 ;
        RECT 39.125 138.255 39.295 138.425 ;
        RECT 39.585 138.255 39.755 138.425 ;
        RECT 40.045 138.255 40.215 138.425 ;
        RECT 40.505 138.255 40.675 138.425 ;
        RECT 40.965 138.255 41.135 138.425 ;
        RECT 41.425 138.255 41.595 138.425 ;
        RECT 41.885 138.255 42.055 138.425 ;
        RECT 42.345 138.255 42.515 138.425 ;
        RECT 42.805 138.255 42.975 138.425 ;
        RECT 43.265 138.255 43.435 138.425 ;
        RECT 43.725 138.255 43.895 138.425 ;
        RECT 44.185 138.255 44.355 138.425 ;
        RECT 44.645 138.255 44.815 138.425 ;
        RECT 45.105 138.255 45.275 138.425 ;
        RECT 45.565 138.255 45.735 138.425 ;
        RECT 46.025 138.255 46.195 138.425 ;
        RECT 46.485 138.255 46.655 138.425 ;
        RECT 46.945 138.255 47.115 138.425 ;
        RECT 47.405 138.255 47.575 138.425 ;
        RECT 47.865 138.255 48.035 138.425 ;
        RECT 48.325 138.255 48.495 138.425 ;
        RECT 48.785 138.255 48.955 138.425 ;
        RECT 49.245 138.255 49.415 138.425 ;
        RECT 49.705 138.255 49.875 138.425 ;
        RECT 50.165 138.255 50.335 138.425 ;
        RECT 50.625 138.255 50.795 138.425 ;
        RECT 51.085 138.255 51.255 138.425 ;
        RECT 51.545 138.255 51.715 138.425 ;
        RECT 52.005 138.255 52.175 138.425 ;
        RECT 52.465 138.255 52.635 138.425 ;
        RECT 52.925 138.255 53.095 138.425 ;
        RECT 53.385 138.255 53.555 138.425 ;
        RECT 53.845 138.255 54.015 138.425 ;
        RECT 54.305 138.255 54.475 138.425 ;
        RECT 54.765 138.255 54.935 138.425 ;
        RECT 55.225 138.255 55.395 138.425 ;
        RECT 55.685 138.255 55.855 138.425 ;
        RECT 56.145 138.255 56.315 138.425 ;
        RECT 56.605 138.255 56.775 138.425 ;
        RECT 57.065 138.255 57.235 138.425 ;
        RECT 57.525 138.255 57.695 138.425 ;
        RECT 57.985 138.255 58.155 138.425 ;
        RECT 58.445 138.255 58.615 138.425 ;
        RECT 58.905 138.255 59.075 138.425 ;
        RECT 59.365 138.255 59.535 138.425 ;
        RECT 59.825 138.255 59.995 138.425 ;
        RECT 60.285 138.255 60.455 138.425 ;
        RECT 60.745 138.255 60.915 138.425 ;
        RECT 61.205 138.255 61.375 138.425 ;
        RECT 61.665 138.255 61.835 138.425 ;
        RECT 62.125 138.255 62.295 138.425 ;
        RECT 62.585 138.255 62.755 138.425 ;
        RECT 63.045 138.255 63.215 138.425 ;
        RECT 63.505 138.255 63.675 138.425 ;
        RECT 63.965 138.255 64.135 138.425 ;
        RECT 64.425 138.255 64.595 138.425 ;
        RECT 64.885 138.255 65.055 138.425 ;
        RECT 65.345 138.255 65.515 138.425 ;
        RECT 65.805 138.255 65.975 138.425 ;
        RECT 66.265 138.255 66.435 138.425 ;
        RECT 66.725 138.255 66.895 138.425 ;
        RECT 67.185 138.255 67.355 138.425 ;
        RECT 67.645 138.255 67.815 138.425 ;
        RECT 68.105 138.255 68.275 138.425 ;
        RECT 68.565 138.255 68.735 138.425 ;
        RECT 69.025 138.255 69.195 138.425 ;
        RECT 69.485 138.255 69.655 138.425 ;
        RECT 69.945 138.255 70.115 138.425 ;
        RECT 70.405 138.255 70.575 138.425 ;
        RECT 70.865 138.255 71.035 138.425 ;
        RECT 71.325 138.255 71.495 138.425 ;
        RECT 71.785 138.255 71.955 138.425 ;
        RECT 72.245 138.255 72.415 138.425 ;
        RECT 72.705 138.255 72.875 138.425 ;
        RECT 73.165 138.255 73.335 138.425 ;
        RECT 73.625 138.255 73.795 138.425 ;
        RECT 74.085 138.255 74.255 138.425 ;
        RECT 74.545 138.255 74.715 138.425 ;
        RECT 75.005 138.255 75.175 138.425 ;
        RECT 75.465 138.255 75.635 138.425 ;
        RECT 75.925 138.255 76.095 138.425 ;
        RECT 76.385 138.255 76.555 138.425 ;
        RECT 76.845 138.255 77.015 138.425 ;
        RECT 77.305 138.255 77.475 138.425 ;
        RECT 77.765 138.255 77.935 138.425 ;
        RECT 78.225 138.255 78.395 138.425 ;
        RECT 78.685 138.255 78.855 138.425 ;
        RECT 79.145 138.255 79.315 138.425 ;
        RECT 79.605 138.255 79.775 138.425 ;
        RECT 80.065 138.255 80.235 138.425 ;
        RECT 80.525 138.255 80.695 138.425 ;
        RECT 80.985 138.255 81.155 138.425 ;
        RECT 81.445 138.255 81.615 138.425 ;
        RECT 81.905 138.255 82.075 138.425 ;
        RECT 82.365 138.255 82.535 138.425 ;
        RECT 82.825 138.255 82.995 138.425 ;
        RECT 83.285 138.255 83.455 138.425 ;
        RECT 83.745 138.255 83.915 138.425 ;
        RECT 84.205 138.255 84.375 138.425 ;
        RECT 84.665 138.255 84.835 138.425 ;
        RECT 85.125 138.255 85.295 138.425 ;
        RECT 85.585 138.255 85.755 138.425 ;
        RECT 86.045 138.255 86.215 138.425 ;
        RECT 86.505 138.255 86.675 138.425 ;
        RECT 86.965 138.255 87.135 138.425 ;
        RECT 87.425 138.255 87.595 138.425 ;
        RECT 87.885 138.255 88.055 138.425 ;
        RECT 88.345 138.255 88.515 138.425 ;
        RECT 88.805 138.255 88.975 138.425 ;
        RECT 89.265 138.255 89.435 138.425 ;
        RECT 89.725 138.255 89.895 138.425 ;
        RECT 90.185 138.255 90.355 138.425 ;
        RECT 90.645 138.255 90.815 138.425 ;
        RECT 91.105 138.255 91.275 138.425 ;
        RECT 91.565 138.255 91.735 138.425 ;
        RECT 92.025 138.255 92.195 138.425 ;
        RECT 113.070 136.775 113.260 138.760 ;
        RECT 114.070 136.275 114.260 138.260 ;
        RECT 115.070 136.275 115.260 138.260 ;
        RECT 116.070 136.275 116.260 138.260 ;
        RECT 117.070 136.275 117.260 138.260 ;
        RECT 118.070 136.275 118.260 138.260 ;
        RECT 119.070 136.275 119.260 138.260 ;
        RECT 120.070 136.275 120.260 138.260 ;
        RECT 18.425 135.535 18.595 135.705 ;
        RECT 18.885 135.535 19.055 135.705 ;
        RECT 19.345 135.535 19.515 135.705 ;
        RECT 19.805 135.535 19.975 135.705 ;
        RECT 20.265 135.535 20.435 135.705 ;
        RECT 20.725 135.535 20.895 135.705 ;
        RECT 21.185 135.535 21.355 135.705 ;
        RECT 21.645 135.535 21.815 135.705 ;
        RECT 22.105 135.535 22.275 135.705 ;
        RECT 22.565 135.535 22.735 135.705 ;
        RECT 23.025 135.535 23.195 135.705 ;
        RECT 23.485 135.535 23.655 135.705 ;
        RECT 23.945 135.535 24.115 135.705 ;
        RECT 24.405 135.535 24.575 135.705 ;
        RECT 24.865 135.535 25.035 135.705 ;
        RECT 25.325 135.535 25.495 135.705 ;
        RECT 25.785 135.535 25.955 135.705 ;
        RECT 26.245 135.535 26.415 135.705 ;
        RECT 26.705 135.535 26.875 135.705 ;
        RECT 27.165 135.535 27.335 135.705 ;
        RECT 27.625 135.535 27.795 135.705 ;
        RECT 28.085 135.535 28.255 135.705 ;
        RECT 28.545 135.535 28.715 135.705 ;
        RECT 29.005 135.535 29.175 135.705 ;
        RECT 29.465 135.535 29.635 135.705 ;
        RECT 29.925 135.535 30.095 135.705 ;
        RECT 30.385 135.535 30.555 135.705 ;
        RECT 30.845 135.535 31.015 135.705 ;
        RECT 31.305 135.535 31.475 135.705 ;
        RECT 31.765 135.535 31.935 135.705 ;
        RECT 32.225 135.535 32.395 135.705 ;
        RECT 32.685 135.535 32.855 135.705 ;
        RECT 33.145 135.535 33.315 135.705 ;
        RECT 33.605 135.535 33.775 135.705 ;
        RECT 34.065 135.535 34.235 135.705 ;
        RECT 34.525 135.535 34.695 135.705 ;
        RECT 34.985 135.535 35.155 135.705 ;
        RECT 35.445 135.535 35.615 135.705 ;
        RECT 35.905 135.535 36.075 135.705 ;
        RECT 36.365 135.535 36.535 135.705 ;
        RECT 36.825 135.535 36.995 135.705 ;
        RECT 37.285 135.535 37.455 135.705 ;
        RECT 37.745 135.535 37.915 135.705 ;
        RECT 38.205 135.535 38.375 135.705 ;
        RECT 38.665 135.535 38.835 135.705 ;
        RECT 39.125 135.535 39.295 135.705 ;
        RECT 39.585 135.535 39.755 135.705 ;
        RECT 40.045 135.535 40.215 135.705 ;
        RECT 40.505 135.535 40.675 135.705 ;
        RECT 40.965 135.535 41.135 135.705 ;
        RECT 41.425 135.535 41.595 135.705 ;
        RECT 41.885 135.535 42.055 135.705 ;
        RECT 42.345 135.535 42.515 135.705 ;
        RECT 42.805 135.535 42.975 135.705 ;
        RECT 43.265 135.535 43.435 135.705 ;
        RECT 43.725 135.535 43.895 135.705 ;
        RECT 44.185 135.535 44.355 135.705 ;
        RECT 44.645 135.535 44.815 135.705 ;
        RECT 45.105 135.535 45.275 135.705 ;
        RECT 45.565 135.535 45.735 135.705 ;
        RECT 46.025 135.535 46.195 135.705 ;
        RECT 46.485 135.535 46.655 135.705 ;
        RECT 46.945 135.535 47.115 135.705 ;
        RECT 47.405 135.535 47.575 135.705 ;
        RECT 47.865 135.535 48.035 135.705 ;
        RECT 48.325 135.535 48.495 135.705 ;
        RECT 48.785 135.535 48.955 135.705 ;
        RECT 49.245 135.535 49.415 135.705 ;
        RECT 49.705 135.535 49.875 135.705 ;
        RECT 50.165 135.535 50.335 135.705 ;
        RECT 50.625 135.535 50.795 135.705 ;
        RECT 51.085 135.535 51.255 135.705 ;
        RECT 51.545 135.535 51.715 135.705 ;
        RECT 52.005 135.535 52.175 135.705 ;
        RECT 52.465 135.535 52.635 135.705 ;
        RECT 52.925 135.535 53.095 135.705 ;
        RECT 53.385 135.535 53.555 135.705 ;
        RECT 53.845 135.535 54.015 135.705 ;
        RECT 54.305 135.535 54.475 135.705 ;
        RECT 54.765 135.535 54.935 135.705 ;
        RECT 55.225 135.535 55.395 135.705 ;
        RECT 55.685 135.535 55.855 135.705 ;
        RECT 56.145 135.535 56.315 135.705 ;
        RECT 56.605 135.535 56.775 135.705 ;
        RECT 57.065 135.535 57.235 135.705 ;
        RECT 57.525 135.535 57.695 135.705 ;
        RECT 57.985 135.535 58.155 135.705 ;
        RECT 58.445 135.535 58.615 135.705 ;
        RECT 58.905 135.535 59.075 135.705 ;
        RECT 59.365 135.535 59.535 135.705 ;
        RECT 59.825 135.535 59.995 135.705 ;
        RECT 60.285 135.535 60.455 135.705 ;
        RECT 60.745 135.535 60.915 135.705 ;
        RECT 61.205 135.535 61.375 135.705 ;
        RECT 61.665 135.535 61.835 135.705 ;
        RECT 62.125 135.535 62.295 135.705 ;
        RECT 62.585 135.535 62.755 135.705 ;
        RECT 63.045 135.535 63.215 135.705 ;
        RECT 63.505 135.535 63.675 135.705 ;
        RECT 63.965 135.535 64.135 135.705 ;
        RECT 64.425 135.535 64.595 135.705 ;
        RECT 64.885 135.535 65.055 135.705 ;
        RECT 65.345 135.535 65.515 135.705 ;
        RECT 65.805 135.535 65.975 135.705 ;
        RECT 66.265 135.535 66.435 135.705 ;
        RECT 66.725 135.535 66.895 135.705 ;
        RECT 67.185 135.535 67.355 135.705 ;
        RECT 67.645 135.535 67.815 135.705 ;
        RECT 68.105 135.535 68.275 135.705 ;
        RECT 68.565 135.535 68.735 135.705 ;
        RECT 69.025 135.535 69.195 135.705 ;
        RECT 69.485 135.535 69.655 135.705 ;
        RECT 69.945 135.535 70.115 135.705 ;
        RECT 70.405 135.535 70.575 135.705 ;
        RECT 70.865 135.535 71.035 135.705 ;
        RECT 71.325 135.535 71.495 135.705 ;
        RECT 71.785 135.535 71.955 135.705 ;
        RECT 72.245 135.535 72.415 135.705 ;
        RECT 72.705 135.535 72.875 135.705 ;
        RECT 73.165 135.535 73.335 135.705 ;
        RECT 73.625 135.535 73.795 135.705 ;
        RECT 74.085 135.535 74.255 135.705 ;
        RECT 74.545 135.535 74.715 135.705 ;
        RECT 75.005 135.535 75.175 135.705 ;
        RECT 75.465 135.535 75.635 135.705 ;
        RECT 75.925 135.535 76.095 135.705 ;
        RECT 76.385 135.535 76.555 135.705 ;
        RECT 76.845 135.535 77.015 135.705 ;
        RECT 77.305 135.535 77.475 135.705 ;
        RECT 77.765 135.535 77.935 135.705 ;
        RECT 78.225 135.535 78.395 135.705 ;
        RECT 78.685 135.535 78.855 135.705 ;
        RECT 79.145 135.535 79.315 135.705 ;
        RECT 79.605 135.535 79.775 135.705 ;
        RECT 80.065 135.535 80.235 135.705 ;
        RECT 80.525 135.535 80.695 135.705 ;
        RECT 80.985 135.535 81.155 135.705 ;
        RECT 81.445 135.535 81.615 135.705 ;
        RECT 81.905 135.535 82.075 135.705 ;
        RECT 82.365 135.535 82.535 135.705 ;
        RECT 82.825 135.535 82.995 135.705 ;
        RECT 83.285 135.535 83.455 135.705 ;
        RECT 83.745 135.535 83.915 135.705 ;
        RECT 84.205 135.535 84.375 135.705 ;
        RECT 84.665 135.535 84.835 135.705 ;
        RECT 85.125 135.535 85.295 135.705 ;
        RECT 85.585 135.535 85.755 135.705 ;
        RECT 86.045 135.535 86.215 135.705 ;
        RECT 86.505 135.535 86.675 135.705 ;
        RECT 86.965 135.535 87.135 135.705 ;
        RECT 87.425 135.535 87.595 135.705 ;
        RECT 87.885 135.535 88.055 135.705 ;
        RECT 88.345 135.535 88.515 135.705 ;
        RECT 88.805 135.535 88.975 135.705 ;
        RECT 89.265 135.535 89.435 135.705 ;
        RECT 89.725 135.535 89.895 135.705 ;
        RECT 90.185 135.535 90.355 135.705 ;
        RECT 90.645 135.535 90.815 135.705 ;
        RECT 91.105 135.535 91.275 135.705 ;
        RECT 91.565 135.535 91.735 135.705 ;
        RECT 92.025 135.535 92.195 135.705 ;
        RECT 113.070 133.620 113.260 135.605 ;
        RECT 114.070 133.620 114.260 135.605 ;
        RECT 115.070 133.620 115.260 135.605 ;
        RECT 116.070 133.620 116.260 135.605 ;
        RECT 117.070 133.620 117.260 135.605 ;
        RECT 118.070 133.620 118.260 135.605 ;
        RECT 119.070 133.620 119.260 135.605 ;
        RECT 120.070 133.620 120.260 135.605 ;
        RECT 18.425 132.815 18.595 132.985 ;
        RECT 18.885 132.815 19.055 132.985 ;
        RECT 19.345 132.815 19.515 132.985 ;
        RECT 19.805 132.815 19.975 132.985 ;
        RECT 20.265 132.815 20.435 132.985 ;
        RECT 20.725 132.815 20.895 132.985 ;
        RECT 21.185 132.815 21.355 132.985 ;
        RECT 21.645 132.815 21.815 132.985 ;
        RECT 22.105 132.815 22.275 132.985 ;
        RECT 22.565 132.815 22.735 132.985 ;
        RECT 23.025 132.815 23.195 132.985 ;
        RECT 23.485 132.815 23.655 132.985 ;
        RECT 23.945 132.815 24.115 132.985 ;
        RECT 24.405 132.815 24.575 132.985 ;
        RECT 24.865 132.815 25.035 132.985 ;
        RECT 25.325 132.815 25.495 132.985 ;
        RECT 25.785 132.815 25.955 132.985 ;
        RECT 26.245 132.815 26.415 132.985 ;
        RECT 26.705 132.815 26.875 132.985 ;
        RECT 27.165 132.815 27.335 132.985 ;
        RECT 27.625 132.815 27.795 132.985 ;
        RECT 28.085 132.815 28.255 132.985 ;
        RECT 28.545 132.815 28.715 132.985 ;
        RECT 29.005 132.815 29.175 132.985 ;
        RECT 29.465 132.815 29.635 132.985 ;
        RECT 29.925 132.815 30.095 132.985 ;
        RECT 30.385 132.815 30.555 132.985 ;
        RECT 30.845 132.815 31.015 132.985 ;
        RECT 31.305 132.815 31.475 132.985 ;
        RECT 31.765 132.815 31.935 132.985 ;
        RECT 32.225 132.815 32.395 132.985 ;
        RECT 32.685 132.815 32.855 132.985 ;
        RECT 33.145 132.815 33.315 132.985 ;
        RECT 33.605 132.815 33.775 132.985 ;
        RECT 34.065 132.815 34.235 132.985 ;
        RECT 34.525 132.815 34.695 132.985 ;
        RECT 34.985 132.815 35.155 132.985 ;
        RECT 35.445 132.815 35.615 132.985 ;
        RECT 35.905 132.815 36.075 132.985 ;
        RECT 36.365 132.815 36.535 132.985 ;
        RECT 36.825 132.815 36.995 132.985 ;
        RECT 37.285 132.815 37.455 132.985 ;
        RECT 37.745 132.815 37.915 132.985 ;
        RECT 38.205 132.815 38.375 132.985 ;
        RECT 38.665 132.815 38.835 132.985 ;
        RECT 39.125 132.815 39.295 132.985 ;
        RECT 39.585 132.815 39.755 132.985 ;
        RECT 40.045 132.815 40.215 132.985 ;
        RECT 40.505 132.815 40.675 132.985 ;
        RECT 40.965 132.815 41.135 132.985 ;
        RECT 41.425 132.815 41.595 132.985 ;
        RECT 41.885 132.815 42.055 132.985 ;
        RECT 42.345 132.815 42.515 132.985 ;
        RECT 42.805 132.815 42.975 132.985 ;
        RECT 43.265 132.815 43.435 132.985 ;
        RECT 43.725 132.815 43.895 132.985 ;
        RECT 44.185 132.815 44.355 132.985 ;
        RECT 44.645 132.815 44.815 132.985 ;
        RECT 45.105 132.815 45.275 132.985 ;
        RECT 45.565 132.815 45.735 132.985 ;
        RECT 46.025 132.815 46.195 132.985 ;
        RECT 46.485 132.815 46.655 132.985 ;
        RECT 46.945 132.815 47.115 132.985 ;
        RECT 47.405 132.815 47.575 132.985 ;
        RECT 47.865 132.815 48.035 132.985 ;
        RECT 48.325 132.815 48.495 132.985 ;
        RECT 48.785 132.815 48.955 132.985 ;
        RECT 49.245 132.815 49.415 132.985 ;
        RECT 49.705 132.815 49.875 132.985 ;
        RECT 50.165 132.815 50.335 132.985 ;
        RECT 50.625 132.815 50.795 132.985 ;
        RECT 51.085 132.815 51.255 132.985 ;
        RECT 51.545 132.815 51.715 132.985 ;
        RECT 52.005 132.815 52.175 132.985 ;
        RECT 52.465 132.815 52.635 132.985 ;
        RECT 52.925 132.815 53.095 132.985 ;
        RECT 53.385 132.815 53.555 132.985 ;
        RECT 53.845 132.815 54.015 132.985 ;
        RECT 54.305 132.815 54.475 132.985 ;
        RECT 54.765 132.815 54.935 132.985 ;
        RECT 55.225 132.815 55.395 132.985 ;
        RECT 55.685 132.815 55.855 132.985 ;
        RECT 56.145 132.815 56.315 132.985 ;
        RECT 56.605 132.815 56.775 132.985 ;
        RECT 57.065 132.815 57.235 132.985 ;
        RECT 57.525 132.815 57.695 132.985 ;
        RECT 57.985 132.815 58.155 132.985 ;
        RECT 58.445 132.815 58.615 132.985 ;
        RECT 58.905 132.815 59.075 132.985 ;
        RECT 59.365 132.815 59.535 132.985 ;
        RECT 59.825 132.815 59.995 132.985 ;
        RECT 60.285 132.815 60.455 132.985 ;
        RECT 60.745 132.815 60.915 132.985 ;
        RECT 61.205 132.815 61.375 132.985 ;
        RECT 61.665 132.815 61.835 132.985 ;
        RECT 62.125 132.815 62.295 132.985 ;
        RECT 62.585 132.815 62.755 132.985 ;
        RECT 63.045 132.815 63.215 132.985 ;
        RECT 63.505 132.815 63.675 132.985 ;
        RECT 63.965 132.815 64.135 132.985 ;
        RECT 64.425 132.815 64.595 132.985 ;
        RECT 64.885 132.815 65.055 132.985 ;
        RECT 65.345 132.815 65.515 132.985 ;
        RECT 65.805 132.815 65.975 132.985 ;
        RECT 66.265 132.815 66.435 132.985 ;
        RECT 66.725 132.815 66.895 132.985 ;
        RECT 67.185 132.815 67.355 132.985 ;
        RECT 67.645 132.815 67.815 132.985 ;
        RECT 68.105 132.815 68.275 132.985 ;
        RECT 68.565 132.815 68.735 132.985 ;
        RECT 69.025 132.815 69.195 132.985 ;
        RECT 69.485 132.815 69.655 132.985 ;
        RECT 69.945 132.815 70.115 132.985 ;
        RECT 70.405 132.815 70.575 132.985 ;
        RECT 70.865 132.815 71.035 132.985 ;
        RECT 71.325 132.815 71.495 132.985 ;
        RECT 71.785 132.815 71.955 132.985 ;
        RECT 72.245 132.815 72.415 132.985 ;
        RECT 72.705 132.815 72.875 132.985 ;
        RECT 73.165 132.815 73.335 132.985 ;
        RECT 73.625 132.815 73.795 132.985 ;
        RECT 74.085 132.815 74.255 132.985 ;
        RECT 74.545 132.815 74.715 132.985 ;
        RECT 75.005 132.815 75.175 132.985 ;
        RECT 75.465 132.815 75.635 132.985 ;
        RECT 75.925 132.815 76.095 132.985 ;
        RECT 76.385 132.815 76.555 132.985 ;
        RECT 76.845 132.815 77.015 132.985 ;
        RECT 77.305 132.815 77.475 132.985 ;
        RECT 77.765 132.815 77.935 132.985 ;
        RECT 78.225 132.815 78.395 132.985 ;
        RECT 78.685 132.815 78.855 132.985 ;
        RECT 79.145 132.815 79.315 132.985 ;
        RECT 79.605 132.815 79.775 132.985 ;
        RECT 80.065 132.815 80.235 132.985 ;
        RECT 80.525 132.815 80.695 132.985 ;
        RECT 80.985 132.815 81.155 132.985 ;
        RECT 81.445 132.815 81.615 132.985 ;
        RECT 81.905 132.815 82.075 132.985 ;
        RECT 82.365 132.815 82.535 132.985 ;
        RECT 82.825 132.815 82.995 132.985 ;
        RECT 83.285 132.815 83.455 132.985 ;
        RECT 83.745 132.815 83.915 132.985 ;
        RECT 84.205 132.815 84.375 132.985 ;
        RECT 84.665 132.815 84.835 132.985 ;
        RECT 85.125 132.815 85.295 132.985 ;
        RECT 85.585 132.815 85.755 132.985 ;
        RECT 86.045 132.815 86.215 132.985 ;
        RECT 86.505 132.815 86.675 132.985 ;
        RECT 86.965 132.815 87.135 132.985 ;
        RECT 87.425 132.815 87.595 132.985 ;
        RECT 87.885 132.815 88.055 132.985 ;
        RECT 88.345 132.815 88.515 132.985 ;
        RECT 88.805 132.815 88.975 132.985 ;
        RECT 89.265 132.815 89.435 132.985 ;
        RECT 89.725 132.815 89.895 132.985 ;
        RECT 90.185 132.815 90.355 132.985 ;
        RECT 90.645 132.815 90.815 132.985 ;
        RECT 91.105 132.815 91.275 132.985 ;
        RECT 91.565 132.815 91.735 132.985 ;
        RECT 92.025 132.815 92.195 132.985 ;
      LAYER met1 ;
        RECT 40.430 206.920 40.750 206.980 ;
        RECT 76.310 206.920 76.630 206.980 ;
        RECT 40.430 206.780 76.630 206.920 ;
        RECT 40.430 206.720 40.750 206.780 ;
        RECT 76.310 206.720 76.630 206.780 ;
        RECT 18.280 206.100 92.340 206.580 ;
        RECT 45.950 205.700 46.270 205.960 ;
        RECT 46.870 205.700 47.190 205.960 ;
        RECT 47.790 205.900 48.110 205.960 ;
        RECT 59.305 205.900 59.595 205.945 ;
        RECT 65.285 205.900 65.575 205.945 ;
        RECT 72.630 205.900 72.950 205.960 ;
        RECT 73.105 205.900 73.395 205.945 ;
        RECT 47.790 205.760 73.395 205.900 ;
        RECT 47.790 205.700 48.110 205.760 ;
        RECT 59.305 205.715 59.595 205.760 ;
        RECT 65.285 205.715 65.575 205.760 ;
        RECT 72.630 205.700 72.950 205.760 ;
        RECT 73.105 205.715 73.395 205.760 ;
        RECT 46.960 205.220 47.100 205.700 ;
        RECT 65.730 205.360 66.050 205.620 ;
        RECT 71.250 205.560 71.570 205.620 ;
        RECT 79.530 205.560 79.850 205.620 ;
        RECT 89.665 205.560 89.955 205.605 ;
        RECT 71.250 205.420 75.620 205.560 ;
        RECT 71.250 205.360 71.570 205.420 ;
        RECT 58.845 205.220 59.135 205.265 ;
        RECT 64.825 205.220 65.115 205.265 ;
        RECT 46.960 205.080 48.020 205.220 ;
        RECT 26.170 204.880 26.490 204.940 ;
        RECT 27.565 204.880 27.855 204.925 ;
        RECT 26.170 204.740 27.855 204.880 ;
        RECT 26.170 204.680 26.490 204.740 ;
        RECT 27.565 204.695 27.855 204.740 ;
        RECT 32.610 204.880 32.930 204.940 ;
        RECT 33.545 204.880 33.835 204.925 ;
        RECT 32.610 204.740 33.835 204.880 ;
        RECT 32.610 204.680 32.930 204.740 ;
        RECT 33.545 204.695 33.835 204.740 ;
        RECT 39.050 204.880 39.370 204.940 ;
        RECT 39.985 204.880 40.275 204.925 ;
        RECT 39.050 204.740 40.275 204.880 ;
        RECT 39.050 204.680 39.370 204.740 ;
        RECT 39.985 204.695 40.275 204.740 ;
        RECT 40.905 204.880 41.195 204.925 ;
        RECT 45.490 204.880 45.810 204.940 ;
        RECT 40.905 204.740 45.810 204.880 ;
        RECT 40.905 204.695 41.195 204.740 ;
        RECT 45.490 204.680 45.810 204.740 ;
        RECT 45.965 204.880 46.255 204.925 ;
        RECT 46.870 204.880 47.190 204.940 ;
        RECT 45.965 204.740 47.190 204.880 ;
        RECT 45.965 204.695 46.255 204.740 ;
        RECT 46.870 204.680 47.190 204.740 ;
        RECT 47.330 204.680 47.650 204.940 ;
        RECT 47.880 204.925 48.020 205.080 ;
        RECT 58.000 205.080 65.115 205.220 ;
        RECT 65.820 205.220 65.960 205.360 ;
        RECT 73.565 205.220 73.855 205.265 ;
        RECT 65.820 205.080 66.880 205.220 ;
        RECT 47.805 204.695 48.095 204.925 ;
        RECT 51.930 204.880 52.250 204.940 ;
        RECT 52.405 204.880 52.695 204.925 ;
        RECT 51.930 204.740 52.695 204.880 ;
        RECT 51.930 204.680 52.250 204.740 ;
        RECT 52.405 204.695 52.695 204.740 ;
        RECT 57.450 204.680 57.770 204.940 ;
        RECT 34.465 204.540 34.755 204.585 ;
        RECT 40.430 204.540 40.750 204.600 ;
        RECT 45.580 204.540 45.720 204.680 ;
        RECT 58.000 204.600 58.140 205.080 ;
        RECT 58.845 205.035 59.135 205.080 ;
        RECT 64.825 205.035 65.115 205.080 ;
        RECT 58.370 204.680 58.690 204.940 ;
        RECT 61.605 204.695 61.895 204.925 ;
        RECT 57.910 204.540 58.230 204.600 ;
        RECT 34.465 204.400 40.750 204.540 ;
        RECT 34.465 204.355 34.755 204.400 ;
        RECT 40.430 204.340 40.750 204.400 ;
        RECT 44.200 204.400 45.260 204.540 ;
        RECT 45.580 204.400 58.230 204.540 ;
        RECT 58.460 204.540 58.600 204.680 ;
        RECT 61.680 204.540 61.820 204.695 ;
        RECT 58.460 204.400 61.820 204.540 ;
        RECT 64.900 204.540 65.040 205.035 ;
        RECT 66.190 204.680 66.510 204.940 ;
        RECT 66.740 204.925 66.880 205.080 ;
        RECT 67.200 205.080 73.855 205.220 ;
        RECT 66.665 204.695 66.955 204.925 ;
        RECT 67.200 204.540 67.340 205.080 ;
        RECT 73.565 205.035 73.855 205.080 ;
        RECT 75.480 204.925 75.620 205.420 ;
        RECT 79.530 205.420 89.955 205.560 ;
        RECT 79.530 205.360 79.850 205.420 ;
        RECT 89.665 205.375 89.955 205.420 ;
        RECT 74.945 204.695 75.235 204.925 ;
        RECT 75.405 204.695 75.695 204.925 ;
        RECT 77.690 204.880 78.010 204.940 ;
        RECT 78.165 204.880 78.455 204.925 ;
        RECT 77.690 204.740 78.455 204.880 ;
        RECT 64.900 204.400 67.340 204.540 ;
        RECT 75.020 204.540 75.160 204.695 ;
        RECT 77.690 204.680 78.010 204.740 ;
        RECT 78.165 204.695 78.455 204.740 ;
        RECT 81.370 204.680 81.690 204.940 ;
        RECT 82.305 204.695 82.595 204.925 ;
        RECT 84.130 204.880 84.450 204.940 ;
        RECT 84.605 204.880 84.895 204.925 ;
        RECT 84.130 204.740 84.895 204.880 ;
        RECT 82.380 204.540 82.520 204.695 ;
        RECT 84.130 204.680 84.450 204.740 ;
        RECT 84.605 204.695 84.895 204.740 ;
        RECT 90.570 204.680 90.890 204.940 ;
        RECT 75.020 204.400 75.620 204.540 ;
        RECT 82.380 204.400 84.820 204.540 ;
        RECT 44.200 204.260 44.340 204.400 ;
        RECT 26.170 204.000 26.490 204.260 ;
        RECT 28.470 204.000 28.790 204.260 ;
        RECT 44.110 204.000 44.430 204.260 ;
        RECT 44.570 204.000 44.890 204.260 ;
        RECT 45.120 204.200 45.260 204.400 ;
        RECT 57.910 204.340 58.230 204.400 ;
        RECT 75.480 204.260 75.620 204.400 ;
        RECT 84.680 204.260 84.820 204.400 ;
        RECT 48.725 204.200 49.015 204.245 ;
        RECT 45.120 204.060 49.015 204.200 ;
        RECT 48.725 204.015 49.015 204.060 ;
        RECT 53.310 204.000 53.630 204.260 ;
        RECT 60.210 204.000 60.530 204.260 ;
        RECT 60.670 204.000 60.990 204.260 ;
        RECT 62.970 204.200 63.290 204.260 ;
        RECT 63.445 204.200 63.735 204.245 ;
        RECT 62.970 204.060 63.735 204.200 ;
        RECT 62.970 204.000 63.290 204.060 ;
        RECT 63.445 204.015 63.735 204.060 ;
        RECT 67.570 204.000 67.890 204.260 ;
        RECT 72.170 204.000 72.490 204.260 ;
        RECT 75.390 204.000 75.710 204.260 ;
        RECT 76.325 204.200 76.615 204.245 ;
        RECT 76.770 204.200 77.090 204.260 ;
        RECT 76.325 204.060 77.090 204.200 ;
        RECT 76.325 204.015 76.615 204.060 ;
        RECT 76.770 204.000 77.090 204.060 ;
        RECT 79.070 204.000 79.390 204.260 ;
        RECT 81.830 204.000 82.150 204.260 ;
        RECT 84.590 204.000 84.910 204.260 ;
        RECT 85.525 204.200 85.815 204.245 ;
        RECT 86.430 204.200 86.750 204.260 ;
        RECT 85.525 204.060 86.750 204.200 ;
        RECT 85.525 204.015 85.815 204.060 ;
        RECT 86.430 204.000 86.750 204.060 ;
        RECT 18.280 203.380 93.120 203.860 ;
        RECT 26.170 202.980 26.490 203.240 ;
        RECT 33.085 202.995 33.375 203.225 ;
        RECT 44.570 203.180 44.890 203.240 ;
        RECT 45.045 203.180 45.335 203.225 ;
        RECT 44.570 203.040 45.335 203.180 ;
        RECT 25.725 202.840 26.015 202.885 ;
        RECT 26.260 202.840 26.400 202.980 ;
        RECT 25.725 202.700 26.400 202.840 ;
        RECT 28.005 202.840 28.655 202.885 ;
        RECT 28.930 202.840 29.250 202.900 ;
        RECT 31.605 202.840 31.895 202.885 ;
        RECT 28.005 202.700 31.895 202.840 ;
        RECT 33.160 202.840 33.300 202.995 ;
        RECT 44.570 202.980 44.890 203.040 ;
        RECT 45.045 202.995 45.335 203.040 ;
        RECT 50.565 203.180 50.855 203.225 ;
        RECT 52.390 203.180 52.710 203.240 ;
        RECT 57.450 203.180 57.770 203.240 ;
        RECT 50.565 203.040 57.770 203.180 ;
        RECT 50.565 202.995 50.855 203.040 ;
        RECT 52.390 202.980 52.710 203.040 ;
        RECT 57.450 202.980 57.770 203.040 ;
        RECT 60.225 203.180 60.515 203.225 ;
        RECT 62.510 203.180 62.830 203.240 ;
        RECT 66.190 203.180 66.510 203.240 ;
        RECT 60.225 203.040 66.510 203.180 ;
        RECT 60.225 202.995 60.515 203.040 ;
        RECT 62.510 202.980 62.830 203.040 ;
        RECT 66.190 202.980 66.510 203.040 ;
        RECT 70.345 203.180 70.635 203.225 ;
        RECT 75.390 203.180 75.710 203.240 ;
        RECT 70.345 203.040 75.710 203.180 ;
        RECT 70.345 202.995 70.635 203.040 ;
        RECT 75.390 202.980 75.710 203.040 ;
        RECT 81.370 203.180 81.690 203.240 ;
        RECT 81.845 203.180 82.135 203.225 ;
        RECT 81.370 203.040 82.135 203.180 ;
        RECT 81.370 202.980 81.690 203.040 ;
        RECT 81.845 202.995 82.135 203.040 ;
        RECT 34.465 202.840 34.755 202.885 ;
        RECT 47.790 202.840 48.110 202.900 ;
        RECT 83.230 202.840 83.520 202.885 ;
        RECT 84.630 202.840 84.920 202.885 ;
        RECT 86.470 202.840 86.760 202.885 ;
        RECT 33.160 202.700 48.110 202.840 ;
        RECT 25.725 202.655 26.015 202.700 ;
        RECT 28.005 202.655 28.655 202.700 ;
        RECT 28.930 202.640 29.250 202.700 ;
        RECT 31.305 202.655 31.895 202.700 ;
        RECT 34.465 202.655 34.755 202.700 ;
        RECT 24.810 202.500 25.100 202.545 ;
        RECT 26.645 202.500 26.935 202.545 ;
        RECT 30.225 202.500 30.515 202.545 ;
        RECT 24.810 202.360 30.515 202.500 ;
        RECT 24.810 202.315 25.100 202.360 ;
        RECT 26.645 202.315 26.935 202.360 ;
        RECT 30.225 202.315 30.515 202.360 ;
        RECT 31.305 202.340 31.595 202.655 ;
        RECT 47.790 202.640 48.110 202.700 ;
        RECT 57.540 202.700 82.520 202.840 ;
        RECT 38.100 202.500 38.390 202.545 ;
        RECT 43.190 202.500 43.510 202.560 ;
        RECT 38.100 202.360 43.510 202.500 ;
        RECT 38.100 202.315 38.390 202.360 ;
        RECT 43.190 202.300 43.510 202.360 ;
        RECT 45.490 202.500 45.810 202.560 ;
        RECT 48.725 202.500 49.015 202.545 ;
        RECT 53.310 202.500 53.630 202.560 ;
        RECT 45.490 202.360 49.015 202.500 ;
        RECT 45.490 202.300 45.810 202.360 ;
        RECT 48.725 202.315 49.015 202.360 ;
        RECT 52.480 202.360 53.630 202.500 ;
        RECT 24.345 202.160 24.635 202.205 ;
        RECT 32.150 202.160 32.470 202.220 ;
        RECT 36.765 202.160 37.055 202.205 ;
        RECT 24.345 202.020 37.055 202.160 ;
        RECT 24.345 201.975 24.635 202.020 ;
        RECT 32.150 201.960 32.470 202.020 ;
        RECT 36.765 201.975 37.055 202.020 ;
        RECT 37.645 202.160 37.935 202.205 ;
        RECT 38.835 202.160 39.125 202.205 ;
        RECT 41.355 202.160 41.645 202.205 ;
        RECT 37.645 202.020 41.645 202.160 ;
        RECT 37.645 201.975 37.935 202.020 ;
        RECT 38.835 201.975 39.125 202.020 ;
        RECT 41.355 201.975 41.645 202.020 ;
        RECT 46.870 201.960 47.190 202.220 ;
        RECT 47.345 202.160 47.635 202.205 ;
        RECT 52.480 202.160 52.620 202.360 ;
        RECT 53.310 202.300 53.630 202.360 ;
        RECT 56.185 202.500 56.475 202.545 ;
        RECT 56.990 202.500 57.310 202.560 ;
        RECT 57.540 202.545 57.680 202.700 ;
        RECT 67.200 202.560 67.340 202.700 ;
        RECT 56.185 202.360 57.310 202.500 ;
        RECT 56.185 202.315 56.475 202.360 ;
        RECT 56.990 202.300 57.310 202.360 ;
        RECT 57.465 202.315 57.755 202.545 ;
        RECT 65.845 202.500 66.135 202.545 ;
        RECT 66.650 202.500 66.970 202.560 ;
        RECT 65.845 202.360 66.970 202.500 ;
        RECT 65.845 202.315 66.135 202.360 ;
        RECT 66.650 202.300 66.970 202.360 ;
        RECT 67.110 202.300 67.430 202.560 ;
        RECT 75.850 202.545 76.170 202.560 ;
        RECT 77.320 202.545 77.460 202.700 ;
        RECT 79.530 202.545 79.850 202.560 ;
        RECT 75.850 202.315 76.200 202.545 ;
        RECT 77.245 202.315 77.535 202.545 ;
        RECT 79.415 202.315 79.850 202.545 ;
        RECT 75.850 202.300 76.170 202.315 ;
        RECT 79.530 202.300 79.850 202.315 ;
        RECT 79.990 202.300 80.310 202.560 ;
        RECT 80.450 202.300 80.770 202.560 ;
        RECT 80.910 202.300 81.230 202.560 ;
        RECT 82.380 202.545 82.520 202.700 ;
        RECT 83.230 202.700 86.760 202.840 ;
        RECT 83.230 202.655 83.520 202.700 ;
        RECT 84.630 202.655 84.920 202.700 ;
        RECT 86.470 202.655 86.760 202.700 ;
        RECT 82.305 202.315 82.595 202.545 ;
        RECT 90.570 202.300 90.890 202.560 ;
        RECT 47.345 202.020 52.620 202.160 ;
        RECT 52.875 202.160 53.165 202.205 ;
        RECT 55.395 202.160 55.685 202.205 ;
        RECT 56.585 202.160 56.875 202.205 ;
        RECT 52.875 202.020 56.875 202.160 ;
        RECT 47.345 201.975 47.635 202.020 ;
        RECT 52.875 201.975 53.165 202.020 ;
        RECT 55.395 201.975 55.685 202.020 ;
        RECT 56.585 201.975 56.875 202.020 ;
        RECT 62.535 202.160 62.825 202.205 ;
        RECT 65.055 202.160 65.345 202.205 ;
        RECT 66.245 202.160 66.535 202.205 ;
        RECT 62.535 202.020 66.535 202.160 ;
        RECT 62.535 201.975 62.825 202.020 ;
        RECT 65.055 201.975 65.345 202.020 ;
        RECT 66.245 201.975 66.535 202.020 ;
        RECT 72.655 202.160 72.945 202.205 ;
        RECT 75.175 202.160 75.465 202.205 ;
        RECT 76.365 202.160 76.655 202.205 ;
        RECT 72.655 202.020 76.655 202.160 ;
        RECT 72.655 201.975 72.945 202.020 ;
        RECT 75.175 201.975 75.465 202.020 ;
        RECT 76.365 201.975 76.655 202.020 ;
        RECT 78.625 201.975 78.915 202.205 ;
        RECT 83.685 202.160 83.975 202.205 ;
        RECT 84.130 202.160 84.450 202.220 ;
        RECT 83.685 202.020 84.450 202.160 ;
        RECT 83.685 201.975 83.975 202.020 ;
        RECT 25.215 201.820 25.505 201.865 ;
        RECT 27.105 201.820 27.395 201.865 ;
        RECT 30.225 201.820 30.515 201.865 ;
        RECT 34.910 201.820 35.230 201.880 ;
        RECT 35.385 201.820 35.675 201.865 ;
        RECT 25.215 201.680 30.515 201.820 ;
        RECT 25.215 201.635 25.505 201.680 ;
        RECT 27.105 201.635 27.395 201.680 ;
        RECT 30.225 201.635 30.515 201.680 ;
        RECT 31.320 201.680 35.675 201.820 ;
        RECT 31.320 201.540 31.460 201.680 ;
        RECT 34.910 201.620 35.230 201.680 ;
        RECT 35.385 201.635 35.675 201.680 ;
        RECT 37.250 201.820 37.540 201.865 ;
        RECT 39.350 201.820 39.640 201.865 ;
        RECT 40.920 201.820 41.210 201.865 ;
        RECT 37.250 201.680 41.210 201.820 ;
        RECT 46.960 201.820 47.100 201.960 ;
        RECT 53.310 201.820 53.600 201.865 ;
        RECT 54.880 201.820 55.170 201.865 ;
        RECT 56.980 201.820 57.270 201.865 ;
        RECT 46.960 201.680 49.860 201.820 ;
        RECT 37.250 201.635 37.540 201.680 ;
        RECT 39.350 201.635 39.640 201.680 ;
        RECT 40.920 201.635 41.210 201.680 ;
        RECT 31.230 201.280 31.550 201.540 ;
        RECT 43.665 201.480 43.955 201.525 ;
        RECT 44.570 201.480 44.890 201.540 ;
        RECT 43.665 201.340 44.890 201.480 ;
        RECT 43.665 201.295 43.955 201.340 ;
        RECT 44.570 201.280 44.890 201.340 ;
        RECT 45.950 201.480 46.270 201.540 ;
        RECT 46.870 201.480 47.190 201.540 ;
        RECT 45.950 201.340 47.190 201.480 ;
        RECT 45.950 201.280 46.270 201.340 ;
        RECT 46.870 201.280 47.190 201.340 ;
        RECT 48.250 201.280 48.570 201.540 ;
        RECT 49.720 201.525 49.860 201.680 ;
        RECT 53.310 201.680 57.270 201.820 ;
        RECT 53.310 201.635 53.600 201.680 ;
        RECT 54.880 201.635 55.170 201.680 ;
        RECT 56.980 201.635 57.270 201.680 ;
        RECT 62.970 201.820 63.260 201.865 ;
        RECT 64.540 201.820 64.830 201.865 ;
        RECT 66.640 201.820 66.930 201.865 ;
        RECT 62.970 201.680 66.930 201.820 ;
        RECT 62.970 201.635 63.260 201.680 ;
        RECT 64.540 201.635 64.830 201.680 ;
        RECT 66.640 201.635 66.930 201.680 ;
        RECT 73.090 201.820 73.380 201.865 ;
        RECT 74.660 201.820 74.950 201.865 ;
        RECT 76.760 201.820 77.050 201.865 ;
        RECT 73.090 201.680 77.050 201.820 ;
        RECT 73.090 201.635 73.380 201.680 ;
        RECT 74.660 201.635 74.950 201.680 ;
        RECT 76.760 201.635 77.050 201.680 ;
        RECT 49.645 201.480 49.935 201.525 ;
        RECT 50.090 201.480 50.410 201.540 ;
        RECT 49.645 201.340 50.410 201.480 ;
        RECT 49.645 201.295 49.935 201.340 ;
        RECT 50.090 201.280 50.410 201.340 ;
        RECT 77.690 201.480 78.010 201.540 ;
        RECT 78.700 201.480 78.840 201.975 ;
        RECT 84.130 201.960 84.450 202.020 ;
        RECT 82.770 201.820 83.060 201.865 ;
        RECT 85.090 201.820 85.380 201.865 ;
        RECT 86.470 201.820 86.760 201.865 ;
        RECT 82.770 201.680 86.760 201.820 ;
        RECT 82.770 201.635 83.060 201.680 ;
        RECT 85.090 201.635 85.380 201.680 ;
        RECT 86.470 201.635 86.760 201.680 ;
        RECT 85.510 201.480 85.830 201.540 ;
        RECT 77.690 201.340 85.830 201.480 ;
        RECT 77.690 201.280 78.010 201.340 ;
        RECT 85.510 201.280 85.830 201.340 ;
        RECT 18.280 200.660 92.340 201.140 ;
        RECT 28.470 200.260 28.790 200.520 ;
        RECT 28.930 200.260 29.250 200.520 ;
        RECT 34.910 200.460 35.230 200.520 ;
        RECT 46.870 200.460 47.190 200.520 ;
        RECT 49.185 200.460 49.475 200.505 ;
        RECT 34.910 200.320 49.475 200.460 ;
        RECT 34.910 200.260 35.230 200.320 ;
        RECT 46.870 200.260 47.190 200.320 ;
        RECT 49.185 200.275 49.475 200.320 ;
        RECT 56.990 200.460 57.310 200.520 ;
        RECT 57.465 200.460 57.755 200.505 ;
        RECT 56.990 200.320 57.755 200.460 ;
        RECT 28.560 199.440 28.700 200.260 ;
        RECT 29.020 199.780 29.160 200.260 ;
        RECT 33.570 200.120 33.860 200.165 ;
        RECT 35.670 200.120 35.960 200.165 ;
        RECT 37.240 200.120 37.530 200.165 ;
        RECT 33.570 199.980 37.530 200.120 ;
        RECT 33.570 199.935 33.860 199.980 ;
        RECT 35.670 199.935 35.960 199.980 ;
        RECT 37.240 199.935 37.530 199.980 ;
        RECT 39.985 200.120 40.275 200.165 ;
        RECT 43.650 200.120 43.970 200.180 ;
        RECT 47.330 200.120 47.650 200.180 ;
        RECT 39.985 199.980 47.650 200.120 ;
        RECT 39.985 199.935 40.275 199.980 ;
        RECT 43.650 199.920 43.970 199.980 ;
        RECT 47.330 199.920 47.650 199.980 ;
        RECT 48.250 199.920 48.570 200.180 ;
        RECT 49.260 200.120 49.400 200.275 ;
        RECT 56.990 200.260 57.310 200.320 ;
        RECT 57.465 200.275 57.755 200.320 ;
        RECT 58.370 200.260 58.690 200.520 ;
        RECT 66.650 200.260 66.970 200.520 ;
        RECT 75.405 200.460 75.695 200.505 ;
        RECT 75.850 200.460 76.170 200.520 ;
        RECT 75.405 200.320 76.170 200.460 ;
        RECT 75.405 200.275 75.695 200.320 ;
        RECT 75.850 200.260 76.170 200.320 ;
        RECT 80.910 200.460 81.230 200.520 ;
        RECT 81.385 200.460 81.675 200.505 ;
        RECT 80.910 200.320 81.675 200.460 ;
        RECT 80.910 200.260 81.230 200.320 ;
        RECT 81.385 200.275 81.675 200.320 ;
        RECT 83.225 200.460 83.515 200.505 ;
        RECT 84.130 200.460 84.450 200.520 ;
        RECT 83.225 200.320 84.450 200.460 ;
        RECT 83.225 200.275 83.515 200.320 ;
        RECT 84.130 200.260 84.450 200.320 ;
        RECT 58.460 200.120 58.600 200.260 ;
        RECT 76.770 200.120 77.090 200.180 ;
        RECT 49.260 199.980 58.600 200.120 ;
        RECT 65.820 199.980 77.090 200.120 ;
        RECT 33.965 199.780 34.255 199.825 ;
        RECT 35.155 199.780 35.445 199.825 ;
        RECT 37.675 199.780 37.965 199.825 ;
        RECT 48.340 199.780 48.480 199.920 ;
        RECT 50.090 199.780 50.410 199.840 ;
        RECT 60.210 199.780 60.530 199.840 ;
        RECT 60.685 199.780 60.975 199.825 ;
        RECT 29.020 199.640 29.620 199.780 ;
        RECT 28.945 199.440 29.235 199.485 ;
        RECT 28.560 199.300 29.235 199.440 ;
        RECT 28.945 199.255 29.235 199.300 ;
        RECT 28.485 199.100 28.775 199.145 ;
        RECT 29.480 199.100 29.620 199.640 ;
        RECT 33.965 199.640 37.965 199.780 ;
        RECT 33.965 199.595 34.255 199.640 ;
        RECT 35.155 199.595 35.445 199.640 ;
        RECT 37.675 199.595 37.965 199.640 ;
        RECT 41.440 199.640 48.480 199.780 ;
        RECT 49.260 199.640 59.060 199.780 ;
        RECT 32.150 199.440 32.470 199.500 ;
        RECT 33.085 199.440 33.375 199.485 ;
        RECT 32.150 199.300 33.375 199.440 ;
        RECT 32.150 199.240 32.470 199.300 ;
        RECT 33.085 199.255 33.375 199.300 ;
        RECT 34.420 199.440 34.710 199.485 ;
        RECT 41.440 199.440 41.580 199.640 ;
        RECT 34.420 199.300 41.580 199.440 ;
        RECT 34.420 199.255 34.710 199.300 ;
        RECT 43.190 199.240 43.510 199.500 ;
        RECT 44.110 199.240 44.430 199.500 ;
        RECT 44.585 199.440 44.875 199.485 ;
        RECT 48.265 199.440 48.555 199.485 ;
        RECT 49.260 199.440 49.400 199.640 ;
        RECT 50.090 199.580 50.410 199.640 ;
        RECT 58.920 199.500 59.060 199.640 ;
        RECT 60.210 199.640 60.975 199.780 ;
        RECT 60.210 199.580 60.530 199.640 ;
        RECT 60.685 199.595 60.975 199.640 ;
        RECT 62.970 199.780 63.290 199.840 ;
        RECT 65.820 199.825 65.960 199.980 ;
        RECT 76.770 199.920 77.090 199.980 ;
        RECT 63.445 199.780 63.735 199.825 ;
        RECT 62.970 199.640 63.735 199.780 ;
        RECT 62.970 199.580 63.290 199.640 ;
        RECT 63.445 199.595 63.735 199.640 ;
        RECT 65.745 199.595 66.035 199.825 ;
        RECT 72.170 199.580 72.490 199.840 ;
        RECT 74.025 199.780 74.315 199.825 ;
        RECT 79.530 199.780 79.850 199.840 ;
        RECT 89.205 199.780 89.495 199.825 ;
        RECT 90.570 199.780 90.890 199.840 ;
        RECT 74.025 199.640 79.850 199.780 ;
        RECT 74.025 199.595 74.315 199.640 ;
        RECT 79.530 199.580 79.850 199.640 ;
        RECT 81.460 199.640 90.890 199.780 ;
        RECT 44.585 199.300 49.400 199.440 ;
        RECT 44.585 199.255 44.875 199.300 ;
        RECT 48.265 199.255 48.555 199.300 ;
        RECT 49.645 199.255 49.935 199.485 ;
        RECT 58.385 199.255 58.675 199.485 ;
        RECT 58.830 199.440 59.150 199.500 ;
        RECT 65.270 199.440 65.590 199.500 ;
        RECT 58.830 199.300 65.590 199.440 ;
        RECT 49.720 199.100 49.860 199.255 ;
        RECT 28.485 198.960 29.620 199.100 ;
        RECT 44.660 198.960 49.860 199.100 ;
        RECT 58.460 199.100 58.600 199.255 ;
        RECT 58.830 199.240 59.150 199.300 ;
        RECT 65.270 199.240 65.590 199.300 ;
        RECT 67.570 199.240 67.890 199.500 ;
        RECT 74.485 199.440 74.775 199.485 ;
        RECT 74.930 199.440 75.250 199.500 ;
        RECT 74.485 199.300 75.250 199.440 ;
        RECT 74.485 199.255 74.775 199.300 ;
        RECT 74.930 199.240 75.250 199.300 ;
        RECT 76.310 199.440 76.630 199.500 ;
        RECT 81.460 199.485 81.600 199.640 ;
        RECT 89.205 199.595 89.495 199.640 ;
        RECT 90.570 199.580 90.890 199.640 ;
        RECT 80.465 199.440 80.755 199.485 ;
        RECT 76.310 199.300 80.755 199.440 ;
        RECT 76.310 199.240 76.630 199.300 ;
        RECT 80.465 199.255 80.755 199.300 ;
        RECT 81.385 199.255 81.675 199.485 ;
        RECT 81.830 199.440 82.150 199.500 ;
        RECT 84.145 199.440 84.435 199.485 ;
        RECT 81.830 199.300 84.435 199.440 ;
        RECT 81.830 199.240 82.150 199.300 ;
        RECT 84.145 199.255 84.435 199.300 ;
        RECT 84.590 199.240 84.910 199.500 ;
        RECT 67.660 199.100 67.800 199.240 ;
        RECT 83.225 199.100 83.515 199.145 ;
        RECT 58.460 198.960 67.800 199.100 ;
        RECT 81.920 198.960 83.515 199.100 ;
        RECT 28.485 198.915 28.775 198.960 ;
        RECT 44.660 198.820 44.800 198.960 ;
        RECT 81.920 198.820 82.060 198.960 ;
        RECT 83.225 198.915 83.515 198.960 ;
        RECT 44.570 198.560 44.890 198.820 ;
        RECT 46.425 198.760 46.715 198.805 ;
        RECT 46.885 198.760 47.175 198.805 ;
        RECT 46.425 198.620 47.175 198.760 ;
        RECT 46.425 198.575 46.715 198.620 ;
        RECT 46.885 198.575 47.175 198.620 ;
        RECT 53.310 198.760 53.630 198.820 ;
        RECT 68.030 198.760 68.350 198.820 ;
        RECT 53.310 198.620 68.350 198.760 ;
        RECT 53.310 198.560 53.630 198.620 ;
        RECT 68.030 198.560 68.350 198.620 ;
        RECT 81.830 198.560 82.150 198.820 ;
        RECT 82.290 198.760 82.610 198.820 ;
        RECT 85.985 198.760 86.275 198.805 ;
        RECT 82.290 198.620 86.275 198.760 ;
        RECT 82.290 198.560 82.610 198.620 ;
        RECT 85.985 198.575 86.275 198.620 ;
        RECT 18.280 197.940 93.120 198.420 ;
        RECT 56.545 197.740 56.835 197.785 ;
        RECT 57.005 197.740 57.295 197.785 ;
        RECT 79.070 197.740 79.390 197.800 ;
        RECT 56.545 197.600 57.295 197.740 ;
        RECT 56.545 197.555 56.835 197.600 ;
        RECT 57.005 197.555 57.295 197.600 ;
        RECT 64.900 197.600 79.390 197.740 ;
        RECT 47.790 196.860 48.110 197.120 ;
        RECT 54.705 197.060 54.995 197.105 ;
        RECT 58.830 197.060 59.150 197.120 ;
        RECT 54.705 196.920 59.150 197.060 ;
        RECT 54.705 196.875 54.995 196.920 ;
        RECT 58.830 196.860 59.150 196.920 ;
        RECT 59.750 196.860 60.070 197.120 ;
        RECT 64.900 197.105 65.040 197.600 ;
        RECT 79.070 197.540 79.390 197.600 ;
        RECT 81.385 197.740 81.675 197.785 ;
        RECT 84.590 197.740 84.910 197.800 ;
        RECT 81.385 197.600 84.910 197.740 ;
        RECT 81.385 197.555 81.675 197.600 ;
        RECT 84.590 197.540 84.910 197.600 ;
        RECT 84.130 197.400 84.450 197.460 ;
        RECT 83.300 197.260 84.450 197.400 ;
        RECT 64.825 196.875 65.115 197.105 ;
        RECT 65.270 197.060 65.590 197.120 ;
        RECT 73.565 197.060 73.855 197.105 ;
        RECT 74.930 197.060 75.250 197.120 ;
        RECT 65.270 196.920 75.250 197.060 ;
        RECT 65.270 196.860 65.590 196.920 ;
        RECT 73.565 196.875 73.855 196.920 ;
        RECT 74.930 196.860 75.250 196.920 ;
        RECT 78.610 197.060 78.930 197.120 ;
        RECT 83.300 197.105 83.440 197.260 ;
        RECT 84.130 197.200 84.450 197.260 ;
        RECT 85.140 197.260 88.040 197.400 ;
        RECT 80.005 197.060 80.295 197.105 ;
        RECT 81.845 197.060 82.135 197.105 ;
        RECT 78.610 196.920 80.295 197.060 ;
        RECT 78.610 196.860 78.930 196.920 ;
        RECT 80.005 196.875 80.295 196.920 ;
        RECT 80.540 196.920 82.135 197.060 ;
        RECT 54.245 196.535 54.535 196.765 ;
        RECT 57.910 196.720 58.230 196.780 ;
        RECT 58.385 196.720 58.675 196.765 ;
        RECT 57.910 196.580 58.675 196.720 ;
        RECT 54.320 196.380 54.460 196.535 ;
        RECT 57.910 196.520 58.230 196.580 ;
        RECT 58.385 196.535 58.675 196.580 ;
        RECT 66.190 196.720 66.510 196.780 ;
        RECT 67.125 196.720 67.415 196.765 ;
        RECT 66.190 196.580 67.415 196.720 ;
        RECT 66.190 196.520 66.510 196.580 ;
        RECT 67.125 196.535 67.415 196.580 ;
        RECT 71.710 196.520 72.030 196.780 ;
        RECT 74.025 196.535 74.315 196.765 ;
        RECT 77.230 196.720 77.550 196.780 ;
        RECT 80.540 196.720 80.680 196.920 ;
        RECT 81.845 196.875 82.135 196.920 ;
        RECT 82.765 196.875 83.055 197.105 ;
        RECT 83.225 196.875 83.515 197.105 ;
        RECT 83.685 197.060 83.975 197.105 ;
        RECT 85.140 197.060 85.280 197.260 ;
        RECT 87.900 197.120 88.040 197.260 ;
        RECT 83.685 196.920 85.280 197.060 ;
        RECT 83.685 196.875 83.975 196.920 ;
        RECT 77.230 196.580 80.680 196.720 ;
        RECT 81.385 196.720 81.675 196.765 ;
        RECT 82.290 196.720 82.610 196.780 ;
        RECT 81.385 196.580 82.610 196.720 ;
        RECT 82.840 196.720 82.980 196.875 ;
        RECT 85.510 196.860 85.830 197.120 ;
        RECT 86.430 196.860 86.750 197.120 ;
        RECT 87.810 196.860 88.130 197.120 ;
        RECT 84.130 196.720 84.450 196.780 ;
        RECT 82.840 196.580 84.450 196.720 ;
        RECT 60.670 196.380 60.990 196.440 ;
        RECT 54.320 196.240 60.990 196.380 ;
        RECT 74.100 196.380 74.240 196.535 ;
        RECT 77.230 196.520 77.550 196.580 ;
        RECT 81.385 196.535 81.675 196.580 ;
        RECT 82.290 196.520 82.610 196.580 ;
        RECT 84.130 196.520 84.450 196.580 ;
        RECT 86.520 196.380 86.660 196.860 ;
        RECT 74.100 196.240 86.660 196.380 ;
        RECT 58.460 196.100 58.600 196.240 ;
        RECT 60.670 196.180 60.990 196.240 ;
        RECT 47.790 196.040 48.110 196.100 ;
        RECT 48.265 196.040 48.555 196.085 ;
        RECT 47.790 195.900 48.555 196.040 ;
        RECT 47.790 195.840 48.110 195.900 ;
        RECT 48.265 195.855 48.555 195.900 ;
        RECT 53.325 196.040 53.615 196.085 ;
        RECT 53.770 196.040 54.090 196.100 ;
        RECT 53.325 195.900 54.090 196.040 ;
        RECT 53.325 195.855 53.615 195.900 ;
        RECT 53.770 195.840 54.090 195.900 ;
        RECT 58.370 195.840 58.690 196.100 ;
        RECT 58.830 196.040 59.150 196.100 ;
        RECT 59.305 196.040 59.595 196.085 ;
        RECT 62.970 196.040 63.290 196.100 ;
        RECT 58.830 195.900 63.290 196.040 ;
        RECT 58.830 195.840 59.150 195.900 ;
        RECT 59.305 195.855 59.595 195.900 ;
        RECT 62.970 195.840 63.290 195.900 ;
        RECT 63.905 196.040 64.195 196.085 ;
        RECT 65.730 196.040 66.050 196.100 ;
        RECT 63.905 195.900 66.050 196.040 ;
        RECT 63.905 195.855 64.195 195.900 ;
        RECT 65.730 195.840 66.050 195.900 ;
        RECT 74.930 195.840 75.250 196.100 ;
        RECT 80.450 195.840 80.770 196.100 ;
        RECT 85.050 195.840 85.370 196.100 ;
        RECT 86.430 196.040 86.750 196.100 ;
        RECT 87.365 196.040 87.655 196.085 ;
        RECT 86.430 195.900 87.655 196.040 ;
        RECT 86.430 195.840 86.750 195.900 ;
        RECT 87.365 195.855 87.655 195.900 ;
        RECT 18.280 195.220 92.340 195.700 ;
        RECT 43.205 195.020 43.495 195.065 ;
        RECT 43.650 195.020 43.970 195.080 ;
        RECT 43.205 194.880 43.970 195.020 ;
        RECT 43.205 194.835 43.495 194.880 ;
        RECT 43.650 194.820 43.970 194.880 ;
        RECT 44.110 195.020 44.430 195.080 ;
        RECT 44.110 194.880 62.280 195.020 ;
        RECT 44.110 194.820 44.430 194.880 ;
        RECT 33.110 194.680 33.400 194.725 ;
        RECT 35.210 194.680 35.500 194.725 ;
        RECT 36.780 194.680 37.070 194.725 ;
        RECT 33.110 194.540 37.070 194.680 ;
        RECT 43.740 194.680 43.880 194.820 ;
        RECT 62.140 194.740 62.280 194.880 ;
        RECT 80.450 194.820 80.770 195.080 ;
        RECT 83.225 195.020 83.515 195.065 ;
        RECT 84.130 195.020 84.450 195.080 ;
        RECT 83.225 194.880 84.450 195.020 ;
        RECT 83.225 194.835 83.515 194.880 ;
        RECT 84.130 194.820 84.450 194.880 ;
        RECT 45.965 194.680 46.255 194.725 ;
        RECT 43.740 194.540 46.255 194.680 ;
        RECT 33.110 194.495 33.400 194.540 ;
        RECT 35.210 194.495 35.500 194.540 ;
        RECT 36.780 194.495 37.070 194.540 ;
        RECT 45.965 194.495 46.255 194.540 ;
        RECT 51.010 194.680 51.300 194.725 ;
        RECT 52.580 194.680 52.870 194.725 ;
        RECT 54.680 194.680 54.970 194.725 ;
        RECT 51.010 194.540 54.970 194.680 ;
        RECT 51.010 194.495 51.300 194.540 ;
        RECT 52.580 194.495 52.870 194.540 ;
        RECT 54.680 194.495 54.970 194.540 ;
        RECT 62.050 194.480 62.370 194.740 ;
        RECT 62.970 194.680 63.260 194.725 ;
        RECT 64.540 194.680 64.830 194.725 ;
        RECT 66.640 194.680 66.930 194.725 ;
        RECT 62.970 194.540 66.930 194.680 ;
        RECT 62.970 194.495 63.260 194.540 ;
        RECT 64.540 194.495 64.830 194.540 ;
        RECT 66.640 194.495 66.930 194.540 ;
        RECT 72.170 194.680 72.460 194.725 ;
        RECT 73.740 194.680 74.030 194.725 ;
        RECT 75.840 194.680 76.130 194.725 ;
        RECT 72.170 194.540 76.130 194.680 ;
        RECT 72.170 194.495 72.460 194.540 ;
        RECT 73.740 194.495 74.030 194.540 ;
        RECT 75.840 194.495 76.130 194.540 ;
        RECT 78.610 194.680 78.930 194.740 ;
        RECT 78.610 194.540 85.740 194.680 ;
        RECT 78.610 194.480 78.930 194.540 ;
        RECT 33.505 194.340 33.795 194.385 ;
        RECT 34.695 194.340 34.985 194.385 ;
        RECT 37.215 194.340 37.505 194.385 ;
        RECT 33.505 194.200 37.505 194.340 ;
        RECT 33.505 194.155 33.795 194.200 ;
        RECT 34.695 194.155 34.985 194.200 ;
        RECT 37.215 194.155 37.505 194.200 ;
        RECT 50.575 194.340 50.865 194.385 ;
        RECT 53.095 194.340 53.385 194.385 ;
        RECT 54.285 194.340 54.575 194.385 ;
        RECT 50.575 194.200 54.575 194.340 ;
        RECT 50.575 194.155 50.865 194.200 ;
        RECT 53.095 194.155 53.385 194.200 ;
        RECT 54.285 194.155 54.575 194.200 ;
        RECT 55.165 194.340 55.455 194.385 ;
        RECT 62.535 194.340 62.825 194.385 ;
        RECT 65.055 194.340 65.345 194.385 ;
        RECT 66.245 194.340 66.535 194.385 ;
        RECT 55.165 194.200 62.280 194.340 ;
        RECT 55.165 194.155 55.455 194.200 ;
        RECT 32.150 194.000 32.470 194.060 ;
        RECT 53.770 194.045 54.090 194.060 ;
        RECT 32.625 194.000 32.915 194.045 ;
        RECT 41.825 194.000 42.115 194.045 ;
        RECT 44.585 194.000 44.875 194.045 ;
        RECT 32.150 193.860 32.915 194.000 ;
        RECT 32.150 193.800 32.470 193.860 ;
        RECT 32.625 193.815 32.915 193.860 ;
        RECT 39.600 193.860 44.875 194.000 ;
        RECT 33.960 193.660 34.250 193.705 ;
        RECT 34.450 193.660 34.770 193.720 ;
        RECT 33.960 193.520 34.770 193.660 ;
        RECT 33.960 193.475 34.250 193.520 ;
        RECT 34.450 193.460 34.770 193.520 ;
        RECT 39.050 193.320 39.370 193.380 ;
        RECT 39.600 193.365 39.740 193.860 ;
        RECT 41.825 193.815 42.115 193.860 ;
        RECT 44.585 193.815 44.875 193.860 ;
        RECT 53.770 194.000 54.120 194.045 ;
        RECT 59.765 194.000 60.055 194.045 ;
        RECT 62.140 194.000 62.280 194.200 ;
        RECT 62.535 194.200 66.535 194.340 ;
        RECT 62.535 194.155 62.825 194.200 ;
        RECT 65.055 194.155 65.345 194.200 ;
        RECT 66.245 194.155 66.535 194.200 ;
        RECT 67.110 194.140 67.430 194.400 ;
        RECT 71.735 194.340 72.025 194.385 ;
        RECT 74.255 194.340 74.545 194.385 ;
        RECT 75.445 194.340 75.735 194.385 ;
        RECT 71.735 194.200 75.735 194.340 ;
        RECT 71.735 194.155 72.025 194.200 ;
        RECT 74.255 194.155 74.545 194.200 ;
        RECT 75.445 194.155 75.735 194.200 ;
        RECT 82.380 194.200 85.280 194.340 ;
        RECT 67.200 194.000 67.340 194.140 ;
        RECT 76.310 194.000 76.630 194.060 ;
        RECT 53.770 193.860 54.285 194.000 ;
        RECT 59.765 193.860 60.440 194.000 ;
        RECT 62.140 193.860 76.630 194.000 ;
        RECT 53.770 193.815 54.120 193.860 ;
        RECT 59.765 193.815 60.055 193.860 ;
        RECT 53.770 193.800 54.090 193.815 ;
        RECT 39.525 193.320 39.815 193.365 ;
        RECT 39.050 193.180 39.815 193.320 ;
        RECT 39.050 193.120 39.370 193.180 ;
        RECT 39.525 193.135 39.815 193.180 ;
        RECT 44.110 193.120 44.430 193.380 ;
        RECT 45.030 193.320 45.350 193.380 ;
        RECT 46.885 193.320 47.175 193.365 ;
        RECT 45.030 193.180 47.175 193.320 ;
        RECT 45.030 193.120 45.350 193.180 ;
        RECT 46.885 193.135 47.175 193.180 ;
        RECT 48.265 193.320 48.555 193.365 ;
        RECT 53.310 193.320 53.630 193.380 ;
        RECT 48.265 193.180 53.630 193.320 ;
        RECT 48.265 193.135 48.555 193.180 ;
        RECT 53.310 193.120 53.630 193.180 ;
        RECT 59.290 193.120 59.610 193.380 ;
        RECT 60.300 193.365 60.440 193.860 ;
        RECT 76.310 193.800 76.630 193.860 ;
        RECT 79.085 194.000 79.375 194.045 ;
        RECT 80.450 194.000 80.770 194.060 ;
        RECT 82.380 194.045 82.520 194.200 ;
        RECT 79.085 193.860 80.770 194.000 ;
        RECT 79.085 193.815 79.375 193.860 ;
        RECT 80.450 193.800 80.770 193.860 ;
        RECT 81.385 193.815 81.675 194.045 ;
        RECT 82.305 193.815 82.595 194.045 ;
        RECT 65.730 193.705 66.050 193.720 ;
        RECT 74.930 193.705 75.250 193.720 ;
        RECT 65.730 193.660 66.080 193.705 ;
        RECT 74.930 193.660 75.280 193.705 ;
        RECT 78.165 193.660 78.455 193.705 ;
        RECT 80.910 193.660 81.230 193.720 ;
        RECT 65.730 193.520 66.245 193.660 ;
        RECT 74.930 193.520 75.445 193.660 ;
        RECT 78.165 193.520 81.230 193.660 ;
        RECT 81.460 193.660 81.600 193.815 ;
        RECT 84.130 193.800 84.450 194.060 ;
        RECT 85.140 194.045 85.280 194.200 ;
        RECT 85.065 193.815 85.355 194.045 ;
        RECT 85.600 194.000 85.740 194.540 ;
        RECT 85.985 194.000 86.275 194.045 ;
        RECT 85.600 193.860 86.275 194.000 ;
        RECT 85.985 193.815 86.275 193.860 ;
        RECT 86.430 193.850 86.750 194.110 ;
        RECT 86.890 194.045 87.210 194.060 ;
        RECT 86.890 194.000 87.225 194.045 ;
        RECT 87.810 194.000 88.130 194.060 ;
        RECT 86.890 193.860 87.405 194.000 ;
        RECT 87.810 193.860 90.800 194.000 ;
        RECT 86.890 193.815 87.225 193.860 ;
        RECT 82.750 193.660 83.070 193.720 ;
        RECT 81.460 193.520 83.070 193.660 ;
        RECT 65.730 193.475 66.080 193.520 ;
        RECT 74.930 193.475 75.280 193.520 ;
        RECT 78.165 193.475 78.455 193.520 ;
        RECT 65.730 193.460 66.050 193.475 ;
        RECT 74.930 193.460 75.250 193.475 ;
        RECT 80.910 193.460 81.230 193.520 ;
        RECT 82.750 193.460 83.070 193.520 ;
        RECT 84.605 193.475 84.895 193.705 ;
        RECT 85.140 193.660 85.280 193.815 ;
        RECT 86.890 193.800 87.210 193.815 ;
        RECT 87.810 193.800 88.130 193.860 ;
        RECT 90.660 193.720 90.800 193.860 ;
        RECT 85.140 193.520 88.040 193.660 ;
        RECT 60.225 193.320 60.515 193.365 ;
        RECT 60.670 193.320 60.990 193.380 ;
        RECT 60.225 193.180 60.990 193.320 ;
        RECT 60.225 193.135 60.515 193.180 ;
        RECT 60.670 193.120 60.990 193.180 ;
        RECT 68.490 193.320 68.810 193.380 ;
        RECT 69.425 193.320 69.715 193.365 ;
        RECT 68.490 193.180 69.715 193.320 ;
        RECT 68.490 193.120 68.810 193.180 ;
        RECT 69.425 193.135 69.715 193.180 ;
        RECT 80.005 193.320 80.295 193.365 ;
        RECT 83.210 193.320 83.530 193.380 ;
        RECT 80.005 193.180 83.530 193.320 ;
        RECT 84.680 193.320 84.820 193.475 ;
        RECT 87.900 193.380 88.040 193.520 ;
        RECT 90.570 193.460 90.890 193.720 ;
        RECT 85.510 193.320 85.830 193.380 ;
        RECT 87.365 193.320 87.655 193.365 ;
        RECT 84.680 193.180 87.655 193.320 ;
        RECT 80.005 193.135 80.295 193.180 ;
        RECT 83.210 193.120 83.530 193.180 ;
        RECT 85.510 193.120 85.830 193.180 ;
        RECT 87.365 193.135 87.655 193.180 ;
        RECT 87.810 193.120 88.130 193.380 ;
        RECT 18.280 192.500 93.120 192.980 ;
        RECT 19.730 192.300 20.050 192.360 ;
        RECT 51.930 192.300 52.250 192.360 ;
        RECT 19.730 192.160 52.250 192.300 ;
        RECT 19.730 192.100 20.050 192.160 ;
        RECT 51.930 192.100 52.250 192.160 ;
        RECT 64.825 192.300 65.115 192.345 ;
        RECT 66.190 192.300 66.510 192.360 ;
        RECT 64.825 192.160 66.510 192.300 ;
        RECT 64.825 192.115 65.115 192.160 ;
        RECT 66.190 192.100 66.510 192.160 ;
        RECT 71.265 192.300 71.555 192.345 ;
        RECT 71.710 192.300 72.030 192.360 ;
        RECT 71.265 192.160 72.030 192.300 ;
        RECT 71.265 192.115 71.555 192.160 ;
        RECT 71.710 192.100 72.030 192.160 ;
        RECT 80.910 192.300 81.230 192.360 ;
        RECT 86.890 192.300 87.210 192.360 ;
        RECT 80.910 192.160 87.210 192.300 ;
        RECT 80.910 192.100 81.230 192.160 ;
        RECT 86.890 192.100 87.210 192.160 ;
        RECT 27.520 191.960 27.810 192.005 ;
        RECT 28.470 191.960 28.790 192.020 ;
        RECT 27.520 191.820 28.790 191.960 ;
        RECT 27.520 191.775 27.810 191.820 ;
        RECT 28.470 191.760 28.790 191.820 ;
        RECT 34.450 191.760 34.770 192.020 ;
        RECT 44.110 191.960 44.430 192.020 ;
        RECT 46.425 191.960 46.715 192.005 ;
        RECT 83.230 191.960 83.520 192.005 ;
        RECT 84.630 191.960 84.920 192.005 ;
        RECT 86.470 191.960 86.760 192.005 ;
        RECT 44.110 191.820 46.715 191.960 ;
        RECT 44.110 191.760 44.430 191.820 ;
        RECT 46.425 191.775 46.715 191.820 ;
        RECT 51.100 191.820 53.540 191.960 ;
        RECT 33.530 191.620 33.850 191.680 ;
        RECT 34.005 191.620 34.295 191.665 ;
        RECT 33.530 191.480 34.295 191.620 ;
        RECT 33.530 191.420 33.850 191.480 ;
        RECT 34.005 191.435 34.295 191.480 ;
        RECT 34.910 191.420 35.230 191.680 ;
        RECT 36.765 191.435 37.055 191.665 ;
        RECT 26.170 191.080 26.490 191.340 ;
        RECT 27.065 191.280 27.355 191.325 ;
        RECT 28.255 191.280 28.545 191.325 ;
        RECT 30.775 191.280 31.065 191.325 ;
        RECT 36.840 191.280 36.980 191.435 ;
        RECT 45.030 191.420 45.350 191.680 ;
        RECT 45.510 191.435 45.800 191.665 ;
        RECT 27.065 191.140 31.065 191.280 ;
        RECT 27.065 191.095 27.355 191.140 ;
        RECT 28.255 191.095 28.545 191.140 ;
        RECT 30.775 191.095 31.065 191.140 ;
        RECT 33.160 191.140 36.980 191.280 ;
        RECT 39.050 191.280 39.370 191.340 ;
        RECT 39.985 191.280 40.275 191.325 ;
        RECT 39.050 191.140 40.275 191.280 ;
        RECT 33.160 191.000 33.300 191.140 ;
        RECT 39.050 191.080 39.370 191.140 ;
        RECT 39.985 191.095 40.275 191.140 ;
        RECT 43.650 191.280 43.970 191.340 ;
        RECT 45.580 191.280 45.720 191.435 ;
        RECT 46.870 191.420 47.190 191.680 ;
        RECT 47.575 191.620 47.865 191.665 ;
        RECT 51.100 191.620 51.240 191.820 ;
        RECT 53.400 191.680 53.540 191.820 ;
        RECT 83.230 191.820 86.760 191.960 ;
        RECT 83.230 191.775 83.520 191.820 ;
        RECT 84.630 191.775 84.920 191.820 ;
        RECT 86.470 191.775 86.760 191.820 ;
        RECT 90.570 191.760 90.890 192.020 ;
        RECT 47.575 191.480 51.240 191.620 ;
        RECT 47.575 191.435 47.865 191.480 ;
        RECT 51.485 191.435 51.775 191.665 ;
        RECT 43.650 191.140 45.720 191.280 ;
        RECT 43.650 191.080 43.970 191.140 ;
        RECT 26.670 190.940 26.960 190.985 ;
        RECT 28.770 190.940 29.060 190.985 ;
        RECT 30.340 190.940 30.630 190.985 ;
        RECT 26.670 190.800 30.630 190.940 ;
        RECT 26.670 190.755 26.960 190.800 ;
        RECT 28.770 190.755 29.060 190.800 ;
        RECT 30.340 190.755 30.630 190.800 ;
        RECT 33.070 190.740 33.390 191.000 ;
        RECT 37.210 190.940 37.530 191.000 ;
        RECT 51.560 190.940 51.700 191.435 ;
        RECT 52.850 191.420 53.170 191.680 ;
        RECT 53.310 191.620 53.630 191.680 ;
        RECT 59.750 191.620 60.070 191.680 ;
        RECT 53.310 191.480 60.070 191.620 ;
        RECT 53.310 191.420 53.630 191.480 ;
        RECT 59.750 191.420 60.070 191.480 ;
        RECT 62.970 191.620 63.290 191.680 ;
        RECT 66.650 191.620 66.970 191.680 ;
        RECT 62.970 191.480 66.970 191.620 ;
        RECT 62.970 191.420 63.290 191.480 ;
        RECT 66.650 191.420 66.970 191.480 ;
        RECT 68.490 191.620 68.810 191.680 ;
        RECT 74.025 191.620 74.315 191.665 ;
        RECT 68.490 191.480 74.315 191.620 ;
        RECT 68.490 191.420 68.810 191.480 ;
        RECT 74.025 191.435 74.315 191.480 ;
        RECT 76.310 191.620 76.630 191.680 ;
        RECT 81.830 191.620 82.150 191.680 ;
        RECT 82.305 191.620 82.595 191.665 ;
        RECT 76.310 191.480 82.595 191.620 ;
        RECT 76.310 191.420 76.630 191.480 ;
        RECT 81.830 191.420 82.150 191.480 ;
        RECT 82.305 191.435 82.595 191.480 ;
        RECT 83.685 191.620 83.975 191.665 ;
        RECT 85.050 191.620 85.370 191.680 ;
        RECT 83.685 191.480 85.370 191.620 ;
        RECT 83.685 191.435 83.975 191.480 ;
        RECT 85.050 191.420 85.370 191.480 ;
        RECT 57.910 191.280 58.230 191.340 ;
        RECT 63.445 191.280 63.735 191.325 ;
        RECT 72.645 191.280 72.935 191.325 ;
        RECT 57.910 191.140 72.935 191.280 ;
        RECT 57.910 191.080 58.230 191.140 ;
        RECT 63.445 191.095 63.735 191.140 ;
        RECT 72.645 191.095 72.935 191.140 ;
        RECT 85.970 191.280 86.290 191.340 ;
        RECT 87.810 191.280 88.130 191.340 ;
        RECT 85.970 191.140 88.130 191.280 ;
        RECT 85.970 191.080 86.290 191.140 ;
        RECT 87.810 191.080 88.130 191.140 ;
        RECT 53.770 190.940 54.090 191.000 ;
        RECT 37.210 190.800 54.090 190.940 ;
        RECT 37.210 190.740 37.530 190.800 ;
        RECT 53.770 190.740 54.090 190.800 ;
        RECT 56.070 190.940 56.390 191.000 ;
        RECT 62.510 190.940 62.830 191.000 ;
        RECT 56.070 190.800 62.830 190.940 ;
        RECT 56.070 190.740 56.390 190.800 ;
        RECT 62.510 190.740 62.830 190.800 ;
        RECT 82.770 190.940 83.060 190.985 ;
        RECT 85.090 190.940 85.380 190.985 ;
        RECT 86.470 190.940 86.760 190.985 ;
        RECT 82.770 190.800 86.760 190.940 ;
        RECT 82.770 190.755 83.060 190.800 ;
        RECT 85.090 190.755 85.380 190.800 ;
        RECT 86.470 190.755 86.760 190.800 ;
        RECT 43.190 190.400 43.510 190.660 ;
        RECT 48.265 190.600 48.555 190.645 ;
        RECT 51.470 190.600 51.790 190.660 ;
        RECT 48.265 190.460 51.790 190.600 ;
        RECT 48.265 190.415 48.555 190.460 ;
        RECT 51.470 190.400 51.790 190.460 ;
        RECT 51.945 190.600 52.235 190.645 ;
        RECT 52.390 190.600 52.710 190.660 ;
        RECT 51.945 190.460 52.710 190.600 ;
        RECT 51.945 190.415 52.235 190.460 ;
        RECT 52.390 190.400 52.710 190.460 ;
        RECT 54.245 190.600 54.535 190.645 ;
        RECT 56.530 190.600 56.850 190.660 ;
        RECT 54.245 190.460 56.850 190.600 ;
        RECT 54.245 190.415 54.535 190.460 ;
        RECT 56.530 190.400 56.850 190.460 ;
        RECT 59.290 190.600 59.610 190.660 ;
        RECT 62.970 190.600 63.290 190.660 ;
        RECT 59.290 190.460 63.290 190.600 ;
        RECT 59.290 190.400 59.610 190.460 ;
        RECT 62.970 190.400 63.290 190.460 ;
        RECT 72.630 190.400 72.950 190.660 ;
        RECT 18.280 189.780 92.340 190.260 ;
        RECT 28.025 189.580 28.315 189.625 ;
        RECT 28.470 189.580 28.790 189.640 ;
        RECT 28.025 189.440 28.790 189.580 ;
        RECT 28.025 189.395 28.315 189.440 ;
        RECT 28.470 189.380 28.790 189.440 ;
        RECT 33.070 189.580 33.390 189.640 ;
        RECT 33.070 189.440 37.900 189.580 ;
        RECT 33.070 189.380 33.390 189.440 ;
        RECT 33.990 189.240 34.310 189.300 ;
        RECT 35.370 189.240 35.690 189.300 ;
        RECT 37.760 189.285 37.900 189.440 ;
        RECT 43.650 189.380 43.970 189.640 ;
        RECT 44.585 189.580 44.875 189.625 ;
        RECT 46.870 189.580 47.190 189.640 ;
        RECT 52.850 189.580 53.170 189.640 ;
        RECT 44.585 189.440 53.170 189.580 ;
        RECT 44.585 189.395 44.875 189.440 ;
        RECT 46.870 189.380 47.190 189.440 ;
        RECT 52.850 189.380 53.170 189.440 ;
        RECT 56.545 189.580 56.835 189.625 ;
        RECT 59.765 189.580 60.055 189.625 ;
        RECT 56.545 189.440 60.055 189.580 ;
        RECT 56.545 189.395 56.835 189.440 ;
        RECT 59.765 189.395 60.055 189.440 ;
        RECT 60.670 189.580 60.990 189.640 ;
        RECT 60.670 189.440 62.280 189.580 ;
        RECT 60.670 189.380 60.990 189.440 ;
        RECT 33.990 189.100 35.690 189.240 ;
        RECT 33.990 189.040 34.310 189.100 ;
        RECT 35.370 189.040 35.690 189.100 ;
        RECT 37.685 189.240 37.975 189.285 ;
        RECT 39.970 189.240 40.290 189.300 ;
        RECT 37.685 189.100 40.290 189.240 ;
        RECT 37.685 189.055 37.975 189.100 ;
        RECT 39.970 189.040 40.290 189.100 ;
        RECT 42.745 189.240 43.035 189.285 ;
        RECT 44.110 189.240 44.430 189.300 ;
        RECT 42.745 189.100 44.430 189.240 ;
        RECT 42.745 189.055 43.035 189.100 ;
        RECT 44.110 189.040 44.430 189.100 ;
        RECT 59.305 189.240 59.595 189.285 ;
        RECT 61.605 189.240 61.895 189.285 ;
        RECT 59.305 189.100 61.895 189.240 ;
        RECT 62.140 189.240 62.280 189.440 ;
        RECT 74.930 189.380 75.250 189.640 ;
        RECT 75.850 189.380 76.170 189.640 ;
        RECT 65.745 189.240 66.035 189.285 ;
        RECT 62.140 189.100 66.035 189.240 ;
        RECT 59.305 189.055 59.595 189.100 ;
        RECT 61.605 189.055 61.895 189.100 ;
        RECT 65.745 189.055 66.035 189.100 ;
        RECT 68.490 189.240 68.810 189.300 ;
        RECT 70.345 189.240 70.635 189.285 ;
        RECT 68.490 189.100 70.635 189.240 ;
        RECT 68.490 189.040 68.810 189.100 ;
        RECT 70.345 189.055 70.635 189.100 ;
        RECT 33.085 188.900 33.375 188.945 ;
        RECT 28.100 188.760 33.375 188.900 ;
        RECT 28.100 188.605 28.240 188.760 ;
        RECT 33.085 188.715 33.375 188.760 ;
        RECT 34.465 188.900 34.755 188.945 ;
        RECT 35.830 188.900 36.150 188.960 ;
        RECT 34.465 188.760 36.150 188.900 ;
        RECT 34.465 188.715 34.755 188.760 ;
        RECT 35.830 188.700 36.150 188.760 ;
        RECT 53.400 188.760 61.360 188.900 ;
        RECT 28.025 188.375 28.315 188.605 ;
        RECT 28.945 188.560 29.235 188.605 ;
        RECT 33.530 188.560 33.850 188.620 ;
        RECT 28.945 188.420 33.850 188.560 ;
        RECT 28.945 188.375 29.235 188.420 ;
        RECT 33.530 188.360 33.850 188.420 ;
        RECT 34.005 188.375 34.295 188.605 ;
        RECT 34.925 188.375 35.215 188.605 ;
        RECT 34.080 188.220 34.220 188.375 ;
        RECT 34.450 188.220 34.770 188.280 ;
        RECT 34.080 188.080 34.770 188.220 ;
        RECT 35.000 188.220 35.140 188.375 ;
        RECT 35.370 188.360 35.690 188.620 ;
        RECT 36.305 188.560 36.595 188.605 ;
        RECT 37.210 188.560 37.530 188.620 ;
        RECT 36.305 188.420 37.530 188.560 ;
        RECT 36.305 188.375 36.595 188.420 ;
        RECT 37.210 188.360 37.530 188.420 ;
        RECT 39.510 188.560 39.830 188.620 ;
        RECT 40.445 188.560 40.735 188.605 ;
        RECT 44.125 188.560 44.415 188.605 ;
        RECT 39.510 188.420 40.735 188.560 ;
        RECT 39.510 188.360 39.830 188.420 ;
        RECT 40.445 188.375 40.735 188.420 ;
        RECT 40.980 188.420 44.415 188.560 ;
        RECT 40.980 188.220 41.120 188.420 ;
        RECT 44.125 188.375 44.415 188.420 ;
        RECT 48.250 188.360 48.570 188.620 ;
        RECT 51.470 188.360 51.790 188.620 ;
        RECT 52.390 188.360 52.710 188.620 ;
        RECT 53.400 188.605 53.540 188.760 ;
        RECT 53.325 188.375 53.615 188.605 ;
        RECT 53.770 188.560 54.090 188.620 ;
        RECT 56.070 188.605 56.390 188.620 ;
        RECT 53.770 188.420 54.285 188.560 ;
        RECT 53.770 188.360 54.090 188.420 ;
        RECT 55.855 188.375 56.390 188.605 ;
        RECT 56.070 188.360 56.390 188.375 ;
        RECT 56.530 188.560 56.850 188.620 ;
        RECT 57.465 188.560 57.755 188.605 ;
        RECT 56.530 188.420 57.755 188.560 ;
        RECT 56.530 188.360 56.850 188.420 ;
        RECT 57.465 188.375 57.755 188.420 ;
        RECT 58.830 188.360 59.150 188.620 ;
        RECT 61.220 188.560 61.360 188.760 ;
        RECT 62.510 188.700 62.830 188.960 ;
        RECT 63.430 188.900 63.750 188.960 ;
        RECT 64.365 188.900 64.655 188.945 ;
        RECT 75.940 188.900 76.080 189.380 ;
        RECT 63.430 188.760 64.655 188.900 ;
        RECT 63.430 188.700 63.750 188.760 ;
        RECT 64.365 188.715 64.655 188.760 ;
        RECT 72.720 188.760 76.080 188.900 ;
        RECT 62.985 188.560 63.275 188.605 ;
        RECT 63.890 188.560 64.210 188.620 ;
        RECT 72.720 188.605 72.860 188.760 ;
        RECT 61.220 188.420 61.820 188.560 ;
        RECT 35.000 188.080 35.600 188.220 ;
        RECT 34.450 188.020 34.770 188.080 ;
        RECT 35.460 187.880 35.600 188.080 ;
        RECT 38.680 188.080 41.120 188.220 ;
        RECT 41.365 188.220 41.655 188.265 ;
        RECT 42.730 188.220 43.050 188.280 ;
        RECT 41.365 188.080 43.050 188.220 ;
        RECT 38.680 187.940 38.820 188.080 ;
        RECT 41.365 188.035 41.655 188.080 ;
        RECT 38.130 187.880 38.450 187.940 ;
        RECT 35.460 187.740 38.450 187.880 ;
        RECT 38.130 187.680 38.450 187.740 ;
        RECT 38.590 187.680 38.910 187.940 ;
        RECT 39.050 187.680 39.370 187.940 ;
        RECT 39.525 187.880 39.815 187.925 ;
        RECT 41.440 187.880 41.580 188.035 ;
        RECT 42.730 188.020 43.050 188.080 ;
        RECT 39.525 187.740 41.580 187.880 ;
        RECT 39.525 187.695 39.815 187.740 ;
        RECT 47.330 187.680 47.650 187.940 ;
        RECT 51.560 187.880 51.700 188.360 ;
        RECT 52.480 188.220 52.620 188.360 ;
        RECT 54.705 188.220 54.995 188.265 ;
        RECT 52.480 188.080 54.995 188.220 ;
        RECT 54.705 188.035 54.995 188.080 ;
        RECT 55.165 188.220 55.455 188.265 ;
        RECT 56.990 188.220 57.310 188.280 ;
        RECT 55.165 188.080 57.310 188.220 ;
        RECT 55.165 188.035 55.455 188.080 ;
        RECT 56.990 188.020 57.310 188.080 ;
        RECT 57.925 187.880 58.215 187.925 ;
        RECT 51.560 187.740 58.215 187.880 ;
        RECT 57.925 187.695 58.215 187.740 ;
        RECT 61.130 187.680 61.450 187.940 ;
        RECT 61.680 187.880 61.820 188.420 ;
        RECT 62.985 188.420 64.210 188.560 ;
        RECT 62.985 188.375 63.275 188.420 ;
        RECT 63.890 188.360 64.210 188.420 ;
        RECT 72.645 188.375 72.935 188.605 ;
        RECT 75.865 188.560 76.155 188.605 ;
        RECT 75.480 188.420 76.155 188.560 ;
        RECT 63.430 188.220 63.750 188.280 ;
        RECT 64.825 188.220 65.115 188.265 ;
        RECT 67.585 188.220 67.875 188.265 ;
        RECT 63.430 188.080 67.875 188.220 ;
        RECT 63.430 188.020 63.750 188.080 ;
        RECT 64.825 188.035 65.115 188.080 ;
        RECT 67.585 188.035 67.875 188.080 ;
        RECT 68.950 188.020 69.270 188.280 ;
        RECT 75.480 187.940 75.620 188.420 ;
        RECT 75.865 188.375 76.155 188.420 ;
        RECT 65.270 187.880 65.590 187.940 ;
        RECT 61.680 187.740 65.590 187.880 ;
        RECT 65.270 187.680 65.590 187.740 ;
        RECT 71.250 187.680 71.570 187.940 ;
        RECT 72.170 187.680 72.490 187.940 ;
        RECT 72.630 187.880 72.950 187.940 ;
        RECT 73.565 187.880 73.855 187.925 ;
        RECT 72.630 187.740 73.855 187.880 ;
        RECT 72.630 187.680 72.950 187.740 ;
        RECT 73.565 187.695 73.855 187.740 ;
        RECT 75.390 187.680 75.710 187.940 ;
        RECT 18.280 187.060 93.120 187.540 ;
        RECT 26.170 186.860 26.490 186.920 ;
        RECT 34.910 186.860 35.230 186.920 ;
        RECT 36.305 186.860 36.595 186.905 ;
        RECT 40.475 186.860 40.765 186.905 ;
        RECT 26.170 186.720 27.780 186.860 ;
        RECT 26.170 186.660 26.490 186.720 ;
        RECT 26.170 186.225 26.490 186.240 ;
        RECT 27.640 186.225 27.780 186.720 ;
        RECT 34.910 186.720 36.595 186.860 ;
        RECT 34.910 186.660 35.230 186.720 ;
        RECT 36.305 186.675 36.595 186.720 ;
        RECT 37.300 186.720 40.765 186.860 ;
        RECT 35.370 186.520 35.690 186.580 ;
        RECT 37.300 186.520 37.440 186.720 ;
        RECT 40.475 186.675 40.765 186.720 ;
        RECT 40.905 186.860 41.195 186.905 ;
        RECT 41.810 186.860 42.130 186.920 ;
        RECT 40.905 186.720 42.130 186.860 ;
        RECT 40.905 186.675 41.195 186.720 ;
        RECT 41.810 186.660 42.130 186.720 ;
        RECT 58.830 186.860 59.150 186.920 ;
        RECT 70.345 186.860 70.635 186.905 ;
        RECT 58.830 186.720 70.635 186.860 ;
        RECT 58.830 186.660 59.150 186.720 ;
        RECT 32.700 186.380 35.140 186.520 ;
        RECT 26.170 186.180 26.520 186.225 ;
        RECT 27.565 186.180 27.855 186.225 ;
        RECT 32.150 186.180 32.470 186.240 ;
        RECT 32.700 186.225 32.840 186.380 ;
        RECT 26.170 186.040 26.685 186.180 ;
        RECT 27.565 186.040 32.470 186.180 ;
        RECT 26.170 185.995 26.520 186.040 ;
        RECT 27.565 185.995 27.855 186.040 ;
        RECT 26.170 185.980 26.490 185.995 ;
        RECT 32.150 185.980 32.470 186.040 ;
        RECT 32.625 185.995 32.915 186.225 ;
        RECT 33.070 185.980 33.390 186.240 ;
        RECT 34.005 185.995 34.295 186.225 ;
        RECT 22.975 185.840 23.265 185.885 ;
        RECT 25.495 185.840 25.785 185.885 ;
        RECT 26.685 185.840 26.975 185.885 ;
        RECT 30.785 185.840 31.075 185.885 ;
        RECT 22.975 185.700 26.975 185.840 ;
        RECT 22.975 185.655 23.265 185.700 ;
        RECT 25.495 185.655 25.785 185.700 ;
        RECT 26.685 185.655 26.975 185.700 ;
        RECT 27.640 185.700 31.075 185.840 ;
        RECT 23.410 185.500 23.700 185.545 ;
        RECT 24.980 185.500 25.270 185.545 ;
        RECT 27.080 185.500 27.370 185.545 ;
        RECT 23.410 185.360 27.370 185.500 ;
        RECT 23.410 185.315 23.700 185.360 ;
        RECT 24.980 185.315 25.270 185.360 ;
        RECT 27.080 185.315 27.370 185.360 ;
        RECT 20.665 185.160 20.955 185.205 ;
        RECT 27.640 185.160 27.780 185.700 ;
        RECT 30.785 185.655 31.075 185.700 ;
        RECT 30.860 185.500 31.000 185.655 ;
        RECT 33.160 185.500 33.300 185.980 ;
        RECT 30.860 185.360 33.300 185.500 ;
        RECT 20.665 185.020 27.780 185.160 ;
        RECT 28.025 185.160 28.315 185.205 ;
        RECT 28.930 185.160 29.250 185.220 ;
        RECT 28.025 185.020 29.250 185.160 ;
        RECT 20.665 184.975 20.955 185.020 ;
        RECT 28.025 184.975 28.315 185.020 ;
        RECT 28.930 184.960 29.250 185.020 ;
        RECT 31.690 184.960 32.010 185.220 ;
        RECT 34.080 185.160 34.220 185.995 ;
        RECT 34.450 185.980 34.770 186.240 ;
        RECT 35.000 186.225 35.140 186.380 ;
        RECT 35.370 186.380 37.440 186.520 ;
        RECT 46.840 186.520 47.130 186.565 ;
        RECT 47.330 186.520 47.650 186.580 ;
        RECT 63.890 186.520 64.210 186.580 ;
        RECT 35.370 186.320 35.690 186.380 ;
        RECT 34.925 186.180 35.215 186.225 ;
        RECT 34.925 186.040 35.600 186.180 ;
        RECT 34.925 185.995 35.215 186.040 ;
        RECT 35.460 185.840 35.600 186.040 ;
        RECT 35.830 185.980 36.150 186.240 ;
        RECT 37.225 185.995 37.515 186.225 ;
        RECT 39.480 186.180 39.770 186.225 ;
        RECT 39.140 186.040 39.770 186.180 ;
        RECT 39.970 186.150 40.290 186.410 ;
        RECT 46.840 186.380 47.650 186.520 ;
        RECT 46.840 186.335 47.130 186.380 ;
        RECT 47.330 186.320 47.650 186.380 ;
        RECT 57.080 186.380 64.210 186.520 ;
        RECT 57.080 186.240 57.220 186.380 ;
        RECT 37.300 185.840 37.440 185.995 ;
        RECT 35.460 185.700 36.060 185.840 ;
        RECT 34.925 185.160 35.215 185.205 ;
        RECT 34.080 185.020 35.215 185.160 ;
        RECT 34.925 184.975 35.215 185.020 ;
        RECT 35.370 185.160 35.690 185.220 ;
        RECT 35.920 185.160 36.060 185.700 ;
        RECT 36.840 185.700 37.440 185.840 ;
        RECT 36.840 185.560 36.980 185.700 ;
        RECT 38.130 185.640 38.450 185.900 ;
        RECT 38.590 185.640 38.910 185.900 ;
        RECT 36.750 185.300 37.070 185.560 ;
        RECT 37.670 185.300 37.990 185.560 ;
        RECT 38.220 185.160 38.360 185.640 ;
        RECT 39.140 185.500 39.280 186.040 ;
        RECT 39.480 185.995 39.770 186.040 ;
        RECT 41.365 185.995 41.655 186.225 ;
        RECT 42.745 186.180 43.035 186.225 ;
        RECT 43.190 186.180 43.510 186.240 ;
        RECT 42.745 186.040 43.510 186.180 ;
        RECT 42.745 185.995 43.035 186.040 ;
        RECT 40.430 185.840 40.750 185.900 ;
        RECT 41.440 185.840 41.580 185.995 ;
        RECT 43.190 185.980 43.510 186.040 ;
        RECT 56.990 185.980 57.310 186.240 ;
        RECT 60.210 185.980 60.530 186.240 ;
        RECT 61.680 186.225 61.820 186.380 ;
        RECT 63.890 186.320 64.210 186.380 ;
        RECT 61.605 185.995 61.895 186.225 ;
        RECT 62.065 186.180 62.355 186.225 ;
        RECT 62.510 186.180 62.830 186.240 ;
        RECT 64.440 186.225 64.580 186.720 ;
        RECT 70.345 186.675 70.635 186.720 ;
        RECT 79.070 186.860 79.390 186.920 ;
        RECT 79.070 186.720 81.140 186.860 ;
        RECT 79.070 186.660 79.390 186.720 ;
        RECT 68.950 186.320 69.270 186.580 ;
        RECT 77.705 186.520 77.995 186.565 ;
        RECT 77.705 186.380 79.300 186.520 ;
        RECT 77.705 186.335 77.995 186.380 ;
        RECT 62.065 186.040 62.830 186.180 ;
        RECT 62.065 185.995 62.355 186.040 ;
        RECT 62.510 185.980 62.830 186.040 ;
        RECT 64.365 185.995 64.655 186.225 ;
        RECT 65.270 185.980 65.590 186.240 ;
        RECT 65.730 185.980 66.050 186.240 ;
        RECT 67.125 186.180 67.415 186.225 ;
        RECT 69.040 186.180 69.180 186.320 ;
        RECT 67.125 186.040 69.180 186.180 ;
        RECT 67.125 185.995 67.415 186.040 ;
        RECT 71.250 185.980 71.570 186.240 ;
        RECT 73.105 185.995 73.395 186.225 ;
        RECT 40.430 185.700 41.580 185.840 ;
        RECT 44.110 185.840 44.430 185.900 ;
        RECT 45.505 185.840 45.795 185.885 ;
        RECT 44.110 185.700 45.795 185.840 ;
        RECT 40.430 185.640 40.750 185.700 ;
        RECT 44.110 185.640 44.430 185.700 ;
        RECT 45.505 185.655 45.795 185.700 ;
        RECT 46.385 185.840 46.675 185.885 ;
        RECT 47.575 185.840 47.865 185.885 ;
        RECT 50.095 185.840 50.385 185.885 ;
        RECT 46.385 185.700 50.385 185.840 ;
        RECT 46.385 185.655 46.675 185.700 ;
        RECT 47.575 185.655 47.865 185.700 ;
        RECT 50.095 185.655 50.385 185.700 ;
        RECT 60.670 185.640 60.990 185.900 ;
        RECT 69.425 185.840 69.715 185.885 ;
        RECT 69.870 185.840 70.190 185.900 ;
        RECT 73.180 185.840 73.320 185.995 ;
        RECT 75.390 185.980 75.710 186.240 ;
        RECT 77.245 185.995 77.535 186.225 ;
        RECT 78.165 185.995 78.455 186.225 ;
        RECT 69.425 185.700 73.320 185.840 ;
        RECT 69.425 185.655 69.715 185.700 ;
        RECT 69.870 185.640 70.190 185.700 ;
        RECT 74.930 185.640 75.250 185.900 ;
        RECT 77.320 185.840 77.460 185.995 ;
        RECT 77.690 185.840 78.010 185.900 ;
        RECT 77.320 185.700 78.010 185.840 ;
        RECT 78.240 185.840 78.380 185.995 ;
        RECT 78.610 185.980 78.930 186.240 ;
        RECT 79.160 186.225 79.300 186.380 ;
        RECT 79.090 185.995 79.380 186.225 ;
        RECT 79.990 185.980 80.310 186.240 ;
        RECT 80.450 185.980 80.770 186.240 ;
        RECT 81.000 186.225 81.140 186.720 ;
        RECT 83.230 186.520 83.520 186.565 ;
        RECT 84.630 186.520 84.920 186.565 ;
        RECT 86.470 186.520 86.760 186.565 ;
        RECT 83.230 186.380 86.760 186.520 ;
        RECT 83.230 186.335 83.520 186.380 ;
        RECT 84.630 186.335 84.920 186.380 ;
        RECT 86.470 186.335 86.760 186.380 ;
        RECT 80.950 185.995 81.240 186.225 ;
        RECT 81.830 186.180 82.150 186.240 ;
        RECT 82.305 186.180 82.595 186.225 ;
        RECT 86.890 186.180 87.210 186.240 ;
        RECT 81.830 186.040 82.595 186.180 ;
        RECT 81.830 185.980 82.150 186.040 ;
        RECT 82.305 185.995 82.595 186.040 ;
        RECT 82.840 186.040 87.210 186.180 ;
        RECT 82.840 185.840 82.980 186.040 ;
        RECT 86.890 185.980 87.210 186.040 ;
        RECT 78.240 185.700 82.980 185.840 ;
        RECT 77.690 185.640 78.010 185.700 ;
        RECT 83.670 185.640 83.990 185.900 ;
        RECT 45.990 185.500 46.280 185.545 ;
        RECT 48.090 185.500 48.380 185.545 ;
        RECT 49.660 185.500 49.950 185.545 ;
        RECT 39.140 185.360 40.200 185.500 ;
        RECT 35.370 185.020 38.360 185.160 ;
        RECT 40.060 185.160 40.200 185.360 ;
        RECT 45.990 185.360 49.950 185.500 ;
        RECT 45.990 185.315 46.280 185.360 ;
        RECT 48.090 185.315 48.380 185.360 ;
        RECT 49.660 185.315 49.950 185.360 ;
        RECT 62.985 185.500 63.275 185.545 ;
        RECT 64.825 185.500 65.115 185.545 ;
        RECT 62.985 185.360 65.115 185.500 ;
        RECT 62.985 185.315 63.275 185.360 ;
        RECT 64.825 185.315 65.115 185.360 ;
        RECT 82.770 185.500 83.060 185.545 ;
        RECT 85.090 185.500 85.380 185.545 ;
        RECT 86.470 185.500 86.760 185.545 ;
        RECT 82.770 185.360 86.760 185.500 ;
        RECT 82.770 185.315 83.060 185.360 ;
        RECT 85.090 185.315 85.380 185.360 ;
        RECT 86.470 185.315 86.760 185.360 ;
        RECT 42.270 185.160 42.590 185.220 ;
        RECT 40.060 185.020 42.590 185.160 ;
        RECT 35.370 184.960 35.690 185.020 ;
        RECT 42.270 184.960 42.590 185.020 ;
        RECT 44.570 185.160 44.890 185.220 ;
        RECT 50.090 185.160 50.410 185.220 ;
        RECT 52.405 185.160 52.695 185.205 ;
        RECT 44.570 185.020 52.695 185.160 ;
        RECT 44.570 184.960 44.890 185.020 ;
        RECT 50.090 184.960 50.410 185.020 ;
        RECT 52.405 184.975 52.695 185.020 ;
        RECT 62.050 185.160 62.370 185.220 ;
        RECT 63.445 185.160 63.735 185.205 ;
        RECT 62.050 185.020 63.735 185.160 ;
        RECT 62.050 184.960 62.370 185.020 ;
        RECT 63.445 184.975 63.735 185.020 ;
        RECT 68.490 184.960 68.810 185.220 ;
        RECT 70.790 185.160 71.110 185.220 ;
        RECT 71.265 185.160 71.555 185.205 ;
        RECT 73.565 185.160 73.855 185.205 ;
        RECT 70.790 185.020 73.855 185.160 ;
        RECT 70.790 184.960 71.110 185.020 ;
        RECT 71.265 184.975 71.555 185.020 ;
        RECT 73.565 184.975 73.855 185.020 ;
        RECT 81.845 185.160 82.135 185.205 ;
        RECT 85.510 185.160 85.830 185.220 ;
        RECT 81.845 185.020 85.830 185.160 ;
        RECT 81.845 184.975 82.135 185.020 ;
        RECT 85.510 184.960 85.830 185.020 ;
        RECT 90.110 184.960 90.430 185.220 ;
        RECT 18.280 184.340 92.340 184.820 ;
        RECT 26.170 184.140 26.490 184.200 ;
        RECT 27.105 184.140 27.395 184.185 ;
        RECT 31.690 184.140 32.010 184.200 ;
        RECT 26.170 184.000 27.395 184.140 ;
        RECT 26.170 183.940 26.490 184.000 ;
        RECT 27.105 183.955 27.395 184.000 ;
        RECT 29.250 184.000 32.010 184.140 ;
        RECT 29.250 183.460 29.390 184.000 ;
        RECT 31.690 183.940 32.010 184.000 ;
        RECT 32.150 184.140 32.470 184.200 ;
        RECT 34.005 184.140 34.295 184.185 ;
        RECT 37.670 184.140 37.990 184.200 ;
        RECT 40.905 184.140 41.195 184.185 ;
        RECT 44.110 184.140 44.430 184.200 ;
        RECT 32.150 184.000 37.440 184.140 ;
        RECT 32.150 183.940 32.470 184.000 ;
        RECT 34.005 183.955 34.295 184.000 ;
        RECT 34.450 183.800 34.770 183.860 ;
        RECT 36.750 183.800 37.070 183.860 ;
        RECT 34.450 183.660 37.070 183.800 ;
        RECT 37.300 183.800 37.440 184.000 ;
        RECT 37.670 184.000 41.195 184.140 ;
        RECT 37.670 183.940 37.990 184.000 ;
        RECT 40.905 183.955 41.195 184.000 ;
        RECT 41.440 184.000 44.430 184.140 ;
        RECT 41.440 183.800 41.580 184.000 ;
        RECT 44.110 183.940 44.430 184.000 ;
        RECT 47.345 184.140 47.635 184.185 ;
        RECT 48.250 184.140 48.570 184.200 ;
        RECT 56.085 184.140 56.375 184.185 ;
        RECT 56.990 184.140 57.310 184.200 ;
        RECT 47.345 184.000 48.570 184.140 ;
        RECT 47.345 183.955 47.635 184.000 ;
        RECT 48.250 183.940 48.570 184.000 ;
        RECT 51.560 184.000 55.840 184.140 ;
        RECT 37.300 183.660 41.580 183.800 ;
        RECT 41.810 183.800 42.130 183.860 ;
        RECT 42.730 183.800 43.050 183.860 ;
        RECT 44.570 183.800 44.890 183.860 ;
        RECT 51.560 183.800 51.700 184.000 ;
        RECT 41.810 183.660 44.890 183.800 ;
        RECT 34.450 183.600 34.770 183.660 ;
        RECT 36.750 183.600 37.070 183.660 ;
        RECT 41.810 183.600 42.130 183.660 ;
        RECT 42.730 183.600 43.050 183.660 ;
        RECT 44.570 183.600 44.890 183.660 ;
        RECT 45.580 183.660 51.700 183.800 ;
        RECT 28.560 183.320 29.390 183.460 ;
        RECT 33.990 183.460 34.310 183.520 ;
        RECT 38.590 183.460 38.910 183.520 ;
        RECT 45.580 183.460 45.720 183.660 ;
        RECT 47.330 183.460 47.650 183.520 ;
        RECT 33.990 183.320 38.910 183.460 ;
        RECT 28.560 183.165 28.700 183.320 ;
        RECT 33.990 183.260 34.310 183.320 ;
        RECT 38.590 183.260 38.910 183.320 ;
        RECT 40.520 183.320 45.720 183.460 ;
        RECT 46.040 183.320 47.650 183.460 ;
        RECT 55.700 183.460 55.840 184.000 ;
        RECT 56.085 184.000 57.310 184.140 ;
        RECT 56.085 183.955 56.375 184.000 ;
        RECT 56.990 183.940 57.310 184.000 ;
        RECT 64.825 184.140 65.115 184.185 ;
        RECT 67.110 184.140 67.430 184.200 ;
        RECT 64.825 184.000 67.430 184.140 ;
        RECT 64.825 183.955 65.115 184.000 ;
        RECT 67.110 183.940 67.430 184.000 ;
        RECT 79.990 183.940 80.310 184.200 ;
        RECT 83.225 184.140 83.515 184.185 ;
        RECT 84.130 184.140 84.450 184.200 ;
        RECT 83.225 184.000 84.450 184.140 ;
        RECT 83.225 183.955 83.515 184.000 ;
        RECT 84.130 183.940 84.450 184.000 ;
        RECT 86.890 183.940 87.210 184.200 ;
        RECT 87.825 184.140 88.115 184.185 ;
        RECT 88.270 184.140 88.590 184.200 ;
        RECT 87.825 184.000 88.590 184.140 ;
        RECT 87.825 183.955 88.115 184.000 ;
        RECT 65.730 183.800 66.050 183.860 ;
        RECT 68.045 183.800 68.335 183.845 ;
        RECT 73.565 183.800 73.855 183.845 ;
        RECT 85.970 183.800 86.290 183.860 ;
        RECT 65.730 183.660 68.335 183.800 ;
        RECT 65.730 183.600 66.050 183.660 ;
        RECT 68.045 183.615 68.335 183.660 ;
        RECT 68.580 183.660 86.290 183.800 ;
        RECT 59.750 183.460 60.070 183.520 ;
        RECT 68.580 183.460 68.720 183.660 ;
        RECT 73.565 183.615 73.855 183.660 ;
        RECT 85.970 183.600 86.290 183.660 ;
        RECT 70.790 183.460 71.110 183.520 ;
        RECT 87.900 183.460 88.040 183.955 ;
        RECT 88.270 183.940 88.590 184.000 ;
        RECT 55.700 183.320 57.680 183.460 ;
        RECT 40.520 183.180 40.660 183.320 ;
        RECT 28.485 182.935 28.775 183.165 ;
        RECT 28.930 182.920 29.250 183.180 ;
        RECT 29.390 183.120 29.710 183.180 ;
        RECT 29.865 183.120 30.155 183.165 ;
        RECT 29.390 182.980 30.155 183.120 ;
        RECT 29.390 182.920 29.710 182.980 ;
        RECT 29.865 182.935 30.155 182.980 ;
        RECT 40.430 182.920 40.750 183.180 ;
        RECT 41.825 182.935 42.115 183.165 ;
        RECT 27.105 182.780 27.395 182.825 ;
        RECT 31.230 182.780 31.550 182.840 ;
        RECT 27.105 182.640 31.550 182.780 ;
        RECT 41.900 182.780 42.040 182.935 ;
        RECT 42.270 182.920 42.590 183.180 ;
        RECT 44.570 183.120 44.890 183.180 ;
        RECT 46.040 183.165 46.180 183.320 ;
        RECT 47.330 183.260 47.650 183.320 ;
        RECT 57.540 183.180 57.680 183.320 ;
        RECT 59.750 183.320 68.720 183.460 ;
        RECT 69.500 183.320 71.110 183.460 ;
        RECT 59.750 183.260 60.070 183.320 ;
        RECT 44.200 182.980 44.890 183.120 ;
        RECT 42.730 182.780 43.050 182.840 ;
        RECT 44.200 182.825 44.340 182.980 ;
        RECT 44.570 182.920 44.890 182.980 ;
        RECT 45.965 182.935 46.255 183.165 ;
        RECT 46.425 183.120 46.715 183.165 ;
        RECT 47.805 183.120 48.095 183.165 ;
        RECT 46.425 182.980 48.095 183.120 ;
        RECT 46.425 182.935 46.715 182.980 ;
        RECT 47.805 182.935 48.095 182.980 ;
        RECT 48.710 182.920 49.030 183.180 ;
        RECT 50.090 183.165 50.410 183.180 ;
        RECT 50.090 182.935 50.525 183.165 ;
        RECT 51.025 183.120 51.315 183.165 ;
        RECT 52.850 183.120 53.170 183.180 ;
        RECT 51.025 182.980 53.170 183.120 ;
        RECT 51.025 182.935 51.315 182.980 ;
        RECT 50.090 182.920 50.410 182.935 ;
        RECT 52.850 182.920 53.170 182.980 ;
        RECT 56.545 182.935 56.835 183.165 ;
        RECT 43.205 182.780 43.495 182.825 ;
        RECT 41.900 182.640 42.500 182.780 ;
        RECT 27.105 182.595 27.395 182.640 ;
        RECT 31.230 182.580 31.550 182.640 ;
        RECT 42.360 182.500 42.500 182.640 ;
        RECT 42.730 182.640 43.495 182.780 ;
        RECT 42.730 182.580 43.050 182.640 ;
        RECT 43.205 182.595 43.495 182.640 ;
        RECT 44.125 182.595 44.415 182.825 ;
        RECT 45.045 182.780 45.335 182.825 ;
        RECT 49.185 182.780 49.475 182.825 ;
        RECT 45.045 182.640 49.475 182.780 ;
        RECT 45.045 182.595 45.335 182.640 ;
        RECT 49.185 182.595 49.475 182.640 ;
        RECT 49.630 182.580 49.950 182.840 ;
        RECT 56.620 182.500 56.760 182.935 ;
        RECT 57.450 182.920 57.770 183.180 ;
        RECT 69.500 183.165 69.640 183.320 ;
        RECT 70.790 183.260 71.110 183.320 ;
        RECT 81.920 183.320 88.040 183.460 ;
        RECT 69.425 182.935 69.715 183.165 ;
        RECT 69.870 182.920 70.190 183.180 ;
        RECT 70.345 182.935 70.635 183.165 ;
        RECT 71.265 183.120 71.555 183.165 ;
        RECT 72.630 183.120 72.950 183.180 ;
        RECT 81.920 183.165 82.060 183.320 ;
        RECT 71.265 182.980 72.950 183.120 ;
        RECT 71.265 182.935 71.555 182.980 ;
        RECT 70.420 182.780 70.560 182.935 ;
        RECT 72.630 182.920 72.950 182.980 ;
        RECT 80.925 182.935 81.215 183.165 ;
        RECT 81.845 182.935 82.135 183.165 ;
        RECT 82.305 183.120 82.595 183.165 ;
        RECT 84.130 183.120 84.450 183.180 ;
        RECT 82.305 182.980 84.450 183.120 ;
        RECT 82.305 182.935 82.595 182.980 ;
        RECT 72.170 182.780 72.490 182.840 ;
        RECT 70.420 182.640 72.490 182.780 ;
        RECT 81.000 182.780 81.140 182.935 ;
        RECT 84.130 182.920 84.450 182.980 ;
        RECT 84.605 182.935 84.895 183.165 ;
        RECT 84.680 182.780 84.820 182.935 ;
        RECT 85.050 182.920 85.370 183.180 ;
        RECT 85.510 182.920 85.830 183.180 ;
        RECT 86.430 182.920 86.750 183.180 ;
        RECT 88.745 182.780 89.035 182.825 ;
        RECT 90.110 182.780 90.430 182.840 ;
        RECT 81.000 182.640 90.430 182.780 ;
        RECT 72.170 182.580 72.490 182.640 ;
        RECT 88.745 182.595 89.035 182.640 ;
        RECT 90.110 182.580 90.430 182.640 ;
        RECT 28.025 182.440 28.315 182.485 ;
        RECT 29.405 182.440 29.695 182.485 ;
        RECT 28.025 182.300 29.695 182.440 ;
        RECT 28.025 182.255 28.315 182.300 ;
        RECT 29.405 182.255 29.695 182.300 ;
        RECT 42.270 182.240 42.590 182.500 ;
        RECT 56.530 182.240 56.850 182.500 ;
        RECT 84.130 182.440 84.450 182.500 ;
        RECT 86.890 182.440 87.210 182.500 ;
        RECT 87.695 182.440 87.985 182.485 ;
        RECT 84.130 182.300 87.985 182.440 ;
        RECT 84.130 182.240 84.450 182.300 ;
        RECT 86.890 182.240 87.210 182.300 ;
        RECT 87.695 182.255 87.985 182.300 ;
        RECT 18.280 181.620 93.120 182.100 ;
        RECT 35.370 181.420 35.690 181.480 ;
        RECT 37.225 181.420 37.515 181.465 ;
        RECT 35.370 181.280 37.515 181.420 ;
        RECT 35.370 181.220 35.690 181.280 ;
        RECT 37.225 181.235 37.515 181.280 ;
        RECT 41.810 181.220 42.130 181.480 ;
        RECT 42.270 181.420 42.590 181.480 ;
        RECT 48.710 181.420 49.030 181.480 ;
        RECT 42.270 181.280 49.030 181.420 ;
        RECT 42.270 181.220 42.590 181.280 ;
        RECT 48.710 181.220 49.030 181.280 ;
        RECT 61.130 181.220 61.450 181.480 ;
        RECT 62.050 181.220 62.370 181.480 ;
        RECT 38.065 181.080 38.355 181.125 ;
        RECT 38.065 180.940 38.820 181.080 ;
        RECT 38.065 180.895 38.355 180.940 ;
        RECT 38.680 180.460 38.820 180.940 ;
        RECT 39.050 180.880 39.370 181.140 ;
        RECT 40.890 180.740 41.210 180.800 ;
        RECT 41.900 180.785 42.040 181.220 ;
        RECT 41.825 180.740 42.115 180.785 ;
        RECT 40.890 180.600 42.115 180.740 ;
        RECT 40.890 180.540 41.210 180.600 ;
        RECT 41.825 180.555 42.115 180.600 ;
        RECT 42.730 180.540 43.050 180.800 ;
        RECT 59.305 180.555 59.595 180.785 ;
        RECT 60.225 180.740 60.515 180.785 ;
        RECT 60.685 180.740 60.975 180.785 ;
        RECT 61.220 180.740 61.360 181.220 ;
        RECT 60.225 180.600 61.360 180.740 ;
        RECT 61.605 180.740 61.895 180.785 ;
        RECT 62.140 180.740 62.280 181.220 ;
        RECT 61.605 180.600 62.280 180.740 ;
        RECT 60.225 180.555 60.515 180.600 ;
        RECT 60.685 180.555 60.975 180.600 ;
        RECT 61.605 180.555 61.895 180.600 ;
        RECT 62.525 180.555 62.815 180.785 ;
        RECT 38.590 180.400 38.910 180.460 ;
        RECT 42.820 180.400 42.960 180.540 ;
        RECT 38.590 180.260 42.960 180.400 ;
        RECT 59.380 180.400 59.520 180.555 ;
        RECT 61.680 180.400 61.820 180.555 ;
        RECT 62.600 180.400 62.740 180.555 ;
        RECT 68.950 180.540 69.270 180.800 ;
        RECT 71.725 180.740 72.015 180.785 ;
        RECT 75.390 180.740 75.710 180.800 ;
        RECT 77.690 180.740 78.010 180.800 ;
        RECT 71.725 180.600 78.010 180.740 ;
        RECT 71.725 180.555 72.015 180.600 ;
        RECT 75.390 180.540 75.710 180.600 ;
        RECT 77.690 180.540 78.010 180.600 ;
        RECT 78.610 180.540 78.930 180.800 ;
        RECT 59.380 180.260 61.820 180.400 ;
        RECT 62.140 180.260 62.740 180.400 ;
        RECT 69.040 180.400 69.180 180.540 ;
        RECT 69.040 180.260 70.790 180.400 ;
        RECT 38.590 180.200 38.910 180.260 ;
        RECT 41.900 179.780 42.040 180.260 ;
        RECT 49.630 180.060 49.950 180.120 ;
        RECT 58.385 180.060 58.675 180.105 ;
        RECT 62.140 180.060 62.280 180.260 ;
        RECT 49.630 179.920 62.280 180.060 ;
        RECT 70.650 180.060 70.790 180.260 ;
        RECT 72.185 180.215 72.475 180.445 ;
        RECT 72.645 180.215 72.935 180.445 ;
        RECT 72.260 180.060 72.400 180.215 ;
        RECT 70.650 179.920 72.400 180.060 ;
        RECT 72.720 180.060 72.860 180.215 ;
        RECT 73.090 180.200 73.410 180.460 ;
        RECT 78.700 180.060 78.840 180.540 ;
        RECT 72.720 179.920 78.840 180.060 ;
        RECT 49.630 179.860 49.950 179.920 ;
        RECT 58.385 179.875 58.675 179.920 ;
        RECT 38.145 179.720 38.435 179.765 ;
        RECT 40.890 179.720 41.210 179.780 ;
        RECT 38.145 179.580 41.210 179.720 ;
        RECT 38.145 179.535 38.435 179.580 ;
        RECT 40.890 179.520 41.210 179.580 ;
        RECT 41.810 179.520 42.130 179.780 ;
        RECT 43.650 179.720 43.970 179.780 ;
        RECT 61.130 179.720 61.450 179.780 ;
        RECT 43.650 179.580 61.450 179.720 ;
        RECT 43.650 179.520 43.970 179.580 ;
        RECT 61.130 179.520 61.450 179.580 ;
        RECT 62.050 179.720 62.370 179.780 ;
        RECT 63.905 179.720 64.195 179.765 ;
        RECT 72.720 179.720 72.860 179.920 ;
        RECT 62.050 179.580 72.860 179.720 ;
        RECT 74.025 179.720 74.315 179.765 ;
        RECT 75.390 179.720 75.710 179.780 ;
        RECT 74.025 179.580 75.710 179.720 ;
        RECT 62.050 179.520 62.370 179.580 ;
        RECT 63.905 179.535 64.195 179.580 ;
        RECT 74.025 179.535 74.315 179.580 ;
        RECT 75.390 179.520 75.710 179.580 ;
        RECT 18.280 178.900 92.340 179.380 ;
        RECT 37.670 178.700 37.990 178.760 ;
        RECT 39.985 178.700 40.275 178.745 ;
        RECT 37.670 178.560 40.275 178.700 ;
        RECT 37.670 178.500 37.990 178.560 ;
        RECT 39.985 178.515 40.275 178.560 ;
        RECT 40.905 178.515 41.195 178.745 ;
        RECT 55.150 178.700 55.470 178.760 ;
        RECT 56.530 178.700 56.850 178.760 ;
        RECT 58.385 178.700 58.675 178.745 ;
        RECT 60.670 178.700 60.990 178.760 ;
        RECT 78.165 178.700 78.455 178.745 ;
        RECT 55.150 178.560 60.990 178.700 ;
        RECT 24.370 178.360 24.660 178.405 ;
        RECT 26.470 178.360 26.760 178.405 ;
        RECT 28.040 178.360 28.330 178.405 ;
        RECT 24.370 178.220 28.330 178.360 ;
        RECT 24.370 178.175 24.660 178.220 ;
        RECT 26.470 178.175 26.760 178.220 ;
        RECT 28.040 178.175 28.330 178.220 ;
        RECT 30.785 178.175 31.075 178.405 ;
        RECT 24.765 178.020 25.055 178.065 ;
        RECT 25.955 178.020 26.245 178.065 ;
        RECT 28.475 178.020 28.765 178.065 ;
        RECT 24.765 177.880 28.765 178.020 ;
        RECT 30.860 178.020 31.000 178.175 ;
        RECT 33.070 178.160 33.390 178.420 ;
        RECT 38.590 178.360 38.910 178.420 ;
        RECT 33.620 178.220 38.910 178.360 ;
        RECT 30.860 177.880 33.300 178.020 ;
        RECT 24.765 177.835 25.055 177.880 ;
        RECT 25.955 177.835 26.245 177.880 ;
        RECT 28.475 177.835 28.765 177.880 ;
        RECT 22.950 177.680 23.270 177.740 ;
        RECT 23.885 177.680 24.175 177.725 ;
        RECT 22.950 177.540 24.175 177.680 ;
        RECT 22.950 177.480 23.270 177.540 ;
        RECT 23.885 177.495 24.175 177.540 ;
        RECT 32.625 177.495 32.915 177.725 ;
        RECT 25.220 177.340 25.510 177.385 ;
        RECT 32.150 177.340 32.470 177.400 ;
        RECT 25.220 177.200 32.470 177.340 ;
        RECT 25.220 177.155 25.510 177.200 ;
        RECT 32.150 177.140 32.470 177.200 ;
        RECT 31.690 176.800 32.010 177.060 ;
        RECT 32.700 177.000 32.840 177.495 ;
        RECT 33.160 177.340 33.300 177.880 ;
        RECT 33.620 177.725 33.760 178.220 ;
        RECT 38.590 178.160 38.910 178.220 ;
        RECT 40.980 178.080 41.120 178.515 ;
        RECT 55.150 178.500 55.470 178.560 ;
        RECT 56.530 178.500 56.850 178.560 ;
        RECT 58.385 178.515 58.675 178.560 ;
        RECT 60.670 178.500 60.990 178.560 ;
        RECT 70.650 178.560 78.455 178.700 ;
        RECT 43.665 178.360 43.955 178.405 ;
        RECT 59.290 178.360 59.610 178.420 ;
        RECT 43.665 178.220 56.300 178.360 ;
        RECT 43.665 178.175 43.955 178.220 ;
        RECT 33.990 177.820 34.310 178.080 ;
        RECT 39.970 178.020 40.290 178.080 ;
        RECT 40.890 178.020 41.210 178.080 ;
        RECT 55.625 178.020 55.915 178.065 ;
        RECT 35.000 177.880 40.290 178.020 ;
        RECT 35.000 177.725 35.140 177.880 ;
        RECT 39.970 177.820 40.290 177.880 ;
        RECT 40.520 177.880 41.210 178.020 ;
        RECT 33.545 177.495 33.835 177.725 ;
        RECT 34.925 177.495 35.215 177.725 ;
        RECT 35.845 177.495 36.135 177.725 ;
        RECT 38.130 177.680 38.450 177.740 ;
        RECT 40.520 177.680 40.660 177.880 ;
        RECT 40.890 177.820 41.210 177.880 ;
        RECT 50.180 177.880 55.915 178.020 ;
        RECT 38.130 177.540 40.660 177.680 ;
        RECT 35.370 177.340 35.690 177.400 ;
        RECT 35.920 177.340 36.060 177.495 ;
        RECT 38.130 177.480 38.450 177.540 ;
        RECT 41.810 177.480 42.130 177.740 ;
        RECT 42.745 177.495 43.035 177.725 ;
        RECT 43.650 177.680 43.970 177.740 ;
        RECT 44.125 177.680 44.415 177.725 ;
        RECT 43.650 177.540 44.415 177.680 ;
        RECT 39.065 177.340 39.355 177.385 ;
        RECT 33.160 177.200 39.355 177.340 ;
        RECT 35.370 177.140 35.690 177.200 ;
        RECT 39.065 177.155 39.355 177.200 ;
        RECT 39.510 177.140 39.830 177.400 ;
        RECT 34.450 177.000 34.770 177.060 ;
        RECT 32.700 176.860 34.770 177.000 ;
        RECT 34.450 176.800 34.770 176.860 ;
        RECT 38.590 176.800 38.910 177.060 ;
        RECT 39.600 177.000 39.740 177.140 ;
        RECT 40.065 177.000 40.355 177.045 ;
        RECT 42.820 177.000 42.960 177.495 ;
        RECT 43.650 177.480 43.970 177.540 ;
        RECT 44.125 177.495 44.415 177.540 ;
        RECT 47.790 177.480 48.110 177.740 ;
        RECT 50.180 177.725 50.320 177.880 ;
        RECT 55.625 177.835 55.915 177.880 ;
        RECT 50.105 177.495 50.395 177.725 ;
        RECT 51.010 177.480 51.330 177.740 ;
        RECT 52.405 177.680 52.695 177.725 ;
        RECT 52.850 177.680 53.170 177.740 ;
        RECT 52.405 177.540 53.170 177.680 ;
        RECT 52.405 177.495 52.695 177.540 ;
        RECT 52.850 177.480 53.170 177.540 ;
        RECT 53.310 177.680 53.630 177.740 ;
        RECT 54.705 177.680 54.995 177.725 ;
        RECT 53.310 177.540 54.995 177.680 ;
        RECT 53.310 177.480 53.630 177.540 ;
        RECT 54.705 177.495 54.995 177.540 ;
        RECT 55.150 177.480 55.470 177.740 ;
        RECT 56.160 177.725 56.300 178.220 ;
        RECT 59.290 178.220 69.640 178.360 ;
        RECT 59.290 178.160 59.610 178.220 ;
        RECT 61.130 177.820 61.450 178.080 ;
        RECT 56.085 177.680 56.375 177.725 ;
        RECT 61.220 177.680 61.360 177.820 ;
        RECT 62.525 177.680 62.815 177.725 ;
        RECT 56.085 177.540 60.440 177.680 ;
        RECT 61.220 177.540 62.815 177.680 ;
        RECT 56.085 177.495 56.375 177.540 ;
        RECT 51.470 177.385 51.790 177.400 ;
        RECT 50.565 177.155 50.855 177.385 ;
        RECT 51.470 177.340 52.005 177.385 ;
        RECT 53.770 177.340 54.090 177.400 ;
        RECT 51.470 177.200 54.090 177.340 ;
        RECT 51.470 177.155 52.005 177.200 ;
        RECT 39.600 176.860 42.960 177.000 ;
        RECT 43.190 177.000 43.510 177.060 ;
        RECT 45.045 177.000 45.335 177.045 ;
        RECT 43.190 176.860 45.335 177.000 ;
        RECT 40.065 176.815 40.355 176.860 ;
        RECT 43.190 176.800 43.510 176.860 ;
        RECT 45.045 176.815 45.335 176.860 ;
        RECT 46.870 176.800 47.190 177.060 ;
        RECT 48.250 177.000 48.570 177.060 ;
        RECT 49.185 177.000 49.475 177.045 ;
        RECT 48.250 176.860 49.475 177.000 ;
        RECT 50.640 177.000 50.780 177.155 ;
        RECT 51.470 177.140 51.790 177.155 ;
        RECT 53.770 177.140 54.090 177.200 ;
        RECT 57.465 177.340 57.755 177.385 ;
        RECT 59.765 177.340 60.055 177.385 ;
        RECT 57.465 177.200 60.055 177.340 ;
        RECT 60.300 177.340 60.440 177.540 ;
        RECT 62.525 177.495 62.815 177.540 ;
        RECT 62.970 177.480 63.290 177.740 ;
        RECT 60.765 177.340 61.055 177.385 ;
        RECT 63.060 177.340 63.200 177.480 ;
        RECT 69.500 177.400 69.640 178.220 ;
        RECT 70.650 178.020 70.790 178.560 ;
        RECT 78.165 178.515 78.455 178.560 ;
        RECT 71.290 178.360 71.580 178.405 ;
        RECT 73.390 178.360 73.680 178.405 ;
        RECT 74.960 178.360 75.250 178.405 ;
        RECT 71.290 178.220 75.250 178.360 ;
        RECT 71.290 178.175 71.580 178.220 ;
        RECT 73.390 178.175 73.680 178.220 ;
        RECT 74.960 178.175 75.250 178.220 ;
        RECT 77.690 178.360 78.010 178.420 ;
        RECT 77.690 178.220 81.140 178.360 ;
        RECT 77.690 178.160 78.010 178.220 ;
        RECT 81.000 178.065 81.140 178.220 ;
        RECT 70.420 177.880 70.790 178.020 ;
        RECT 71.685 178.020 71.975 178.065 ;
        RECT 72.875 178.020 73.165 178.065 ;
        RECT 75.395 178.020 75.685 178.065 ;
        RECT 71.685 177.880 75.685 178.020 ;
        RECT 70.420 177.725 70.560 177.880 ;
        RECT 71.685 177.835 71.975 177.880 ;
        RECT 72.875 177.835 73.165 177.880 ;
        RECT 75.395 177.835 75.685 177.880 ;
        RECT 80.925 177.835 81.215 178.065 ;
        RECT 85.970 177.820 86.290 178.080 ;
        RECT 70.345 177.495 70.635 177.725 ;
        RECT 70.805 177.680 71.095 177.725 ;
        RECT 80.450 177.680 80.770 177.740 ;
        RECT 70.805 177.540 80.770 177.680 ;
        RECT 70.805 177.495 71.095 177.540 ;
        RECT 80.450 177.480 80.770 177.540 ;
        RECT 87.365 177.495 87.655 177.725 ;
        RECT 60.300 177.200 61.055 177.340 ;
        RECT 57.465 177.155 57.755 177.200 ;
        RECT 59.765 177.155 60.055 177.200 ;
        RECT 60.765 177.155 61.055 177.200 ;
        RECT 61.220 177.200 63.200 177.340 ;
        RECT 69.410 177.340 69.730 177.400 ;
        RECT 72.140 177.340 72.430 177.385 ;
        RECT 72.630 177.340 72.950 177.400 ;
        RECT 69.410 177.200 70.560 177.340 ;
        RECT 52.865 177.000 53.155 177.045 ;
        RECT 50.640 176.860 53.155 177.000 ;
        RECT 48.250 176.800 48.570 176.860 ;
        RECT 49.185 176.815 49.475 176.860 ;
        RECT 52.865 176.815 53.155 176.860 ;
        RECT 53.310 177.000 53.630 177.060 ;
        RECT 58.465 177.000 58.755 177.045 ;
        RECT 53.310 176.860 58.755 177.000 ;
        RECT 59.840 177.000 59.980 177.155 ;
        RECT 61.220 177.000 61.360 177.200 ;
        RECT 69.410 177.140 69.730 177.200 ;
        RECT 59.840 176.860 61.360 177.000 ;
        RECT 53.310 176.800 53.630 176.860 ;
        RECT 58.465 176.815 58.755 176.860 ;
        RECT 61.590 176.800 61.910 177.060 ;
        RECT 63.905 177.000 64.195 177.045 ;
        RECT 68.490 177.000 68.810 177.060 ;
        RECT 63.905 176.860 68.810 177.000 ;
        RECT 63.905 176.815 64.195 176.860 ;
        RECT 68.490 176.800 68.810 176.860 ;
        RECT 69.870 176.800 70.190 177.060 ;
        RECT 70.420 177.000 70.560 177.200 ;
        RECT 72.140 177.200 72.950 177.340 ;
        RECT 72.140 177.155 72.430 177.200 ;
        RECT 72.630 177.140 72.950 177.200 ;
        RECT 76.770 177.340 77.090 177.400 ;
        RECT 85.065 177.340 85.355 177.385 ;
        RECT 76.770 177.200 85.355 177.340 ;
        RECT 76.770 177.140 77.090 177.200 ;
        RECT 85.065 177.155 85.355 177.200 ;
        RECT 86.890 177.340 87.210 177.400 ;
        RECT 87.440 177.340 87.580 177.495 ;
        RECT 88.270 177.480 88.590 177.740 ;
        RECT 86.890 177.200 87.580 177.340 ;
        RECT 88.360 177.340 88.500 177.480 ;
        RECT 90.570 177.340 90.890 177.400 ;
        RECT 88.360 177.200 90.890 177.340 ;
        RECT 86.890 177.140 87.210 177.200 ;
        RECT 90.570 177.140 90.890 177.200 ;
        RECT 73.090 177.000 73.410 177.060 ;
        RECT 70.420 176.860 73.410 177.000 ;
        RECT 73.090 176.800 73.410 176.860 ;
        RECT 80.910 177.000 81.230 177.060 ;
        RECT 83.225 177.000 83.515 177.045 ;
        RECT 80.910 176.860 83.515 177.000 ;
        RECT 80.910 176.800 81.230 176.860 ;
        RECT 83.225 176.815 83.515 176.860 ;
        RECT 85.525 177.000 85.815 177.045 ;
        RECT 87.825 177.000 88.115 177.045 ;
        RECT 85.525 176.860 88.115 177.000 ;
        RECT 85.525 176.815 85.815 176.860 ;
        RECT 87.825 176.815 88.115 176.860 ;
        RECT 18.280 176.180 93.120 176.660 ;
        RECT 31.690 175.780 32.010 176.040 ;
        RECT 32.150 175.780 32.470 176.040 ;
        RECT 33.070 175.980 33.390 176.040 ;
        RECT 35.385 175.980 35.675 176.025 ;
        RECT 33.070 175.840 35.675 175.980 ;
        RECT 33.070 175.780 33.390 175.840 ;
        RECT 35.385 175.795 35.675 175.840 ;
        RECT 38.590 175.780 38.910 176.040 ;
        RECT 39.970 175.780 40.290 176.040 ;
        RECT 51.470 175.780 51.790 176.040 ;
        RECT 57.450 175.980 57.770 176.040 ;
        RECT 58.385 175.980 58.675 176.025 ;
        RECT 57.450 175.840 58.675 175.980 ;
        RECT 57.450 175.780 57.770 175.840 ;
        RECT 58.385 175.795 58.675 175.840 ;
        RECT 61.590 175.780 61.910 176.040 ;
        RECT 62.050 175.980 62.370 176.040 ;
        RECT 65.730 175.980 66.050 176.040 ;
        RECT 62.050 175.840 66.050 175.980 ;
        RECT 62.050 175.780 62.370 175.840 ;
        RECT 65.730 175.780 66.050 175.840 ;
        RECT 68.505 175.980 68.795 176.025 ;
        RECT 68.950 175.980 69.270 176.040 ;
        RECT 68.505 175.840 69.270 175.980 ;
        RECT 68.505 175.795 68.795 175.840 ;
        RECT 68.950 175.780 69.270 175.840 ;
        RECT 72.630 175.980 72.950 176.040 ;
        RECT 74.025 175.980 74.315 176.025 ;
        RECT 79.990 175.980 80.310 176.040 ;
        RECT 72.630 175.840 74.315 175.980 ;
        RECT 72.630 175.780 72.950 175.840 ;
        RECT 74.025 175.795 74.315 175.840 ;
        RECT 76.860 175.840 80.310 175.980 ;
        RECT 31.780 175.345 31.920 175.780 ;
        RECT 31.705 175.115 31.995 175.345 ;
        RECT 32.625 175.300 32.915 175.345 ;
        RECT 33.530 175.300 33.850 175.360 ;
        RECT 32.625 175.160 33.850 175.300 ;
        RECT 32.625 175.115 32.915 175.160 ;
        RECT 33.530 175.100 33.850 175.160 ;
        RECT 34.925 175.300 35.215 175.345 ;
        RECT 35.370 175.300 35.690 175.360 ;
        RECT 34.925 175.160 35.690 175.300 ;
        RECT 34.925 175.115 35.215 175.160 ;
        RECT 35.370 175.100 35.690 175.160 ;
        RECT 35.845 175.300 36.135 175.345 ;
        RECT 37.670 175.300 37.990 175.360 ;
        RECT 35.845 175.160 37.990 175.300 ;
        RECT 38.680 175.300 38.820 175.780 ;
        RECT 43.190 175.640 43.510 175.700 ;
        RECT 40.060 175.500 43.510 175.640 ;
        RECT 39.525 175.300 39.815 175.345 ;
        RECT 38.680 175.160 39.815 175.300 ;
        RECT 35.845 175.115 36.135 175.160 ;
        RECT 37.670 175.100 37.990 175.160 ;
        RECT 39.525 175.115 39.815 175.160 ;
        RECT 28.485 174.960 28.775 175.005 ;
        RECT 29.850 174.960 30.170 175.020 ;
        RECT 28.485 174.820 30.170 174.960 ;
        RECT 28.485 174.775 28.775 174.820 ;
        RECT 29.850 174.760 30.170 174.820 ;
        RECT 34.450 174.960 34.770 175.020 ;
        RECT 40.060 174.960 40.200 175.500 ;
        RECT 43.190 175.440 43.510 175.500 ;
        RECT 45.920 175.640 46.210 175.685 ;
        RECT 46.870 175.640 47.190 175.700 ;
        RECT 45.920 175.500 47.190 175.640 ;
        RECT 45.920 175.455 46.210 175.500 ;
        RECT 46.870 175.440 47.190 175.500 ;
        RECT 51.930 175.440 52.250 175.700 ;
        RECT 61.680 175.640 61.820 175.780 ;
        RECT 61.220 175.500 61.820 175.640 ;
        RECT 61.220 175.345 61.360 175.500 ;
        RECT 61.145 175.115 61.435 175.345 ;
        RECT 61.605 175.300 61.895 175.345 ;
        RECT 62.140 175.300 62.280 175.780 ;
        RECT 63.445 175.640 63.735 175.685 ;
        RECT 66.650 175.640 66.970 175.700 ;
        RECT 76.860 175.640 77.000 175.840 ;
        RECT 79.990 175.780 80.310 175.840 ;
        RECT 80.910 175.780 81.230 176.040 ;
        RECT 88.270 175.980 88.590 176.040 ;
        RECT 81.460 175.840 88.590 175.980 ;
        RECT 81.000 175.640 81.140 175.780 ;
        RECT 63.445 175.500 65.040 175.640 ;
        RECT 63.445 175.455 63.735 175.500 ;
        RECT 61.605 175.160 62.280 175.300 ;
        RECT 61.605 175.115 61.895 175.160 ;
        RECT 62.525 175.115 62.815 175.345 ;
        RECT 34.450 174.820 40.200 174.960 ;
        RECT 34.450 174.760 34.770 174.820 ;
        RECT 44.570 174.760 44.890 175.020 ;
        RECT 45.465 174.960 45.755 175.005 ;
        RECT 46.655 174.960 46.945 175.005 ;
        RECT 49.175 174.960 49.465 175.005 ;
        RECT 62.600 174.960 62.740 175.115 ;
        RECT 63.890 175.100 64.210 175.360 ;
        RECT 64.900 175.345 65.040 175.500 ;
        RECT 65.820 175.500 77.000 175.640 ;
        RECT 64.825 175.115 65.115 175.345 ;
        RECT 65.270 175.100 65.590 175.360 ;
        RECT 65.820 175.345 65.960 175.500 ;
        RECT 66.650 175.440 66.970 175.500 ;
        RECT 65.745 175.115 66.035 175.345 ;
        RECT 67.585 175.300 67.875 175.345 ;
        RECT 68.490 175.300 68.810 175.360 ;
        RECT 67.585 175.160 68.810 175.300 ;
        RECT 67.585 175.115 67.875 175.160 ;
        RECT 68.490 175.100 68.810 175.160 ;
        RECT 68.965 175.300 69.255 175.345 ;
        RECT 69.410 175.300 69.730 175.360 ;
        RECT 68.965 175.160 69.730 175.300 ;
        RECT 68.965 175.115 69.255 175.160 ;
        RECT 69.410 175.100 69.730 175.160 ;
        RECT 69.870 175.300 70.190 175.360 ;
        RECT 74.945 175.300 75.235 175.345 ;
        RECT 69.870 175.160 75.235 175.300 ;
        RECT 69.870 175.100 70.190 175.160 ;
        RECT 74.945 175.115 75.235 175.160 ;
        RECT 75.390 175.300 75.710 175.360 ;
        RECT 76.325 175.300 76.615 175.345 ;
        RECT 75.390 175.160 76.615 175.300 ;
        RECT 75.390 175.100 75.710 175.160 ;
        RECT 76.325 175.115 76.615 175.160 ;
        RECT 70.345 174.960 70.635 175.005 ;
        RECT 45.465 174.820 49.465 174.960 ;
        RECT 45.465 174.775 45.755 174.820 ;
        RECT 46.655 174.775 46.945 174.820 ;
        RECT 49.175 174.775 49.465 174.820 ;
        RECT 62.140 174.820 62.740 174.960 ;
        RECT 64.440 174.820 70.635 174.960 ;
        RECT 33.990 174.620 34.310 174.680 ;
        RECT 44.110 174.620 44.430 174.680 ;
        RECT 33.990 174.480 44.430 174.620 ;
        RECT 33.990 174.420 34.310 174.480 ;
        RECT 44.110 174.420 44.430 174.480 ;
        RECT 45.070 174.620 45.360 174.665 ;
        RECT 47.170 174.620 47.460 174.665 ;
        RECT 48.740 174.620 49.030 174.665 ;
        RECT 45.070 174.480 49.030 174.620 ;
        RECT 45.070 174.435 45.360 174.480 ;
        RECT 47.170 174.435 47.460 174.480 ;
        RECT 48.740 174.435 49.030 174.480 ;
        RECT 25.250 174.080 25.570 174.340 ;
        RECT 40.890 174.280 41.210 174.340 ;
        RECT 53.310 174.280 53.630 174.340 ;
        RECT 61.130 174.280 61.450 174.340 ;
        RECT 40.890 174.140 61.450 174.280 ;
        RECT 62.140 174.280 62.280 174.820 ;
        RECT 64.440 174.280 64.580 174.820 ;
        RECT 70.345 174.775 70.635 174.820 ;
        RECT 73.105 174.775 73.395 175.005 ;
        RECT 76.860 174.960 77.000 175.500 ;
        RECT 79.160 175.500 81.140 175.640 ;
        RECT 77.245 175.300 77.535 175.345 ;
        RECT 77.690 175.300 78.010 175.360 ;
        RECT 78.165 175.300 78.455 175.345 ;
        RECT 77.245 175.160 78.455 175.300 ;
        RECT 77.245 175.115 77.535 175.160 ;
        RECT 77.690 175.100 78.010 175.160 ;
        RECT 78.165 175.115 78.455 175.160 ;
        RECT 75.480 174.820 77.000 174.960 ;
        RECT 65.270 174.620 65.590 174.680 ;
        RECT 68.950 174.620 69.270 174.680 ;
        RECT 71.710 174.620 72.030 174.680 ;
        RECT 73.180 174.620 73.320 174.775 ;
        RECT 75.480 174.665 75.620 174.820 ;
        RECT 65.270 174.480 67.800 174.620 ;
        RECT 65.270 174.420 65.590 174.480 ;
        RECT 62.140 174.140 64.580 174.280 ;
        RECT 66.190 174.280 66.510 174.340 ;
        RECT 67.660 174.325 67.800 174.480 ;
        RECT 68.950 174.480 73.320 174.620 ;
        RECT 68.950 174.420 69.270 174.480 ;
        RECT 71.710 174.420 72.030 174.480 ;
        RECT 75.405 174.435 75.695 174.665 ;
        RECT 75.865 174.435 76.155 174.665 ;
        RECT 67.125 174.280 67.415 174.325 ;
        RECT 66.190 174.140 67.415 174.280 ;
        RECT 40.890 174.080 41.210 174.140 ;
        RECT 53.310 174.080 53.630 174.140 ;
        RECT 61.130 174.080 61.450 174.140 ;
        RECT 66.190 174.080 66.510 174.140 ;
        RECT 67.125 174.095 67.415 174.140 ;
        RECT 67.585 174.280 67.875 174.325 ;
        RECT 75.940 174.280 76.080 174.435 ;
        RECT 67.585 174.140 76.080 174.280 ;
        RECT 78.240 174.280 78.380 175.115 ;
        RECT 78.610 175.100 78.930 175.360 ;
        RECT 79.160 175.345 79.300 175.500 ;
        RECT 79.085 175.115 79.375 175.345 ;
        RECT 80.925 175.300 81.215 175.345 ;
        RECT 81.460 175.300 81.600 175.840 ;
        RECT 88.270 175.780 88.590 175.840 ;
        RECT 83.230 175.640 83.520 175.685 ;
        RECT 84.630 175.640 84.920 175.685 ;
        RECT 86.470 175.640 86.760 175.685 ;
        RECT 83.230 175.500 86.760 175.640 ;
        RECT 83.230 175.455 83.520 175.500 ;
        RECT 84.630 175.455 84.920 175.500 ;
        RECT 86.470 175.455 86.760 175.500 ;
        RECT 80.925 175.160 81.600 175.300 ;
        RECT 81.845 175.300 82.135 175.345 ;
        RECT 83.685 175.300 83.975 175.345 ;
        RECT 81.845 175.160 83.975 175.300 ;
        RECT 80.925 175.115 81.215 175.160 ;
        RECT 81.845 175.115 82.135 175.160 ;
        RECT 83.685 175.115 83.975 175.160 ;
        RECT 78.700 174.960 78.840 175.100 ;
        RECT 79.545 174.960 79.835 175.005 ;
        RECT 78.700 174.820 79.835 174.960 ;
        RECT 79.545 174.775 79.835 174.820 ;
        RECT 79.990 174.760 80.310 175.020 ;
        RECT 80.450 174.960 80.770 175.020 ;
        RECT 82.305 174.960 82.595 175.005 ;
        RECT 80.450 174.820 82.595 174.960 ;
        RECT 80.450 174.760 80.770 174.820 ;
        RECT 82.305 174.775 82.595 174.820 ;
        RECT 82.770 174.620 83.060 174.665 ;
        RECT 85.090 174.620 85.380 174.665 ;
        RECT 86.470 174.620 86.760 174.665 ;
        RECT 82.770 174.480 86.760 174.620 ;
        RECT 82.770 174.435 83.060 174.480 ;
        RECT 85.090 174.435 85.380 174.480 ;
        RECT 86.470 174.435 86.760 174.480 ;
        RECT 85.970 174.280 86.290 174.340 ;
        RECT 78.240 174.140 86.290 174.280 ;
        RECT 67.585 174.095 67.875 174.140 ;
        RECT 85.970 174.080 86.290 174.140 ;
        RECT 90.125 174.280 90.415 174.325 ;
        RECT 90.570 174.280 90.890 174.340 ;
        RECT 90.125 174.140 90.890 174.280 ;
        RECT 90.125 174.095 90.415 174.140 ;
        RECT 90.570 174.080 90.890 174.140 ;
        RECT 18.280 173.460 92.340 173.940 ;
        RECT 29.850 173.060 30.170 173.320 ;
        RECT 37.685 173.260 37.975 173.305 ;
        RECT 41.365 173.260 41.655 173.305 ;
        RECT 41.810 173.260 42.130 173.320 ;
        RECT 37.685 173.120 41.120 173.260 ;
        RECT 37.685 173.075 37.975 173.120 ;
        RECT 23.450 172.920 23.740 172.965 ;
        RECT 25.550 172.920 25.840 172.965 ;
        RECT 27.120 172.920 27.410 172.965 ;
        RECT 23.450 172.780 27.410 172.920 ;
        RECT 23.450 172.735 23.740 172.780 ;
        RECT 25.550 172.735 25.840 172.780 ;
        RECT 27.120 172.735 27.410 172.780 ;
        RECT 31.705 172.735 31.995 172.965 ;
        RECT 35.385 172.735 35.675 172.965 ;
        RECT 35.830 172.920 36.150 172.980 ;
        RECT 38.605 172.920 38.895 172.965 ;
        RECT 35.830 172.780 38.895 172.920 ;
        RECT 40.980 172.920 41.120 173.120 ;
        RECT 41.365 173.120 42.130 173.260 ;
        RECT 41.365 173.075 41.655 173.120 ;
        RECT 41.810 173.060 42.130 173.120 ;
        RECT 46.885 173.260 47.175 173.305 ;
        RECT 47.790 173.260 48.110 173.320 ;
        RECT 46.885 173.120 48.110 173.260 ;
        RECT 46.885 173.075 47.175 173.120 ;
        RECT 47.790 173.060 48.110 173.120 ;
        RECT 71.710 173.060 72.030 173.320 ;
        RECT 79.990 173.260 80.310 173.320 ;
        RECT 81.385 173.260 81.675 173.305 ;
        RECT 79.990 173.120 81.675 173.260 ;
        RECT 79.990 173.060 80.310 173.120 ;
        RECT 81.385 173.075 81.675 173.120 ;
        RECT 43.650 172.920 43.970 172.980 ;
        RECT 40.980 172.780 43.970 172.920 ;
        RECT 23.845 172.580 24.135 172.625 ;
        RECT 25.035 172.580 25.325 172.625 ;
        RECT 27.555 172.580 27.845 172.625 ;
        RECT 23.845 172.440 27.845 172.580 ;
        RECT 23.845 172.395 24.135 172.440 ;
        RECT 25.035 172.395 25.325 172.440 ;
        RECT 27.555 172.395 27.845 172.440 ;
        RECT 22.950 172.240 23.270 172.300 ;
        RECT 28.930 172.240 29.250 172.300 ;
        RECT 31.780 172.240 31.920 172.735 ;
        RECT 22.950 172.100 29.250 172.240 ;
        RECT 22.950 172.040 23.270 172.100 ;
        RECT 28.930 172.040 29.250 172.100 ;
        RECT 30.400 172.100 31.920 172.240 ;
        RECT 33.085 172.240 33.375 172.285 ;
        RECT 35.460 172.240 35.600 172.735 ;
        RECT 35.830 172.720 36.150 172.780 ;
        RECT 38.605 172.735 38.895 172.780 ;
        RECT 43.650 172.720 43.970 172.780 ;
        RECT 58.845 172.920 59.135 172.965 ;
        RECT 62.525 172.920 62.815 172.965 ;
        RECT 58.845 172.780 62.815 172.920 ;
        RECT 58.845 172.735 59.135 172.780 ;
        RECT 62.525 172.735 62.815 172.780 ;
        RECT 65.310 172.920 65.600 172.965 ;
        RECT 67.410 172.920 67.700 172.965 ;
        RECT 68.980 172.920 69.270 172.965 ;
        RECT 65.310 172.780 69.270 172.920 ;
        RECT 65.310 172.735 65.600 172.780 ;
        RECT 67.410 172.735 67.700 172.780 ;
        RECT 68.980 172.735 69.270 172.780 ;
        RECT 77.230 172.920 77.550 172.980 ;
        RECT 77.230 172.780 84.360 172.920 ;
        RECT 77.230 172.720 77.550 172.780 ;
        RECT 36.765 172.580 37.055 172.625 ;
        RECT 37.670 172.580 37.990 172.640 ;
        RECT 36.765 172.440 37.990 172.580 ;
        RECT 36.765 172.395 37.055 172.440 ;
        RECT 37.670 172.380 37.990 172.440 ;
        RECT 47.330 172.580 47.650 172.640 ;
        RECT 48.725 172.580 49.015 172.625 ;
        RECT 61.590 172.580 61.910 172.640 ;
        RECT 64.825 172.580 65.115 172.625 ;
        RECT 47.330 172.440 49.015 172.580 ;
        RECT 47.330 172.380 47.650 172.440 ;
        RECT 48.725 172.395 49.015 172.440 ;
        RECT 52.480 172.440 65.115 172.580 ;
        RECT 52.480 172.300 52.620 172.440 ;
        RECT 61.590 172.380 61.910 172.440 ;
        RECT 64.825 172.395 65.115 172.440 ;
        RECT 65.705 172.580 65.995 172.625 ;
        RECT 66.895 172.580 67.185 172.625 ;
        RECT 69.415 172.580 69.705 172.625 ;
        RECT 83.685 172.580 83.975 172.625 ;
        RECT 65.705 172.440 69.705 172.580 ;
        RECT 65.705 172.395 65.995 172.440 ;
        RECT 66.895 172.395 67.185 172.440 ;
        RECT 69.415 172.395 69.705 172.440 ;
        RECT 81.460 172.440 83.975 172.580 ;
        RECT 81.460 172.300 81.600 172.440 ;
        RECT 83.685 172.395 83.975 172.440 ;
        RECT 33.085 172.100 35.600 172.240 ;
        RECT 24.300 171.900 24.590 171.945 ;
        RECT 30.400 171.900 30.540 172.100 ;
        RECT 33.085 172.055 33.375 172.100 ;
        RECT 38.130 172.040 38.450 172.300 ;
        RECT 39.510 172.240 39.830 172.300 ;
        RECT 40.445 172.240 40.735 172.285 ;
        RECT 39.510 172.100 40.735 172.240 ;
        RECT 39.510 172.040 39.830 172.100 ;
        RECT 40.445 172.055 40.735 172.100 ;
        RECT 41.350 172.240 41.670 172.300 ;
        RECT 42.745 172.240 43.035 172.285 ;
        RECT 41.350 172.100 43.035 172.240 ;
        RECT 41.350 172.040 41.670 172.100 ;
        RECT 42.745 172.055 43.035 172.100 ;
        RECT 47.805 172.240 48.095 172.285 ;
        RECT 48.250 172.240 48.570 172.300 ;
        RECT 47.805 172.100 48.570 172.240 ;
        RECT 47.805 172.055 48.095 172.100 ;
        RECT 48.250 172.040 48.570 172.100 ;
        RECT 52.390 172.040 52.710 172.300 ;
        RECT 58.385 172.240 58.675 172.285 ;
        RECT 58.000 172.100 58.675 172.240 ;
        RECT 24.300 171.760 30.540 171.900 ;
        RECT 31.230 171.900 31.550 171.960 ;
        RECT 31.705 171.900 31.995 171.945 ;
        RECT 33.990 171.900 34.310 171.960 ;
        RECT 31.230 171.760 34.310 171.900 ;
        RECT 24.300 171.715 24.590 171.760 ;
        RECT 31.230 171.700 31.550 171.760 ;
        RECT 31.705 171.715 31.995 171.760 ;
        RECT 33.990 171.700 34.310 171.760 ;
        RECT 34.450 171.900 34.770 171.960 ;
        RECT 34.450 171.760 43.190 171.900 ;
        RECT 34.450 171.700 34.770 171.760 ;
        RECT 32.610 171.360 32.930 171.620 ;
        RECT 39.050 171.560 39.370 171.620 ;
        RECT 39.525 171.560 39.815 171.605 ;
        RECT 39.050 171.420 39.815 171.560 ;
        RECT 39.050 171.360 39.370 171.420 ;
        RECT 39.525 171.375 39.815 171.420 ;
        RECT 39.970 171.360 40.290 171.620 ;
        RECT 43.050 171.560 43.190 171.760 ;
        RECT 58.000 171.620 58.140 172.100 ;
        RECT 58.385 172.055 58.675 172.100 ;
        RECT 59.290 172.040 59.610 172.300 ;
        RECT 59.750 172.040 60.070 172.300 ;
        RECT 60.210 172.240 60.530 172.300 ;
        RECT 60.685 172.240 60.975 172.285 ;
        RECT 60.210 172.100 60.975 172.240 ;
        RECT 60.210 172.040 60.530 172.100 ;
        RECT 60.685 172.055 60.975 172.100 ;
        RECT 60.760 171.900 60.900 172.055 ;
        RECT 61.130 172.040 61.450 172.300 ;
        RECT 66.190 172.285 66.510 172.300 ;
        RECT 63.445 172.240 63.735 172.285 ;
        RECT 61.680 172.100 63.735 172.240 ;
        RECT 61.680 171.900 61.820 172.100 ;
        RECT 63.445 172.055 63.735 172.100 ;
        RECT 63.905 172.055 64.195 172.285 ;
        RECT 66.160 172.240 66.510 172.285 ;
        RECT 65.995 172.100 66.510 172.240 ;
        RECT 66.160 172.055 66.510 172.100 ;
        RECT 60.760 171.760 61.820 171.900 ;
        RECT 62.525 171.900 62.815 171.945 ;
        RECT 62.970 171.900 63.290 171.960 ;
        RECT 63.980 171.900 64.120 172.055 ;
        RECT 66.190 172.040 66.510 172.055 ;
        RECT 78.610 172.040 78.930 172.300 ;
        RECT 81.370 172.040 81.690 172.300 ;
        RECT 84.220 172.285 84.360 172.780 ;
        RECT 82.305 172.055 82.595 172.285 ;
        RECT 83.225 172.055 83.515 172.285 ;
        RECT 84.145 172.055 84.435 172.285 ;
        RECT 62.525 171.760 64.120 171.900 ;
        RECT 78.700 171.900 78.840 172.040 ;
        RECT 82.380 171.900 82.520 172.055 ;
        RECT 78.700 171.760 82.520 171.900 ;
        RECT 83.300 171.900 83.440 172.055 ;
        RECT 86.890 172.040 87.210 172.300 ;
        RECT 86.980 171.900 87.120 172.040 ;
        RECT 83.300 171.760 87.120 171.900 ;
        RECT 62.525 171.715 62.815 171.760 ;
        RECT 62.970 171.700 63.290 171.760 ;
        RECT 43.650 171.560 43.970 171.620 ;
        RECT 43.050 171.420 43.970 171.560 ;
        RECT 43.650 171.360 43.970 171.420 ;
        RECT 56.530 171.560 56.850 171.620 ;
        RECT 57.465 171.560 57.755 171.605 ;
        RECT 56.530 171.420 57.755 171.560 ;
        RECT 56.530 171.360 56.850 171.420 ;
        RECT 57.465 171.375 57.755 171.420 ;
        RECT 57.910 171.360 58.230 171.620 ;
        RECT 60.670 171.560 60.990 171.620 ;
        RECT 61.605 171.560 61.895 171.605 ;
        RECT 60.670 171.420 61.895 171.560 ;
        RECT 60.670 171.360 60.990 171.420 ;
        RECT 61.605 171.375 61.895 171.420 ;
        RECT 75.390 171.560 75.710 171.620 ;
        RECT 85.050 171.560 85.370 171.620 ;
        RECT 75.390 171.420 85.370 171.560 ;
        RECT 75.390 171.360 75.710 171.420 ;
        RECT 85.050 171.360 85.370 171.420 ;
        RECT 18.280 170.740 93.120 171.220 ;
        RECT 25.250 170.340 25.570 170.600 ;
        RECT 28.025 170.540 28.315 170.585 ;
        RECT 32.610 170.540 32.930 170.600 ;
        RECT 28.025 170.400 32.930 170.540 ;
        RECT 28.025 170.355 28.315 170.400 ;
        RECT 32.610 170.340 32.930 170.400 ;
        RECT 59.305 170.540 59.595 170.585 ;
        RECT 62.970 170.540 63.290 170.600 ;
        RECT 59.305 170.400 63.290 170.540 ;
        RECT 59.305 170.355 59.595 170.400 ;
        RECT 62.970 170.340 63.290 170.400 ;
        RECT 66.650 170.340 66.970 170.600 ;
        RECT 67.570 170.540 67.890 170.600 ;
        RECT 67.570 170.400 82.520 170.540 ;
        RECT 67.570 170.340 67.890 170.400 ;
        RECT 25.340 169.860 25.480 170.340 ;
        RECT 29.390 170.200 29.710 170.260 ;
        RECT 28.100 170.060 29.710 170.200 ;
        RECT 28.100 169.905 28.240 170.060 ;
        RECT 29.390 170.000 29.710 170.060 ;
        RECT 37.225 170.200 37.515 170.245 ;
        RECT 40.430 170.200 40.750 170.260 ;
        RECT 37.225 170.060 40.750 170.200 ;
        RECT 37.225 170.015 37.515 170.060 ;
        RECT 40.430 170.000 40.750 170.060 ;
        RECT 43.650 170.200 43.970 170.260 ;
        RECT 43.650 170.060 60.900 170.200 ;
        RECT 43.650 170.000 43.970 170.060 ;
        RECT 60.760 169.920 60.900 170.060 ;
        RECT 27.105 169.860 27.395 169.905 ;
        RECT 25.340 169.720 27.395 169.860 ;
        RECT 27.105 169.675 27.395 169.720 ;
        RECT 28.025 169.675 28.315 169.905 ;
        RECT 39.050 169.660 39.370 169.920 ;
        RECT 52.390 169.660 52.710 169.920 ;
        RECT 53.770 169.905 54.090 169.920 ;
        RECT 53.740 169.675 54.090 169.905 ;
        RECT 53.770 169.660 54.090 169.675 ;
        RECT 58.370 169.860 58.690 169.920 ;
        RECT 59.765 169.860 60.055 169.905 ;
        RECT 58.370 169.720 60.055 169.860 ;
        RECT 58.370 169.660 58.690 169.720 ;
        RECT 59.765 169.675 60.055 169.720 ;
        RECT 60.670 169.860 60.990 169.920 ;
        RECT 66.740 169.860 66.880 170.340 ;
        RECT 75.850 170.000 76.170 170.260 ;
        RECT 78.610 170.200 78.930 170.260 ;
        RECT 78.610 170.060 80.220 170.200 ;
        RECT 78.610 170.000 78.930 170.060 ;
        RECT 60.670 169.720 66.880 169.860 ;
        RECT 68.490 169.860 68.810 169.920 ;
        RECT 72.170 169.860 72.490 169.920 ;
        RECT 75.390 169.860 75.710 169.920 ;
        RECT 68.490 169.720 75.710 169.860 ;
        RECT 75.940 169.860 76.080 170.000 ;
        RECT 78.150 169.860 78.470 169.920 ;
        RECT 80.080 169.905 80.220 170.060 ;
        RECT 81.370 170.000 81.690 170.260 ;
        RECT 80.910 169.905 81.230 169.920 ;
        RECT 82.380 169.905 82.520 170.400 ;
        RECT 79.545 169.860 79.835 169.905 ;
        RECT 75.940 169.720 77.460 169.860 ;
        RECT 60.670 169.660 60.990 169.720 ;
        RECT 68.490 169.660 68.810 169.720 ;
        RECT 72.170 169.660 72.490 169.720 ;
        RECT 75.390 169.660 75.710 169.720 ;
        RECT 35.830 169.520 36.150 169.580 ;
        RECT 38.145 169.520 38.435 169.565 ;
        RECT 35.830 169.380 38.435 169.520 ;
        RECT 35.830 169.320 36.150 169.380 ;
        RECT 38.145 169.335 38.435 169.380 ;
        RECT 38.590 169.320 38.910 169.580 ;
        RECT 39.525 169.520 39.815 169.565 ;
        RECT 39.970 169.520 40.290 169.580 ;
        RECT 39.525 169.380 40.290 169.520 ;
        RECT 39.525 169.335 39.815 169.380 ;
        RECT 39.970 169.320 40.290 169.380 ;
        RECT 53.285 169.520 53.575 169.565 ;
        RECT 54.475 169.520 54.765 169.565 ;
        RECT 56.995 169.520 57.285 169.565 ;
        RECT 53.285 169.380 57.285 169.520 ;
        RECT 53.285 169.335 53.575 169.380 ;
        RECT 54.475 169.335 54.765 169.380 ;
        RECT 56.995 169.335 57.285 169.380 ;
        RECT 74.930 169.320 75.250 169.580 ;
        RECT 75.865 169.335 76.155 169.565 ;
        RECT 76.325 169.335 76.615 169.565 ;
        RECT 77.320 169.520 77.460 169.720 ;
        RECT 78.150 169.720 79.835 169.860 ;
        RECT 78.150 169.660 78.470 169.720 ;
        RECT 79.545 169.675 79.835 169.720 ;
        RECT 80.005 169.675 80.295 169.905 ;
        RECT 80.745 169.675 81.230 169.905 ;
        RECT 81.845 169.675 82.135 169.905 ;
        RECT 82.330 169.675 82.620 169.905 ;
        RECT 80.910 169.660 81.230 169.675 ;
        RECT 79.070 169.520 79.390 169.580 ;
        RECT 81.920 169.520 82.060 169.675 ;
        RECT 77.320 169.380 79.390 169.520 ;
        RECT 28.930 169.180 29.250 169.240 ;
        RECT 30.785 169.180 31.075 169.225 ;
        RECT 32.150 169.180 32.470 169.240 ;
        RECT 44.570 169.180 44.890 169.240 ;
        RECT 28.930 169.040 44.890 169.180 ;
        RECT 28.930 168.980 29.250 169.040 ;
        RECT 30.785 168.995 31.075 169.040 ;
        RECT 32.150 168.980 32.470 169.040 ;
        RECT 44.570 168.980 44.890 169.040 ;
        RECT 52.890 169.180 53.180 169.225 ;
        RECT 54.990 169.180 55.280 169.225 ;
        RECT 56.560 169.180 56.850 169.225 ;
        RECT 52.890 169.040 56.850 169.180 ;
        RECT 52.890 168.995 53.180 169.040 ;
        RECT 54.990 168.995 55.280 169.040 ;
        RECT 56.560 168.995 56.850 169.040 ;
        RECT 60.225 169.180 60.515 169.225 ;
        RECT 75.940 169.180 76.080 169.335 ;
        RECT 60.225 169.040 76.080 169.180 ;
        RECT 76.400 169.180 76.540 169.335 ;
        RECT 79.070 169.320 79.390 169.380 ;
        RECT 79.620 169.380 82.060 169.520 ;
        RECT 79.620 169.240 79.760 169.380 ;
        RECT 77.705 169.180 77.995 169.225 ;
        RECT 76.400 169.040 77.995 169.180 ;
        RECT 60.225 168.995 60.515 169.040 ;
        RECT 77.705 168.995 77.995 169.040 ;
        RECT 79.530 168.980 79.850 169.240 ;
        RECT 38.130 168.840 38.450 168.900 ;
        RECT 40.445 168.840 40.735 168.885 ;
        RECT 38.130 168.700 40.735 168.840 ;
        RECT 38.130 168.640 38.450 168.700 ;
        RECT 40.445 168.655 40.735 168.700 ;
        RECT 62.050 168.840 62.370 168.900 ;
        RECT 66.650 168.840 66.970 168.900 ;
        RECT 62.050 168.700 66.970 168.840 ;
        RECT 62.050 168.640 62.370 168.700 ;
        RECT 66.650 168.640 66.970 168.700 ;
        RECT 77.230 168.640 77.550 168.900 ;
        RECT 78.610 168.640 78.930 168.900 ;
        RECT 83.225 168.840 83.515 168.885 ;
        RECT 85.510 168.840 85.830 168.900 ;
        RECT 83.225 168.700 85.830 168.840 ;
        RECT 83.225 168.655 83.515 168.700 ;
        RECT 85.510 168.640 85.830 168.700 ;
        RECT 18.280 168.020 92.340 168.500 ;
        RECT 37.225 167.820 37.515 167.865 ;
        RECT 37.670 167.820 37.990 167.880 ;
        RECT 37.225 167.680 37.990 167.820 ;
        RECT 37.225 167.635 37.515 167.680 ;
        RECT 37.670 167.620 37.990 167.680 ;
        RECT 39.510 167.620 39.830 167.880 ;
        RECT 53.770 167.820 54.090 167.880 ;
        RECT 54.705 167.820 54.995 167.865 ;
        RECT 70.330 167.820 70.650 167.880 ;
        RECT 72.645 167.820 72.935 167.865 ;
        RECT 53.770 167.680 54.995 167.820 ;
        RECT 53.770 167.620 54.090 167.680 ;
        RECT 54.705 167.635 54.995 167.680 ;
        RECT 63.520 167.680 72.935 167.820 ;
        RECT 29.850 167.480 30.170 167.540 ;
        RECT 34.465 167.480 34.755 167.525 ;
        RECT 29.850 167.340 34.755 167.480 ;
        RECT 29.850 167.280 30.170 167.340 ;
        RECT 34.465 167.295 34.755 167.340 ;
        RECT 40.930 167.480 41.220 167.525 ;
        RECT 43.030 167.480 43.320 167.525 ;
        RECT 44.600 167.480 44.890 167.525 ;
        RECT 40.930 167.340 44.890 167.480 ;
        RECT 40.930 167.295 41.220 167.340 ;
        RECT 43.030 167.295 43.320 167.340 ;
        RECT 44.600 167.295 44.890 167.340 ;
        RECT 47.330 167.480 47.650 167.540 ;
        RECT 47.330 167.340 49.860 167.480 ;
        RECT 34.540 167.140 34.680 167.295 ;
        RECT 47.330 167.280 47.650 167.340 ;
        RECT 35.830 167.140 36.150 167.200 ;
        RECT 49.720 167.185 49.860 167.340 ;
        RECT 37.685 167.140 37.975 167.185 ;
        RECT 34.540 167.000 37.975 167.140 ;
        RECT 35.830 166.940 36.150 167.000 ;
        RECT 37.685 166.955 37.975 167.000 ;
        RECT 41.325 167.140 41.615 167.185 ;
        RECT 42.515 167.140 42.805 167.185 ;
        RECT 45.035 167.140 45.325 167.185 ;
        RECT 41.325 167.000 45.325 167.140 ;
        RECT 41.325 166.955 41.615 167.000 ;
        RECT 42.515 166.955 42.805 167.000 ;
        RECT 45.035 166.955 45.325 167.000 ;
        RECT 49.645 166.955 49.935 167.185 ;
        RECT 52.865 167.140 53.155 167.185 ;
        RECT 63.520 167.140 63.660 167.680 ;
        RECT 70.330 167.620 70.650 167.680 ;
        RECT 72.645 167.635 72.935 167.680 ;
        RECT 76.325 167.820 76.615 167.865 ;
        RECT 76.770 167.820 77.090 167.880 ;
        RECT 76.325 167.680 77.090 167.820 ;
        RECT 76.325 167.635 76.615 167.680 ;
        RECT 76.770 167.620 77.090 167.680 ;
        RECT 80.910 167.820 81.230 167.880 ;
        RECT 81.845 167.820 82.135 167.865 ;
        RECT 80.910 167.680 82.135 167.820 ;
        RECT 80.910 167.620 81.230 167.680 ;
        RECT 81.845 167.635 82.135 167.680 ;
        RECT 63.905 167.480 64.195 167.525 ;
        RECT 64.825 167.480 65.115 167.525 ;
        RECT 63.905 167.340 65.115 167.480 ;
        RECT 63.905 167.295 64.195 167.340 ;
        RECT 64.825 167.295 65.115 167.340 ;
        RECT 52.865 167.000 55.380 167.140 ;
        RECT 63.520 167.000 64.120 167.140 ;
        RECT 52.865 166.955 53.155 167.000 ;
        RECT 38.590 166.800 38.910 166.860 ;
        RECT 35.460 166.660 38.910 166.800 ;
        RECT 29.850 166.120 30.170 166.180 ;
        RECT 34.910 166.120 35.230 166.180 ;
        RECT 35.460 166.165 35.600 166.660 ;
        RECT 38.590 166.600 38.910 166.660 ;
        RECT 39.050 166.600 39.370 166.860 ;
        RECT 40.445 166.800 40.735 166.845 ;
        RECT 44.570 166.800 44.890 166.860 ;
        RECT 40.445 166.660 44.890 166.800 ;
        RECT 40.445 166.615 40.735 166.660 ;
        RECT 44.570 166.600 44.890 166.660 ;
        RECT 53.785 166.800 54.075 166.845 ;
        RECT 54.230 166.800 54.550 166.860 ;
        RECT 55.240 166.845 55.380 167.000 ;
        RECT 53.785 166.660 54.550 166.800 ;
        RECT 53.785 166.615 54.075 166.660 ;
        RECT 35.845 166.460 36.135 166.505 ;
        RECT 39.140 166.460 39.280 166.600 ;
        RECT 35.845 166.320 39.280 166.460 ;
        RECT 41.780 166.460 42.070 166.505 ;
        RECT 42.270 166.460 42.590 166.520 ;
        RECT 41.780 166.320 42.590 166.460 ;
        RECT 35.845 166.275 36.135 166.320 ;
        RECT 41.780 166.275 42.070 166.320 ;
        RECT 42.270 166.260 42.590 166.320 ;
        RECT 52.850 166.460 53.170 166.520 ;
        RECT 53.860 166.460 54.000 166.615 ;
        RECT 54.230 166.600 54.550 166.660 ;
        RECT 54.705 166.615 54.995 166.845 ;
        RECT 55.165 166.615 55.455 166.845 ;
        RECT 52.850 166.320 54.000 166.460 ;
        RECT 54.780 166.460 54.920 166.615 ;
        RECT 56.530 166.600 56.850 166.860 ;
        RECT 62.510 166.600 62.830 166.860 ;
        RECT 63.980 166.845 64.120 167.000 ;
        RECT 63.905 166.615 64.195 166.845 ;
        RECT 64.365 166.615 64.655 166.845 ;
        RECT 64.900 166.800 65.040 167.295 ;
        RECT 66.190 167.280 66.510 167.540 ;
        RECT 66.650 167.280 66.970 167.540 ;
        RECT 76.860 167.480 77.000 167.620 ;
        RECT 71.340 167.340 74.240 167.480 ;
        RECT 76.860 167.340 78.840 167.480 ;
        RECT 65.745 167.140 66.035 167.185 ;
        RECT 66.740 167.140 66.880 167.280 ;
        RECT 65.745 167.000 66.880 167.140 ;
        RECT 65.745 166.955 66.035 167.000 ;
        RECT 67.585 166.800 67.875 166.845 ;
        RECT 64.900 166.660 67.875 166.800 ;
        RECT 67.585 166.615 67.875 166.660 ;
        RECT 68.030 166.800 68.350 166.860 ;
        RECT 71.340 166.845 71.480 167.340 ;
        RECT 70.345 166.800 70.635 166.845 ;
        RECT 68.030 166.660 70.635 166.800 ;
        RECT 56.620 166.460 56.760 166.600 ;
        RECT 54.780 166.320 56.760 166.460 ;
        RECT 52.850 166.260 53.170 166.320 ;
        RECT 35.385 166.120 35.675 166.165 ;
        RECT 29.850 165.980 35.675 166.120 ;
        RECT 29.850 165.920 30.170 165.980 ;
        RECT 34.910 165.920 35.230 165.980 ;
        RECT 35.385 165.935 35.675 165.980 ;
        RECT 36.305 166.120 36.595 166.165 ;
        RECT 38.130 166.120 38.450 166.180 ;
        RECT 39.970 166.120 40.290 166.180 ;
        RECT 36.305 165.980 40.290 166.120 ;
        RECT 36.305 165.935 36.595 165.980 ;
        RECT 38.130 165.920 38.450 165.980 ;
        RECT 39.970 165.920 40.290 165.980 ;
        RECT 53.310 166.120 53.630 166.180 ;
        RECT 55.625 166.120 55.915 166.165 ;
        RECT 53.310 165.980 55.915 166.120 ;
        RECT 53.310 165.920 53.630 165.980 ;
        RECT 55.625 165.935 55.915 165.980 ;
        RECT 62.970 165.920 63.290 166.180 ;
        RECT 64.440 166.120 64.580 166.615 ;
        RECT 68.030 166.600 68.350 166.660 ;
        RECT 70.345 166.615 70.635 166.660 ;
        RECT 71.265 166.615 71.555 166.845 ;
        RECT 72.185 166.800 72.475 166.845 ;
        RECT 72.630 166.800 72.950 166.860 ;
        RECT 72.185 166.660 72.950 166.800 ;
        RECT 72.185 166.615 72.475 166.660 ;
        RECT 72.630 166.600 72.950 166.660 ;
        RECT 73.565 166.615 73.855 166.845 ;
        RECT 74.100 166.800 74.240 167.340 ;
        RECT 78.165 167.140 78.455 167.185 ;
        RECT 75.940 167.000 78.455 167.140 ;
        RECT 75.940 166.800 76.080 167.000 ;
        RECT 78.165 166.955 78.455 167.000 ;
        RECT 74.100 166.660 76.080 166.800 ;
        RECT 76.785 166.800 77.075 166.845 ;
        RECT 76.785 166.660 77.460 166.800 ;
        RECT 76.785 166.615 77.075 166.660 ;
        RECT 65.745 166.460 66.035 166.505 ;
        RECT 66.205 166.460 66.495 166.505 ;
        RECT 65.745 166.320 66.495 166.460 ;
        RECT 65.745 166.275 66.035 166.320 ;
        RECT 66.205 166.275 66.495 166.320 ;
        RECT 67.125 166.460 67.415 166.505 ;
        RECT 68.490 166.460 68.810 166.520 ;
        RECT 67.125 166.320 68.810 166.460 ;
        RECT 67.125 166.275 67.415 166.320 ;
        RECT 67.200 166.120 67.340 166.275 ;
        RECT 68.490 166.260 68.810 166.320 ;
        RECT 70.790 166.460 71.110 166.520 ;
        RECT 73.640 166.460 73.780 166.615 ;
        RECT 70.790 166.320 77.000 166.460 ;
        RECT 70.790 166.260 71.110 166.320 ;
        RECT 76.860 166.180 77.000 166.320 ;
        RECT 64.440 165.980 67.340 166.120 ;
        RECT 69.425 166.120 69.715 166.165 ;
        RECT 71.710 166.120 72.030 166.180 ;
        RECT 69.425 165.980 72.030 166.120 ;
        RECT 69.425 165.935 69.715 165.980 ;
        RECT 71.710 165.920 72.030 165.980 ;
        RECT 76.770 165.920 77.090 166.180 ;
        RECT 77.320 166.120 77.460 166.660 ;
        RECT 77.690 166.600 78.010 166.860 ;
        RECT 78.700 166.845 78.840 167.340 ;
        RECT 84.680 167.000 90.800 167.140 ;
        RECT 84.680 166.845 84.820 167.000 ;
        RECT 90.660 166.860 90.800 167.000 ;
        RECT 78.625 166.615 78.915 166.845 ;
        RECT 80.925 166.800 81.215 166.845 ;
        RECT 84.605 166.800 84.895 166.845 ;
        RECT 80.925 166.660 84.895 166.800 ;
        RECT 80.925 166.615 81.215 166.660 ;
        RECT 84.605 166.615 84.895 166.660 ;
        RECT 85.050 166.600 85.370 166.860 ;
        RECT 85.510 166.600 85.830 166.860 ;
        RECT 86.430 166.600 86.750 166.860 ;
        RECT 90.570 166.600 90.890 166.860 ;
        RECT 78.150 166.460 78.470 166.520 ;
        RECT 80.005 166.460 80.295 166.505 ;
        RECT 78.150 166.320 80.295 166.460 ;
        RECT 78.150 166.260 78.470 166.320 ;
        RECT 80.005 166.275 80.295 166.320 ;
        RECT 79.070 166.120 79.390 166.180 ;
        RECT 77.320 165.980 79.390 166.120 ;
        RECT 79.070 165.920 79.390 165.980 ;
        RECT 83.225 166.120 83.515 166.165 ;
        RECT 83.670 166.120 83.990 166.180 ;
        RECT 83.225 165.980 83.990 166.120 ;
        RECT 83.225 165.935 83.515 165.980 ;
        RECT 83.670 165.920 83.990 165.980 ;
        RECT 18.280 165.300 93.120 165.780 ;
        RECT 30.325 165.100 30.615 165.145 ;
        RECT 29.940 164.960 30.615 165.100 ;
        RECT 29.940 164.820 30.080 164.960 ;
        RECT 30.325 164.915 30.615 164.960 ;
        RECT 33.530 165.100 33.850 165.160 ;
        RECT 33.530 164.960 39.740 165.100 ;
        RECT 33.530 164.900 33.850 164.960 ;
        RECT 29.850 164.560 30.170 164.820 ;
        RECT 39.050 164.760 39.370 164.820 ;
        RECT 36.380 164.620 39.370 164.760 ;
        RECT 29.390 164.420 29.710 164.480 ;
        RECT 30.310 164.420 30.600 164.465 ;
        RECT 34.450 164.420 34.770 164.480 ;
        RECT 29.390 164.280 34.770 164.420 ;
        RECT 29.390 164.220 29.710 164.280 ;
        RECT 30.310 164.235 30.600 164.280 ;
        RECT 34.450 164.220 34.770 164.280 ;
        RECT 34.910 164.465 35.230 164.480 ;
        RECT 36.380 164.465 36.520 164.620 ;
        RECT 39.050 164.560 39.370 164.620 ;
        RECT 34.910 164.420 35.250 164.465 ;
        RECT 34.910 164.280 35.405 164.420 ;
        RECT 34.910 164.235 35.250 164.280 ;
        RECT 36.305 164.235 36.595 164.465 ;
        RECT 37.225 164.420 37.515 164.465 ;
        RECT 39.600 164.420 39.740 164.960 ;
        RECT 42.270 164.900 42.590 165.160 ;
        RECT 53.310 164.900 53.630 165.160 ;
        RECT 53.770 165.100 54.090 165.160 ;
        RECT 62.970 165.100 63.290 165.160 ;
        RECT 70.790 165.100 71.110 165.160 ;
        RECT 53.770 164.960 71.110 165.100 ;
        RECT 53.770 164.900 54.090 164.960 ;
        RECT 62.970 164.900 63.290 164.960 ;
        RECT 70.790 164.900 71.110 164.960 ;
        RECT 75.865 165.100 76.155 165.145 ;
        RECT 77.690 165.100 78.010 165.160 ;
        RECT 75.865 164.960 78.010 165.100 ;
        RECT 75.865 164.915 76.155 164.960 ;
        RECT 77.690 164.900 78.010 164.960 ;
        RECT 78.150 164.900 78.470 165.160 ;
        RECT 80.080 164.960 88.040 165.100 ;
        RECT 41.825 164.420 42.115 164.465 ;
        RECT 37.225 164.280 38.360 164.420 ;
        RECT 39.600 164.280 42.115 164.420 ;
        RECT 37.225 164.235 37.515 164.280 ;
        RECT 34.910 164.220 35.230 164.235 ;
        RECT 38.220 164.140 38.360 164.280 ;
        RECT 41.825 164.235 42.115 164.280 ;
        RECT 42.745 164.235 43.035 164.465 ;
        RECT 44.570 164.420 44.890 164.480 ;
        RECT 46.425 164.420 46.715 164.465 ;
        RECT 44.570 164.280 46.715 164.420 ;
        RECT 32.625 163.895 32.915 164.125 ;
        RECT 35.385 164.080 35.675 164.125 ;
        RECT 35.385 163.940 36.980 164.080 ;
        RECT 35.385 163.895 35.675 163.940 ;
        RECT 32.700 163.740 32.840 163.895 ;
        RECT 32.700 163.600 36.520 163.740 ;
        RECT 36.380 163.460 36.520 163.600 ;
        RECT 29.390 163.200 29.710 163.460 ;
        RECT 32.165 163.400 32.455 163.445 ;
        RECT 33.085 163.400 33.375 163.445 ;
        RECT 32.165 163.260 33.375 163.400 ;
        RECT 32.165 163.215 32.455 163.260 ;
        RECT 33.085 163.215 33.375 163.260 ;
        RECT 36.290 163.200 36.610 163.460 ;
        RECT 36.840 163.445 36.980 163.940 ;
        RECT 38.130 163.880 38.450 164.140 ;
        RECT 42.820 163.740 42.960 164.235 ;
        RECT 44.570 164.220 44.890 164.280 ;
        RECT 46.425 164.235 46.715 164.280 ;
        RECT 47.330 164.220 47.650 164.480 ;
        RECT 48.710 164.420 49.030 164.480 ;
        RECT 51.025 164.420 51.315 164.465 ;
        RECT 53.400 164.420 53.540 164.900 ;
        RECT 72.630 164.760 72.950 164.820 ;
        RECT 80.080 164.805 80.220 164.960 ;
        RECT 87.900 164.820 88.040 164.960 ;
        RECT 78.925 164.760 79.215 164.805 ;
        RECT 72.630 164.620 79.215 164.760 ;
        RECT 72.630 164.560 72.950 164.620 ;
        RECT 48.710 164.280 50.780 164.420 ;
        RECT 48.710 164.220 49.030 164.280 ;
        RECT 46.885 164.080 47.175 164.125 ;
        RECT 49.645 164.080 49.935 164.125 ;
        RECT 46.885 163.940 49.935 164.080 ;
        RECT 46.885 163.895 47.175 163.940 ;
        RECT 49.645 163.895 49.935 163.940 ;
        RECT 50.105 163.895 50.395 164.125 ;
        RECT 50.640 164.080 50.780 164.280 ;
        RECT 51.025 164.280 53.540 164.420 ;
        RECT 51.025 164.235 51.315 164.280 ;
        RECT 57.910 164.220 58.230 164.480 ;
        RECT 75.480 164.465 75.620 164.620 ;
        RECT 78.925 164.575 79.215 164.620 ;
        RECT 80.005 164.575 80.295 164.805 ;
        RECT 83.230 164.760 83.520 164.805 ;
        RECT 84.630 164.760 84.920 164.805 ;
        RECT 86.470 164.760 86.760 164.805 ;
        RECT 83.230 164.620 86.760 164.760 ;
        RECT 83.230 164.575 83.520 164.620 ;
        RECT 84.630 164.575 84.920 164.620 ;
        RECT 86.470 164.575 86.760 164.620 ;
        RECT 75.405 164.420 75.695 164.465 ;
        RECT 75.195 164.280 75.695 164.420 ;
        RECT 75.405 164.235 75.695 164.280 ;
        RECT 76.785 164.420 77.075 164.465 ;
        RECT 80.080 164.420 80.220 164.575 ;
        RECT 87.810 164.560 88.130 164.820 ;
        RECT 76.785 164.280 80.220 164.420 ;
        RECT 80.450 164.420 80.770 164.480 ;
        RECT 82.305 164.420 82.595 164.465 ;
        RECT 80.450 164.280 82.595 164.420 ;
        RECT 76.785 164.235 77.075 164.280 ;
        RECT 58.000 164.080 58.140 164.220 ;
        RECT 50.640 163.940 58.140 164.080 ;
        RECT 75.480 164.080 75.620 164.235 ;
        RECT 80.450 164.220 80.770 164.280 ;
        RECT 82.305 164.235 82.595 164.280 ;
        RECT 83.670 164.220 83.990 164.480 ;
        RECT 90.570 164.220 90.890 164.480 ;
        RECT 75.480 163.940 79.760 164.080 ;
        RECT 47.805 163.740 48.095 163.785 ;
        RECT 42.820 163.600 48.095 163.740 ;
        RECT 47.805 163.555 48.095 163.600 ;
        RECT 49.170 163.540 49.490 163.800 ;
        RECT 50.180 163.740 50.320 163.895 ;
        RECT 59.750 163.740 60.070 163.800 ;
        RECT 50.180 163.600 60.070 163.740 ;
        RECT 36.765 163.400 37.055 163.445 ;
        RECT 37.670 163.400 37.990 163.460 ;
        RECT 36.765 163.260 37.990 163.400 ;
        RECT 36.765 163.215 37.055 163.260 ;
        RECT 37.670 163.200 37.990 163.260 ;
        RECT 44.110 163.400 44.430 163.460 ;
        RECT 46.870 163.400 47.190 163.460 ;
        RECT 50.180 163.400 50.320 163.600 ;
        RECT 59.750 163.540 60.070 163.600 ;
        RECT 76.785 163.740 77.075 163.785 ;
        RECT 78.610 163.740 78.930 163.800 ;
        RECT 76.785 163.600 78.930 163.740 ;
        RECT 76.785 163.555 77.075 163.600 ;
        RECT 78.610 163.540 78.930 163.600 ;
        RECT 79.620 163.460 79.760 163.940 ;
        RECT 82.770 163.740 83.060 163.785 ;
        RECT 85.090 163.740 85.380 163.785 ;
        RECT 86.470 163.740 86.760 163.785 ;
        RECT 82.770 163.600 86.760 163.740 ;
        RECT 82.770 163.555 83.060 163.600 ;
        RECT 85.090 163.555 85.380 163.600 ;
        RECT 86.470 163.555 86.760 163.600 ;
        RECT 44.110 163.260 50.320 163.400 ;
        RECT 44.110 163.200 44.430 163.260 ;
        RECT 46.870 163.200 47.190 163.260 ;
        RECT 79.070 163.200 79.390 163.460 ;
        RECT 79.530 163.200 79.850 163.460 ;
        RECT 18.280 162.580 92.340 163.060 ;
        RECT 29.390 162.180 29.710 162.440 ;
        RECT 36.290 162.380 36.610 162.440 ;
        RECT 37.225 162.380 37.515 162.425 ;
        RECT 36.290 162.240 37.515 162.380 ;
        RECT 36.290 162.180 36.610 162.240 ;
        RECT 37.225 162.195 37.515 162.240 ;
        RECT 38.130 162.380 38.450 162.440 ;
        RECT 49.170 162.380 49.490 162.440 ;
        RECT 50.565 162.380 50.855 162.425 ;
        RECT 38.130 162.240 50.855 162.380 ;
        RECT 22.990 162.040 23.280 162.085 ;
        RECT 25.090 162.040 25.380 162.085 ;
        RECT 26.660 162.040 26.950 162.085 ;
        RECT 22.990 161.900 26.950 162.040 ;
        RECT 22.990 161.855 23.280 161.900 ;
        RECT 25.090 161.855 25.380 161.900 ;
        RECT 26.660 161.855 26.950 161.900 ;
        RECT 22.490 161.500 22.810 161.760 ;
        RECT 23.385 161.700 23.675 161.745 ;
        RECT 24.575 161.700 24.865 161.745 ;
        RECT 27.095 161.700 27.385 161.745 ;
        RECT 23.385 161.560 27.385 161.700 ;
        RECT 23.385 161.515 23.675 161.560 ;
        RECT 24.575 161.515 24.865 161.560 ;
        RECT 27.095 161.515 27.385 161.560 ;
        RECT 29.480 161.360 29.620 162.180 ;
        RECT 37.300 162.040 37.440 162.195 ;
        RECT 38.130 162.180 38.450 162.240 ;
        RECT 49.170 162.180 49.490 162.240 ;
        RECT 50.565 162.195 50.855 162.240 ;
        RECT 63.905 162.380 64.195 162.425 ;
        RECT 65.730 162.380 66.050 162.440 ;
        RECT 63.905 162.240 66.050 162.380 ;
        RECT 63.905 162.195 64.195 162.240 ;
        RECT 65.730 162.180 66.050 162.240 ;
        RECT 70.330 162.180 70.650 162.440 ;
        RECT 86.890 162.180 87.210 162.440 ;
        RECT 43.190 162.040 43.510 162.100 ;
        RECT 37.300 161.900 43.510 162.040 ;
        RECT 43.050 161.840 43.510 161.900 ;
        RECT 47.330 162.040 47.650 162.100 ;
        RECT 47.805 162.040 48.095 162.085 ;
        RECT 47.330 161.900 48.095 162.040 ;
        RECT 47.330 161.840 47.650 161.900 ;
        RECT 47.805 161.855 48.095 161.900 ;
        RECT 48.710 161.840 49.030 162.100 ;
        RECT 56.085 162.040 56.375 162.085 ;
        RECT 57.925 162.040 58.215 162.085 ;
        RECT 56.085 161.900 58.215 162.040 ;
        RECT 56.085 161.855 56.375 161.900 ;
        RECT 57.925 161.855 58.215 161.900 ;
        RECT 64.350 162.040 64.670 162.100 ;
        RECT 64.825 162.040 65.115 162.085 ;
        RECT 64.350 161.900 65.115 162.040 ;
        RECT 64.350 161.840 64.670 161.900 ;
        RECT 64.825 161.855 65.115 161.900 ;
        RECT 36.305 161.700 36.595 161.745 ;
        RECT 38.605 161.700 38.895 161.745 ;
        RECT 36.305 161.560 38.895 161.700 ;
        RECT 43.050 161.700 43.190 161.840 ;
        RECT 48.800 161.700 48.940 161.840 ;
        RECT 43.050 161.560 48.940 161.700 ;
        RECT 54.690 161.700 55.010 161.760 ;
        RECT 65.820 161.700 65.960 162.180 ;
        RECT 66.650 162.040 66.970 162.100 ;
        RECT 75.850 162.040 76.170 162.100 ;
        RECT 66.650 161.900 76.170 162.040 ;
        RECT 66.650 161.840 66.970 161.900 ;
        RECT 75.850 161.840 76.170 161.900 ;
        RECT 77.690 161.840 78.010 162.100 ;
        RECT 89.665 162.040 89.955 162.085 ;
        RECT 90.570 162.040 90.890 162.100 ;
        RECT 89.665 161.900 90.890 162.040 ;
        RECT 89.665 161.855 89.955 161.900 ;
        RECT 90.570 161.840 90.890 161.900 ;
        RECT 71.265 161.700 71.555 161.745 ;
        RECT 77.780 161.700 77.920 161.840 ;
        RECT 54.690 161.560 62.740 161.700 ;
        RECT 65.820 161.560 70.100 161.700 ;
        RECT 36.305 161.515 36.595 161.560 ;
        RECT 38.605 161.515 38.895 161.560 ;
        RECT 29.865 161.360 30.155 161.405 ;
        RECT 29.480 161.220 30.155 161.360 ;
        RECT 29.865 161.175 30.155 161.220 ;
        RECT 30.785 161.360 31.075 161.405 ;
        RECT 33.530 161.360 33.850 161.420 ;
        RECT 30.785 161.220 33.850 161.360 ;
        RECT 30.785 161.175 31.075 161.220 ;
        RECT 33.530 161.160 33.850 161.220 ;
        RECT 37.670 161.160 37.990 161.420 ;
        RECT 38.130 161.160 38.450 161.420 ;
        RECT 39.050 161.160 39.370 161.420 ;
        RECT 45.120 161.405 45.260 161.560 ;
        RECT 54.690 161.500 55.010 161.560 ;
        RECT 45.045 161.175 45.335 161.405 ;
        RECT 45.490 161.160 45.810 161.420 ;
        RECT 45.950 161.160 46.270 161.420 ;
        RECT 46.425 161.360 46.715 161.405 ;
        RECT 46.870 161.360 47.190 161.420 ;
        RECT 46.425 161.220 47.190 161.360 ;
        RECT 46.425 161.175 46.715 161.220 ;
        RECT 46.870 161.160 47.190 161.220 ;
        RECT 47.345 161.360 47.635 161.405 ;
        RECT 51.945 161.360 52.235 161.405 ;
        RECT 47.345 161.220 52.235 161.360 ;
        RECT 47.345 161.175 47.635 161.220 ;
        RECT 51.945 161.175 52.235 161.220 ;
        RECT 52.390 161.160 52.710 161.420 ;
        RECT 54.245 161.175 54.535 161.405 ;
        RECT 57.465 161.360 57.755 161.405 ;
        RECT 57.910 161.360 58.230 161.420 ;
        RECT 57.465 161.220 58.230 161.360 ;
        RECT 57.465 161.175 57.755 161.220 ;
        RECT 23.840 161.020 24.130 161.065 ;
        RECT 30.325 161.020 30.615 161.065 ;
        RECT 23.840 160.880 30.615 161.020 ;
        RECT 23.840 160.835 24.130 160.880 ;
        RECT 30.325 160.835 30.615 160.880 ;
        RECT 49.170 161.020 49.490 161.080 ;
        RECT 54.320 161.020 54.460 161.175 ;
        RECT 57.910 161.160 58.230 161.220 ;
        RECT 60.060 161.360 60.350 161.405 ;
        RECT 60.670 161.360 60.990 161.420 ;
        RECT 60.060 161.220 60.990 161.360 ;
        RECT 60.060 161.175 60.350 161.220 ;
        RECT 60.670 161.160 60.990 161.220 ;
        RECT 49.170 160.880 59.980 161.020 ;
        RECT 49.170 160.820 49.490 160.880 ;
        RECT 29.405 160.680 29.695 160.725 ;
        RECT 29.850 160.680 30.170 160.740 ;
        RECT 29.405 160.540 30.170 160.680 ;
        RECT 29.405 160.495 29.695 160.540 ;
        RECT 29.850 160.480 30.170 160.540 ;
        RECT 34.910 160.480 35.230 160.740 ;
        RECT 44.110 160.480 44.430 160.740 ;
        RECT 48.710 160.480 49.030 160.740 ;
        RECT 49.630 160.680 49.950 160.740 ;
        RECT 54.690 160.680 55.010 160.740 ;
        RECT 59.840 160.725 59.980 160.880 ;
        RECT 49.630 160.540 55.010 160.680 ;
        RECT 49.630 160.480 49.950 160.540 ;
        RECT 54.690 160.480 55.010 160.540 ;
        RECT 59.765 160.495 60.055 160.725 ;
        RECT 60.670 160.480 60.990 160.740 ;
        RECT 61.130 160.680 61.450 160.740 ;
        RECT 62.065 160.680 62.355 160.725 ;
        RECT 61.130 160.540 62.355 160.680 ;
        RECT 62.600 160.680 62.740 161.560 ;
        RECT 62.985 161.360 63.275 161.405 ;
        RECT 63.890 161.360 64.210 161.420 ;
        RECT 62.985 161.220 64.210 161.360 ;
        RECT 62.985 161.175 63.275 161.220 ;
        RECT 63.890 161.160 64.210 161.220 ;
        RECT 64.350 161.160 64.670 161.420 ;
        RECT 65.730 161.160 66.050 161.420 ;
        RECT 69.960 161.405 70.100 161.560 ;
        RECT 71.265 161.560 77.920 161.700 ;
        RECT 71.265 161.515 71.555 161.560 ;
        RECT 66.205 161.360 66.495 161.405 ;
        RECT 66.205 161.220 67.340 161.360 ;
        RECT 66.205 161.175 66.495 161.220 ;
        RECT 64.825 161.020 65.115 161.065 ;
        RECT 66.650 161.020 66.970 161.080 ;
        RECT 64.825 160.880 66.970 161.020 ;
        RECT 64.825 160.835 65.115 160.880 ;
        RECT 66.650 160.820 66.970 160.880 ;
        RECT 67.200 160.740 67.340 161.220 ;
        RECT 69.885 161.175 70.175 161.405 ;
        RECT 71.710 161.160 72.030 161.420 ;
        RECT 72.630 161.160 72.950 161.420 ;
        RECT 77.230 161.360 77.550 161.420 ;
        RECT 79.085 161.360 79.375 161.405 ;
        RECT 77.230 161.220 79.375 161.360 ;
        RECT 77.230 161.160 77.550 161.220 ;
        RECT 79.085 161.175 79.375 161.220 ;
        RECT 80.465 161.175 80.755 161.405 ;
        RECT 81.385 161.360 81.675 161.405 ;
        RECT 83.225 161.360 83.515 161.405 ;
        RECT 81.385 161.220 83.515 161.360 ;
        RECT 81.385 161.175 81.675 161.220 ;
        RECT 83.225 161.175 83.515 161.220 ;
        RECT 86.445 161.360 86.735 161.405 ;
        RECT 87.810 161.360 88.130 161.420 ;
        RECT 88.745 161.360 89.035 161.405 ;
        RECT 86.445 161.220 89.035 161.360 ;
        RECT 86.445 161.175 86.735 161.220 ;
        RECT 72.720 161.020 72.860 161.160 ;
        RECT 80.540 161.020 80.680 161.175 ;
        RECT 87.810 161.160 88.130 161.220 ;
        RECT 88.745 161.175 89.035 161.220 ;
        RECT 72.720 160.880 80.680 161.020 ;
        RECT 67.110 160.680 67.430 160.740 ;
        RECT 62.600 160.540 67.430 160.680 ;
        RECT 61.130 160.480 61.450 160.540 ;
        RECT 62.065 160.495 62.355 160.540 ;
        RECT 67.110 160.480 67.430 160.540 ;
        RECT 71.250 160.480 71.570 160.740 ;
        RECT 72.170 160.480 72.490 160.740 ;
        RECT 78.150 160.480 78.470 160.740 ;
        RECT 79.530 160.680 79.850 160.740 ;
        RECT 87.825 160.680 88.115 160.725 ;
        RECT 79.530 160.540 88.115 160.680 ;
        RECT 79.530 160.480 79.850 160.540 ;
        RECT 87.825 160.495 88.115 160.540 ;
        RECT 88.270 160.480 88.590 160.740 ;
        RECT 18.280 159.860 93.120 160.340 ;
        RECT 34.910 159.460 35.230 159.720 ;
        RECT 35.370 159.660 35.690 159.720 ;
        RECT 45.490 159.660 45.810 159.720 ;
        RECT 48.250 159.705 48.570 159.720 ;
        RECT 47.345 159.660 47.635 159.705 ;
        RECT 35.370 159.520 36.060 159.660 ;
        RECT 35.370 159.460 35.690 159.520 ;
        RECT 33.990 159.120 34.310 159.380 ;
        RECT 35.000 159.320 35.140 159.460 ;
        RECT 35.000 159.180 35.600 159.320 ;
        RECT 33.530 158.780 33.850 159.040 ;
        RECT 35.460 159.025 35.600 159.180 ;
        RECT 35.920 159.025 36.060 159.520 ;
        RECT 45.490 159.520 47.635 159.660 ;
        RECT 45.490 159.460 45.810 159.520 ;
        RECT 47.345 159.475 47.635 159.520 ;
        RECT 48.160 159.660 48.570 159.705 ;
        RECT 49.630 159.660 49.950 159.720 ;
        RECT 48.160 159.520 49.950 159.660 ;
        RECT 48.160 159.475 48.570 159.520 ;
        RECT 48.250 159.460 48.570 159.475 ;
        RECT 49.630 159.460 49.950 159.520 ;
        RECT 52.390 159.660 52.710 159.720 ;
        RECT 52.865 159.660 53.155 159.705 ;
        RECT 52.390 159.520 53.155 159.660 ;
        RECT 52.390 159.460 52.710 159.520 ;
        RECT 52.865 159.475 53.155 159.520 ;
        RECT 61.145 159.660 61.435 159.705 ;
        RECT 61.590 159.660 61.910 159.720 ;
        RECT 61.145 159.520 61.910 159.660 ;
        RECT 61.145 159.475 61.435 159.520 ;
        RECT 61.590 159.460 61.910 159.520 ;
        RECT 64.350 159.660 64.670 159.720 ;
        RECT 65.745 159.660 66.035 159.705 ;
        RECT 64.350 159.520 66.035 159.660 ;
        RECT 64.350 159.460 64.670 159.520 ;
        RECT 65.745 159.475 66.035 159.520 ;
        RECT 72.170 159.460 72.490 159.720 ;
        RECT 76.310 159.460 76.630 159.720 ;
        RECT 45.580 159.180 48.020 159.320 ;
        RECT 45.580 159.040 45.720 159.180 ;
        RECT 34.925 158.795 35.215 159.025 ;
        RECT 35.385 158.795 35.675 159.025 ;
        RECT 35.845 158.795 36.135 159.025 ;
        RECT 36.765 158.980 37.055 159.025 ;
        RECT 38.145 158.980 38.435 159.025 ;
        RECT 36.765 158.840 38.435 158.980 ;
        RECT 36.765 158.795 37.055 158.840 ;
        RECT 38.145 158.795 38.435 158.840 ;
        RECT 39.050 158.980 39.370 159.040 ;
        RECT 40.905 158.980 41.195 159.025 ;
        RECT 41.825 158.980 42.115 159.025 ;
        RECT 39.050 158.840 41.195 158.980 ;
        RECT 33.620 158.300 33.760 158.780 ;
        RECT 35.000 158.640 35.140 158.795 ;
        RECT 39.050 158.780 39.370 158.840 ;
        RECT 40.905 158.795 41.195 158.840 ;
        RECT 41.440 158.840 42.115 158.980 ;
        RECT 36.305 158.640 36.595 158.685 ;
        RECT 35.000 158.500 36.595 158.640 ;
        RECT 36.305 158.455 36.595 158.500 ;
        RECT 41.440 158.300 41.580 158.840 ;
        RECT 41.825 158.795 42.115 158.840 ;
        RECT 42.745 158.980 43.035 159.025 ;
        RECT 44.110 158.980 44.430 159.040 ;
        RECT 42.745 158.840 44.430 158.980 ;
        RECT 42.745 158.795 43.035 158.840 ;
        RECT 44.110 158.780 44.430 158.840 ;
        RECT 45.490 158.780 45.810 159.040 ;
        RECT 46.425 158.795 46.715 159.025 ;
        RECT 46.885 158.980 47.175 159.025 ;
        RECT 47.330 158.980 47.650 159.040 ;
        RECT 46.885 158.840 47.650 158.980 ;
        RECT 47.880 158.980 48.020 159.180 ;
        RECT 49.185 159.135 49.475 159.365 ;
        RECT 54.705 159.320 54.995 159.365 ;
        RECT 57.450 159.320 57.770 159.380 ;
        RECT 72.260 159.320 72.400 159.460 ;
        RECT 54.705 159.180 57.770 159.320 ;
        RECT 54.705 159.135 54.995 159.180 ;
        RECT 48.710 158.980 49.030 159.040 ;
        RECT 49.260 158.980 49.400 159.135 ;
        RECT 57.450 159.120 57.770 159.180 ;
        RECT 71.800 159.180 72.400 159.320 ;
        RECT 73.105 159.320 73.395 159.365 ;
        RECT 76.400 159.320 76.540 159.460 ;
        RECT 73.105 159.180 76.540 159.320 ;
        RECT 80.470 159.320 80.760 159.365 ;
        RECT 81.870 159.320 82.160 159.365 ;
        RECT 83.710 159.320 84.000 159.365 ;
        RECT 80.470 159.180 84.000 159.320 ;
        RECT 49.645 158.980 49.935 159.025 ;
        RECT 47.880 158.840 49.935 158.980 ;
        RECT 46.885 158.795 47.175 158.840 ;
        RECT 45.950 158.440 46.270 158.700 ;
        RECT 46.500 158.640 46.640 158.795 ;
        RECT 47.330 158.780 47.650 158.840 ;
        RECT 48.710 158.780 49.030 158.840 ;
        RECT 49.645 158.795 49.935 158.840 ;
        RECT 52.850 158.980 53.170 159.040 ;
        RECT 53.325 158.980 53.615 159.025 ;
        RECT 52.850 158.840 53.615 158.980 ;
        RECT 52.850 158.780 53.170 158.840 ;
        RECT 53.325 158.795 53.615 158.840 ;
        RECT 54.245 158.980 54.535 159.025 ;
        RECT 60.670 158.980 60.990 159.040 ;
        RECT 71.800 159.025 71.940 159.180 ;
        RECT 73.105 159.135 73.395 159.180 ;
        RECT 80.470 159.135 80.760 159.180 ;
        RECT 81.870 159.135 82.160 159.180 ;
        RECT 83.710 159.135 84.000 159.180 ;
        RECT 54.245 158.840 60.990 158.980 ;
        RECT 54.245 158.795 54.535 158.840 ;
        RECT 60.670 158.780 60.990 158.840 ;
        RECT 71.725 158.795 72.015 159.025 ;
        RECT 72.185 158.795 72.475 159.025 ;
        RECT 49.170 158.640 49.490 158.700 ;
        RECT 46.500 158.500 49.490 158.640 ;
        RECT 49.170 158.440 49.490 158.500 ;
        RECT 45.505 158.300 45.795 158.345 ;
        RECT 46.040 158.300 46.180 158.440 ;
        RECT 52.940 158.300 53.080 158.780 ;
        RECT 67.110 158.640 67.430 158.700 ;
        RECT 68.505 158.640 68.795 158.685 ;
        RECT 67.110 158.500 68.795 158.640 ;
        RECT 67.110 158.440 67.430 158.500 ;
        RECT 68.505 158.455 68.795 158.500 ;
        RECT 71.250 158.640 71.570 158.700 ;
        RECT 72.260 158.640 72.400 158.795 ;
        RECT 75.850 158.780 76.170 159.040 ;
        RECT 78.150 158.980 78.470 159.040 ;
        RECT 80.925 158.980 81.215 159.025 ;
        RECT 78.150 158.840 81.215 158.980 ;
        RECT 78.150 158.780 78.470 158.840 ;
        RECT 80.925 158.795 81.215 158.840 ;
        RECT 71.250 158.500 72.400 158.640 ;
        RECT 79.545 158.640 79.835 158.685 ;
        RECT 80.450 158.640 80.770 158.700 ;
        RECT 79.545 158.500 80.770 158.640 ;
        RECT 71.250 158.440 71.570 158.500 ;
        RECT 79.545 158.455 79.835 158.500 ;
        RECT 80.450 158.440 80.770 158.500 ;
        RECT 33.620 158.160 45.260 158.300 ;
        RECT 33.990 157.760 34.310 158.020 ;
        RECT 41.810 157.960 42.130 158.020 ;
        RECT 42.745 157.960 43.035 158.005 ;
        RECT 41.810 157.820 43.035 157.960 ;
        RECT 45.120 157.960 45.260 158.160 ;
        RECT 45.505 158.160 46.180 158.300 ;
        RECT 46.500 158.160 53.080 158.300 ;
        RECT 80.010 158.300 80.300 158.345 ;
        RECT 82.330 158.300 82.620 158.345 ;
        RECT 83.710 158.300 84.000 158.345 ;
        RECT 80.010 158.160 84.000 158.300 ;
        RECT 45.505 158.115 45.795 158.160 ;
        RECT 46.500 157.960 46.640 158.160 ;
        RECT 80.010 158.115 80.300 158.160 ;
        RECT 82.330 158.115 82.620 158.160 ;
        RECT 83.710 158.115 84.000 158.160 ;
        RECT 45.120 157.820 46.640 157.960 ;
        RECT 48.265 157.960 48.555 158.005 ;
        RECT 49.170 157.960 49.490 158.020 ;
        RECT 48.265 157.820 49.490 157.960 ;
        RECT 41.810 157.760 42.130 157.820 ;
        RECT 42.745 157.775 43.035 157.820 ;
        RECT 48.265 157.775 48.555 157.820 ;
        RECT 49.170 157.760 49.490 157.820 ;
        RECT 54.230 157.760 54.550 158.020 ;
        RECT 73.105 157.960 73.395 158.005 ;
        RECT 73.550 157.960 73.870 158.020 ;
        RECT 73.105 157.820 73.870 157.960 ;
        RECT 73.105 157.775 73.395 157.820 ;
        RECT 73.550 157.760 73.870 157.820 ;
        RECT 87.365 157.960 87.655 158.005 ;
        RECT 87.810 157.960 88.130 158.020 ;
        RECT 87.365 157.820 88.130 157.960 ;
        RECT 87.365 157.775 87.655 157.820 ;
        RECT 87.810 157.760 88.130 157.820 ;
        RECT 18.280 157.140 92.340 157.620 ;
        RECT 39.050 156.740 39.370 157.000 ;
        RECT 46.870 156.940 47.190 157.000 ;
        RECT 47.345 156.940 47.635 156.985 ;
        RECT 46.870 156.800 47.635 156.940 ;
        RECT 46.870 156.740 47.190 156.800 ;
        RECT 47.345 156.755 47.635 156.800 ;
        RECT 49.170 156.940 49.490 157.000 ;
        RECT 49.645 156.940 49.935 156.985 ;
        RECT 49.170 156.800 49.935 156.940 ;
        RECT 49.170 156.740 49.490 156.800 ;
        RECT 49.645 156.755 49.935 156.800 ;
        RECT 67.110 156.740 67.430 157.000 ;
        RECT 79.070 156.940 79.390 157.000 ;
        RECT 80.005 156.940 80.295 156.985 ;
        RECT 88.270 156.940 88.590 157.000 ;
        RECT 79.070 156.800 88.590 156.940 ;
        RECT 79.070 156.740 79.390 156.800 ;
        RECT 80.005 156.755 80.295 156.800 ;
        RECT 88.270 156.740 88.590 156.800 ;
        RECT 32.650 156.600 32.940 156.645 ;
        RECT 34.750 156.600 35.040 156.645 ;
        RECT 36.320 156.600 36.610 156.645 ;
        RECT 32.650 156.460 36.610 156.600 ;
        RECT 32.650 156.415 32.940 156.460 ;
        RECT 34.750 156.415 35.040 156.460 ;
        RECT 36.320 156.415 36.610 156.460 ;
        RECT 40.930 156.600 41.220 156.645 ;
        RECT 43.030 156.600 43.320 156.645 ;
        RECT 44.600 156.600 44.890 156.645 ;
        RECT 40.930 156.460 44.890 156.600 ;
        RECT 40.930 156.415 41.220 156.460 ;
        RECT 43.030 156.415 43.320 156.460 ;
        RECT 44.600 156.415 44.890 156.460 ;
        RECT 52.390 156.600 52.680 156.645 ;
        RECT 53.960 156.600 54.250 156.645 ;
        RECT 56.060 156.600 56.350 156.645 ;
        RECT 52.390 156.460 56.350 156.600 ;
        RECT 52.390 156.415 52.680 156.460 ;
        RECT 53.960 156.415 54.250 156.460 ;
        RECT 56.060 156.415 56.350 156.460 ;
        RECT 60.710 156.600 61.000 156.645 ;
        RECT 62.810 156.600 63.100 156.645 ;
        RECT 64.380 156.600 64.670 156.645 ;
        RECT 60.710 156.460 64.670 156.600 ;
        RECT 60.710 156.415 61.000 156.460 ;
        RECT 62.810 156.415 63.100 156.460 ;
        RECT 64.380 156.415 64.670 156.460 ;
        RECT 72.650 156.600 72.940 156.645 ;
        RECT 74.970 156.600 75.260 156.645 ;
        RECT 76.350 156.600 76.640 156.645 ;
        RECT 72.650 156.460 76.640 156.600 ;
        RECT 72.650 156.415 72.940 156.460 ;
        RECT 74.970 156.415 75.260 156.460 ;
        RECT 76.350 156.415 76.640 156.460 ;
        RECT 32.150 156.060 32.470 156.320 ;
        RECT 33.045 156.260 33.335 156.305 ;
        RECT 34.235 156.260 34.525 156.305 ;
        RECT 36.755 156.260 37.045 156.305 ;
        RECT 33.045 156.120 37.045 156.260 ;
        RECT 33.045 156.075 33.335 156.120 ;
        RECT 34.235 156.075 34.525 156.120 ;
        RECT 36.755 156.075 37.045 156.120 ;
        RECT 41.325 156.260 41.615 156.305 ;
        RECT 42.515 156.260 42.805 156.305 ;
        RECT 45.035 156.260 45.325 156.305 ;
        RECT 41.325 156.120 45.325 156.260 ;
        RECT 41.325 156.075 41.615 156.120 ;
        RECT 42.515 156.075 42.805 156.120 ;
        RECT 45.035 156.075 45.325 156.120 ;
        RECT 51.955 156.260 52.245 156.305 ;
        RECT 54.475 156.260 54.765 156.305 ;
        RECT 55.665 156.260 55.955 156.305 ;
        RECT 51.955 156.120 55.955 156.260 ;
        RECT 51.955 156.075 52.245 156.120 ;
        RECT 54.475 156.075 54.765 156.120 ;
        RECT 55.665 156.075 55.955 156.120 ;
        RECT 61.105 156.260 61.395 156.305 ;
        RECT 62.295 156.260 62.585 156.305 ;
        RECT 64.815 156.260 65.105 156.305 ;
        RECT 72.185 156.260 72.475 156.305 ;
        RECT 80.450 156.260 80.770 156.320 ;
        RECT 61.105 156.120 65.105 156.260 ;
        RECT 61.105 156.075 61.395 156.120 ;
        RECT 62.295 156.075 62.585 156.120 ;
        RECT 64.815 156.075 65.105 156.120 ;
        RECT 70.650 156.120 80.770 156.260 ;
        RECT 32.240 155.920 32.380 156.060 ;
        RECT 41.810 155.965 42.130 155.980 ;
        RECT 40.445 155.920 40.735 155.965 ;
        RECT 41.780 155.920 42.130 155.965 ;
        RECT 32.240 155.780 40.735 155.920 ;
        RECT 41.615 155.780 42.130 155.920 ;
        RECT 40.445 155.735 40.735 155.780 ;
        RECT 41.780 155.735 42.130 155.780 ;
        RECT 41.810 155.720 42.130 155.735 ;
        RECT 55.150 155.965 55.470 155.980 ;
        RECT 55.150 155.735 55.500 155.965 ;
        RECT 56.545 155.920 56.835 155.965 ;
        RECT 60.225 155.920 60.515 155.965 ;
        RECT 62.970 155.920 63.290 155.980 ;
        RECT 70.650 155.920 70.790 156.120 ;
        RECT 72.185 156.075 72.475 156.120 ;
        RECT 80.450 156.060 80.770 156.120 ;
        RECT 56.545 155.780 70.790 155.920 ;
        RECT 56.545 155.735 56.835 155.780 ;
        RECT 60.225 155.735 60.515 155.780 ;
        RECT 55.150 155.720 55.470 155.735 ;
        RECT 62.970 155.720 63.290 155.780 ;
        RECT 73.550 155.720 73.870 155.980 ;
        RECT 33.500 155.580 33.790 155.625 ;
        RECT 33.990 155.580 34.310 155.640 ;
        RECT 33.500 155.440 34.310 155.580 ;
        RECT 33.500 155.395 33.790 155.440 ;
        RECT 33.990 155.380 34.310 155.440 ;
        RECT 61.560 155.580 61.850 155.625 ;
        RECT 62.050 155.580 62.370 155.640 ;
        RECT 61.560 155.440 62.370 155.580 ;
        RECT 61.560 155.395 61.850 155.440 ;
        RECT 62.050 155.380 62.370 155.440 ;
        RECT 73.110 155.580 73.400 155.625 ;
        RECT 74.510 155.580 74.800 155.625 ;
        RECT 76.350 155.580 76.640 155.625 ;
        RECT 73.110 155.440 76.640 155.580 ;
        RECT 73.110 155.395 73.400 155.440 ;
        RECT 74.510 155.395 74.800 155.440 ;
        RECT 76.350 155.395 76.640 155.440 ;
        RECT 112.400 155.300 113.000 155.330 ;
        RECT 117.370 155.300 118.030 155.900 ;
        RECT 18.280 154.420 93.120 154.900 ;
        RECT 112.400 154.700 114.600 155.300 ;
        RECT 112.400 154.670 113.000 154.700 ;
        RECT 18.280 151.700 92.340 152.180 ;
        RECT 71.725 151.500 72.015 151.545 ;
        RECT 77.230 151.500 77.550 151.560 ;
        RECT 79.530 151.500 79.850 151.560 ;
        RECT 71.725 151.360 79.850 151.500 ;
        RECT 71.725 151.315 72.015 151.360 ;
        RECT 77.230 151.300 77.550 151.360 ;
        RECT 79.530 151.300 79.850 151.360 ;
        RECT 64.370 151.160 64.660 151.205 ;
        RECT 66.690 151.160 66.980 151.205 ;
        RECT 68.070 151.160 68.360 151.205 ;
        RECT 64.370 151.020 68.360 151.160 ;
        RECT 64.370 150.975 64.660 151.020 ;
        RECT 66.690 150.975 66.980 151.020 ;
        RECT 68.070 150.975 68.360 151.020 ;
        RECT 62.970 150.820 63.290 150.880 ;
        RECT 63.905 150.820 64.195 150.865 ;
        RECT 62.970 150.680 64.195 150.820 ;
        RECT 62.970 150.620 63.290 150.680 ;
        RECT 63.905 150.635 64.195 150.680 ;
        RECT 65.270 150.620 65.590 150.880 ;
        RECT 64.830 150.140 65.120 150.185 ;
        RECT 66.230 150.140 66.520 150.185 ;
        RECT 68.070 150.140 68.360 150.185 ;
        RECT 64.830 150.000 68.360 150.140 ;
        RECT 64.830 149.955 65.120 150.000 ;
        RECT 66.230 149.955 66.520 150.000 ;
        RECT 68.070 149.955 68.360 150.000 ;
        RECT 18.280 148.980 93.120 149.460 ;
        RECT 107.000 149.000 107.600 149.030 ;
        RECT 107.000 148.400 113.200 149.000 ;
        RECT 107.000 148.370 107.600 148.400 ;
        RECT 112.600 146.930 113.200 148.400 ;
        RECT 114.000 146.930 114.600 154.700 ;
        RECT 115.870 152.500 116.530 153.100 ;
        RECT 115.900 146.930 116.500 152.500 ;
        RECT 117.400 146.930 118.000 155.300 ;
        RECT 118.870 155.200 119.530 155.800 ;
        RECT 118.900 146.930 119.500 155.200 ;
        RECT 120.370 155.100 121.030 155.700 ;
        RECT 120.400 146.930 121.000 155.100 ;
        RECT 121.770 154.100 122.430 154.700 ;
        RECT 121.800 149.000 122.400 154.100 ;
        RECT 121.800 148.400 122.900 149.000 ;
        RECT 122.300 146.930 122.900 148.400 ;
        RECT 18.280 146.260 92.340 146.740 ;
        RECT 106.700 146.700 107.300 146.730 ;
        RECT 110.780 146.700 111.780 146.930 ;
        RECT 106.700 146.100 111.780 146.700 ;
        RECT 106.700 146.070 107.300 146.100 ;
        RECT 110.780 145.930 111.780 146.100 ;
        RECT 112.380 145.930 113.380 146.930 ;
        RECT 113.880 145.930 114.880 146.930 ;
        RECT 115.480 146.100 116.500 146.930 ;
        RECT 115.480 145.930 116.480 146.100 ;
        RECT 117.080 145.930 118.080 146.930 ;
        RECT 118.680 145.930 119.680 146.930 ;
        RECT 120.280 145.930 121.280 146.930 ;
        RECT 121.980 146.540 122.980 146.930 ;
        RECT 121.970 145.930 122.980 146.540 ;
        RECT 111.350 144.640 111.650 145.930 ;
        RECT 112.820 145.300 113.120 145.930 ;
        RECT 114.530 145.680 114.830 145.930 ;
        RECT 114.530 145.380 115.320 145.680 ;
        RECT 112.820 145.000 114.320 145.300 ;
        RECT 113.040 144.640 113.290 144.820 ;
        RECT 111.350 144.340 113.300 144.640 ;
        RECT 114.020 144.370 114.320 145.000 ;
        RECT 18.280 143.540 93.120 144.020 ;
        RECT 113.040 142.715 113.290 144.340 ;
        RECT 114.040 142.715 114.290 144.370 ;
        RECT 115.020 144.340 115.320 145.380 ;
        RECT 116.010 144.460 116.310 145.930 ;
        RECT 117.310 145.490 117.610 145.930 ;
        RECT 118.770 145.770 119.070 145.930 ;
        RECT 117.010 145.190 117.610 145.490 ;
        RECT 118.300 145.470 119.070 145.770 ;
        RECT 120.470 145.740 120.770 145.930 ;
        RECT 118.300 145.350 118.600 145.470 ;
        RECT 115.040 142.715 115.290 144.340 ;
        RECT 116.040 142.715 116.290 144.460 ;
        RECT 117.010 144.450 117.310 145.190 ;
        RECT 118.040 145.050 118.600 145.350 ;
        RECT 119.620 145.440 120.770 145.740 ;
        RECT 119.620 145.310 119.920 145.440 ;
        RECT 118.040 144.460 118.340 145.050 ;
        RECT 119.030 145.010 119.920 145.310 ;
        RECT 119.030 144.490 119.330 145.010 ;
        RECT 120.040 144.780 120.290 144.820 ;
        RECT 121.970 144.780 122.270 145.930 ;
        RECT 117.040 142.715 117.290 144.450 ;
        RECT 118.040 142.715 118.290 144.460 ;
        RECT 119.040 142.715 119.290 144.490 ;
        RECT 119.980 144.480 122.270 144.780 ;
        RECT 120.040 142.715 120.290 144.480 ;
        RECT 18.280 140.820 92.340 141.300 ;
        RECT 113.040 140.540 113.290 141.665 ;
        RECT 114.040 140.550 114.290 141.665 ;
        RECT 113.900 140.540 114.740 140.550 ;
        RECT 18.280 138.100 93.120 138.580 ;
        RECT 113.030 138.250 113.330 140.540 ;
        RECT 113.900 139.530 114.820 140.540 ;
        RECT 115.040 140.500 115.290 141.665 ;
        RECT 116.040 140.690 116.290 141.665 ;
        RECT 114.040 138.250 114.290 138.320 ;
        RECT 112.940 137.470 114.360 138.250 ;
        RECT 113.040 136.715 113.290 137.470 ;
        RECT 114.040 136.215 114.290 137.470 ;
        RECT 18.280 135.380 92.340 135.860 ;
        RECT 111.380 134.220 112.380 134.530 ;
        RECT 113.040 134.220 113.290 135.665 ;
        RECT 114.040 134.410 114.290 135.665 ;
        RECT 114.510 134.410 114.820 139.530 ;
        RECT 115.000 138.280 115.350 140.500 ;
        RECT 116.020 139.670 116.790 140.690 ;
        RECT 117.040 140.580 117.290 141.665 ;
        RECT 118.040 140.760 118.290 141.665 ;
        RECT 116.040 139.560 116.290 139.670 ;
        RECT 116.040 138.280 116.290 138.320 ;
        RECT 114.980 137.500 116.400 138.280 ;
        RECT 115.040 136.215 115.290 137.500 ;
        RECT 116.040 136.215 116.290 137.500 ;
        RECT 111.380 133.770 113.290 134.220 ;
        RECT 111.380 133.530 112.380 133.770 ;
        RECT 113.040 133.560 113.290 133.770 ;
        RECT 114.010 134.380 114.820 134.410 ;
        RECT 115.040 134.380 115.290 135.665 ;
        RECT 116.040 134.390 116.290 135.665 ;
        RECT 116.540 134.400 116.790 139.670 ;
        RECT 117.000 138.360 117.350 140.580 ;
        RECT 117.970 139.740 118.810 140.760 ;
        RECT 119.040 140.600 119.290 141.665 ;
        RECT 118.040 139.560 118.290 139.740 ;
        RECT 118.490 139.710 118.800 139.740 ;
        RECT 116.950 138.320 118.240 138.360 ;
        RECT 116.950 137.580 118.290 138.320 ;
        RECT 117.040 136.215 117.290 137.580 ;
        RECT 118.040 136.215 118.290 137.580 ;
        RECT 116.540 134.390 116.850 134.400 ;
        RECT 117.040 134.390 117.290 135.665 ;
        RECT 118.040 134.440 118.290 135.665 ;
        RECT 118.000 134.430 118.290 134.440 ;
        RECT 118.530 134.440 118.800 139.710 ;
        RECT 119.000 138.370 119.350 140.600 ;
        RECT 120.040 140.380 120.290 141.665 ;
        RECT 119.920 139.870 120.340 140.380 ;
        RECT 119.920 139.330 121.510 139.870 ;
        RECT 119.920 138.840 125.700 139.330 ;
        RECT 119.990 138.830 125.700 138.840 ;
        RECT 120.760 138.510 125.700 138.830 ;
        RECT 118.950 137.590 120.370 138.370 ;
        RECT 119.040 136.215 119.290 137.590 ;
        RECT 120.040 136.215 120.290 137.590 ;
        RECT 119.040 134.440 119.290 135.665 ;
        RECT 118.530 134.430 119.330 134.440 ;
        RECT 114.010 133.680 115.350 134.380 ;
        RECT 116.010 133.690 117.340 134.390 ;
        RECT 118.000 133.740 119.330 134.430 ;
        RECT 120.040 134.420 120.290 135.665 ;
        RECT 120.810 134.420 121.240 138.510 ;
        RECT 121.480 138.330 125.700 138.510 ;
        RECT 114.010 133.610 114.760 133.680 ;
        RECT 114.040 133.560 114.290 133.610 ;
        RECT 115.040 133.560 115.290 133.680 ;
        RECT 116.040 133.560 116.290 133.690 ;
        RECT 117.040 133.560 117.290 133.690 ;
        RECT 118.040 133.560 118.290 133.740 ;
        RECT 119.040 133.560 119.290 133.740 ;
        RECT 119.960 133.720 121.290 134.420 ;
        RECT 120.040 133.560 120.290 133.720 ;
        RECT 18.280 132.660 93.120 133.140 ;
        RECT 124.715 30.400 125.690 138.330 ;
        RECT 124.715 27.915 125.700 30.400 ;
        RECT 125.100 26.400 125.700 27.915 ;
        RECT 130.300 26.400 130.900 26.430 ;
        RECT 125.100 25.800 130.900 26.400 ;
        RECT 130.300 25.770 130.900 25.800 ;
      LAYER via ;
        RECT 40.460 206.720 40.720 206.980 ;
        RECT 76.340 206.720 76.600 206.980 ;
        RECT 26.765 206.210 27.025 206.470 ;
        RECT 27.085 206.210 27.345 206.470 ;
        RECT 27.405 206.210 27.665 206.470 ;
        RECT 27.725 206.210 27.985 206.470 ;
        RECT 28.045 206.210 28.305 206.470 ;
        RECT 45.275 206.210 45.535 206.470 ;
        RECT 45.595 206.210 45.855 206.470 ;
        RECT 45.915 206.210 46.175 206.470 ;
        RECT 46.235 206.210 46.495 206.470 ;
        RECT 46.555 206.210 46.815 206.470 ;
        RECT 63.785 206.210 64.045 206.470 ;
        RECT 64.105 206.210 64.365 206.470 ;
        RECT 64.425 206.210 64.685 206.470 ;
        RECT 64.745 206.210 65.005 206.470 ;
        RECT 65.065 206.210 65.325 206.470 ;
        RECT 82.295 206.210 82.555 206.470 ;
        RECT 82.615 206.210 82.875 206.470 ;
        RECT 82.935 206.210 83.195 206.470 ;
        RECT 83.255 206.210 83.515 206.470 ;
        RECT 83.575 206.210 83.835 206.470 ;
        RECT 45.980 205.700 46.240 205.960 ;
        RECT 46.900 205.700 47.160 205.960 ;
        RECT 47.820 205.700 48.080 205.960 ;
        RECT 72.660 205.700 72.920 205.960 ;
        RECT 65.760 205.360 66.020 205.620 ;
        RECT 71.280 205.360 71.540 205.620 ;
        RECT 26.200 204.680 26.460 204.940 ;
        RECT 32.640 204.680 32.900 204.940 ;
        RECT 39.080 204.680 39.340 204.940 ;
        RECT 45.520 204.680 45.780 204.940 ;
        RECT 46.900 204.680 47.160 204.940 ;
        RECT 47.360 204.680 47.620 204.940 ;
        RECT 51.960 204.680 52.220 204.940 ;
        RECT 57.480 204.680 57.740 204.940 ;
        RECT 40.460 204.340 40.720 204.600 ;
        RECT 58.400 204.680 58.660 204.940 ;
        RECT 26.200 204.000 26.460 204.260 ;
        RECT 28.500 204.000 28.760 204.260 ;
        RECT 44.140 204.000 44.400 204.260 ;
        RECT 44.600 204.000 44.860 204.260 ;
        RECT 57.940 204.340 58.200 204.600 ;
        RECT 66.220 204.680 66.480 204.940 ;
        RECT 79.560 205.360 79.820 205.620 ;
        RECT 77.720 204.680 77.980 204.940 ;
        RECT 81.400 204.680 81.660 204.940 ;
        RECT 84.160 204.680 84.420 204.940 ;
        RECT 90.600 204.680 90.860 204.940 ;
        RECT 53.340 204.000 53.600 204.260 ;
        RECT 60.240 204.000 60.500 204.260 ;
        RECT 60.700 204.000 60.960 204.260 ;
        RECT 63.000 204.000 63.260 204.260 ;
        RECT 67.600 204.000 67.860 204.260 ;
        RECT 72.200 204.000 72.460 204.260 ;
        RECT 75.420 204.000 75.680 204.260 ;
        RECT 76.800 204.000 77.060 204.260 ;
        RECT 79.100 204.000 79.360 204.260 ;
        RECT 81.860 204.000 82.120 204.260 ;
        RECT 84.620 204.000 84.880 204.260 ;
        RECT 86.460 204.000 86.720 204.260 ;
        RECT 36.020 203.490 36.280 203.750 ;
        RECT 36.340 203.490 36.600 203.750 ;
        RECT 36.660 203.490 36.920 203.750 ;
        RECT 36.980 203.490 37.240 203.750 ;
        RECT 37.300 203.490 37.560 203.750 ;
        RECT 54.530 203.490 54.790 203.750 ;
        RECT 54.850 203.490 55.110 203.750 ;
        RECT 55.170 203.490 55.430 203.750 ;
        RECT 55.490 203.490 55.750 203.750 ;
        RECT 55.810 203.490 56.070 203.750 ;
        RECT 73.040 203.490 73.300 203.750 ;
        RECT 73.360 203.490 73.620 203.750 ;
        RECT 73.680 203.490 73.940 203.750 ;
        RECT 74.000 203.490 74.260 203.750 ;
        RECT 74.320 203.490 74.580 203.750 ;
        RECT 91.550 203.490 91.810 203.750 ;
        RECT 91.870 203.490 92.130 203.750 ;
        RECT 92.190 203.490 92.450 203.750 ;
        RECT 92.510 203.490 92.770 203.750 ;
        RECT 92.830 203.490 93.090 203.750 ;
        RECT 26.200 202.980 26.460 203.240 ;
        RECT 28.960 202.640 29.220 202.900 ;
        RECT 44.600 202.980 44.860 203.240 ;
        RECT 52.420 202.980 52.680 203.240 ;
        RECT 57.480 202.980 57.740 203.240 ;
        RECT 62.540 202.980 62.800 203.240 ;
        RECT 66.220 202.980 66.480 203.240 ;
        RECT 75.420 202.980 75.680 203.240 ;
        RECT 81.400 202.980 81.660 203.240 ;
        RECT 47.820 202.640 48.080 202.900 ;
        RECT 43.220 202.300 43.480 202.560 ;
        RECT 45.520 202.300 45.780 202.560 ;
        RECT 32.180 201.960 32.440 202.220 ;
        RECT 46.900 201.960 47.160 202.220 ;
        RECT 53.340 202.300 53.600 202.560 ;
        RECT 57.020 202.300 57.280 202.560 ;
        RECT 66.680 202.300 66.940 202.560 ;
        RECT 67.140 202.300 67.400 202.560 ;
        RECT 75.880 202.300 76.140 202.560 ;
        RECT 79.560 202.300 79.820 202.560 ;
        RECT 80.020 202.300 80.280 202.560 ;
        RECT 80.480 202.300 80.740 202.560 ;
        RECT 80.940 202.300 81.200 202.560 ;
        RECT 90.600 202.300 90.860 202.560 ;
        RECT 34.940 201.620 35.200 201.880 ;
        RECT 31.260 201.280 31.520 201.540 ;
        RECT 44.600 201.280 44.860 201.540 ;
        RECT 45.980 201.280 46.240 201.540 ;
        RECT 46.900 201.280 47.160 201.540 ;
        RECT 48.280 201.280 48.540 201.540 ;
        RECT 50.120 201.280 50.380 201.540 ;
        RECT 77.720 201.280 77.980 201.540 ;
        RECT 84.160 201.960 84.420 202.220 ;
        RECT 85.540 201.280 85.800 201.540 ;
        RECT 26.765 200.770 27.025 201.030 ;
        RECT 27.085 200.770 27.345 201.030 ;
        RECT 27.405 200.770 27.665 201.030 ;
        RECT 27.725 200.770 27.985 201.030 ;
        RECT 28.045 200.770 28.305 201.030 ;
        RECT 45.275 200.770 45.535 201.030 ;
        RECT 45.595 200.770 45.855 201.030 ;
        RECT 45.915 200.770 46.175 201.030 ;
        RECT 46.235 200.770 46.495 201.030 ;
        RECT 46.555 200.770 46.815 201.030 ;
        RECT 63.785 200.770 64.045 201.030 ;
        RECT 64.105 200.770 64.365 201.030 ;
        RECT 64.425 200.770 64.685 201.030 ;
        RECT 64.745 200.770 65.005 201.030 ;
        RECT 65.065 200.770 65.325 201.030 ;
        RECT 82.295 200.770 82.555 201.030 ;
        RECT 82.615 200.770 82.875 201.030 ;
        RECT 82.935 200.770 83.195 201.030 ;
        RECT 83.255 200.770 83.515 201.030 ;
        RECT 83.575 200.770 83.835 201.030 ;
        RECT 28.500 200.260 28.760 200.520 ;
        RECT 28.960 200.260 29.220 200.520 ;
        RECT 34.940 200.260 35.200 200.520 ;
        RECT 46.900 200.260 47.160 200.520 ;
        RECT 43.680 199.920 43.940 200.180 ;
        RECT 47.360 199.920 47.620 200.180 ;
        RECT 48.280 199.920 48.540 200.180 ;
        RECT 57.020 200.260 57.280 200.520 ;
        RECT 58.400 200.260 58.660 200.520 ;
        RECT 66.680 200.260 66.940 200.520 ;
        RECT 75.880 200.260 76.140 200.520 ;
        RECT 80.940 200.260 81.200 200.520 ;
        RECT 84.160 200.260 84.420 200.520 ;
        RECT 32.180 199.240 32.440 199.500 ;
        RECT 43.220 199.240 43.480 199.500 ;
        RECT 44.140 199.240 44.400 199.500 ;
        RECT 50.120 199.580 50.380 199.840 ;
        RECT 60.240 199.580 60.500 199.840 ;
        RECT 63.000 199.580 63.260 199.840 ;
        RECT 76.800 199.920 77.060 200.180 ;
        RECT 72.200 199.580 72.460 199.840 ;
        RECT 79.560 199.580 79.820 199.840 ;
        RECT 58.860 199.240 59.120 199.500 ;
        RECT 65.300 199.240 65.560 199.500 ;
        RECT 67.600 199.240 67.860 199.500 ;
        RECT 74.960 199.240 75.220 199.500 ;
        RECT 76.340 199.240 76.600 199.500 ;
        RECT 90.600 199.580 90.860 199.840 ;
        RECT 81.860 199.240 82.120 199.500 ;
        RECT 84.620 199.240 84.880 199.500 ;
        RECT 44.600 198.560 44.860 198.820 ;
        RECT 53.340 198.560 53.600 198.820 ;
        RECT 68.060 198.560 68.320 198.820 ;
        RECT 81.860 198.560 82.120 198.820 ;
        RECT 82.320 198.560 82.580 198.820 ;
        RECT 36.020 198.050 36.280 198.310 ;
        RECT 36.340 198.050 36.600 198.310 ;
        RECT 36.660 198.050 36.920 198.310 ;
        RECT 36.980 198.050 37.240 198.310 ;
        RECT 37.300 198.050 37.560 198.310 ;
        RECT 54.530 198.050 54.790 198.310 ;
        RECT 54.850 198.050 55.110 198.310 ;
        RECT 55.170 198.050 55.430 198.310 ;
        RECT 55.490 198.050 55.750 198.310 ;
        RECT 55.810 198.050 56.070 198.310 ;
        RECT 73.040 198.050 73.300 198.310 ;
        RECT 73.360 198.050 73.620 198.310 ;
        RECT 73.680 198.050 73.940 198.310 ;
        RECT 74.000 198.050 74.260 198.310 ;
        RECT 74.320 198.050 74.580 198.310 ;
        RECT 91.550 198.050 91.810 198.310 ;
        RECT 91.870 198.050 92.130 198.310 ;
        RECT 92.190 198.050 92.450 198.310 ;
        RECT 92.510 198.050 92.770 198.310 ;
        RECT 92.830 198.050 93.090 198.310 ;
        RECT 47.820 196.860 48.080 197.120 ;
        RECT 58.860 196.860 59.120 197.120 ;
        RECT 59.780 196.860 60.040 197.120 ;
        RECT 79.100 197.540 79.360 197.800 ;
        RECT 84.620 197.540 84.880 197.800 ;
        RECT 65.300 196.860 65.560 197.120 ;
        RECT 74.960 196.860 75.220 197.120 ;
        RECT 78.640 196.860 78.900 197.120 ;
        RECT 84.160 197.200 84.420 197.460 ;
        RECT 57.940 196.520 58.200 196.780 ;
        RECT 66.220 196.520 66.480 196.780 ;
        RECT 71.740 196.520 72.000 196.780 ;
        RECT 60.700 196.180 60.960 196.440 ;
        RECT 77.260 196.520 77.520 196.780 ;
        RECT 82.320 196.520 82.580 196.780 ;
        RECT 85.540 196.860 85.800 197.120 ;
        RECT 86.460 196.860 86.720 197.120 ;
        RECT 87.840 196.860 88.100 197.120 ;
        RECT 84.160 196.520 84.420 196.780 ;
        RECT 47.820 195.840 48.080 196.100 ;
        RECT 53.800 195.840 54.060 196.100 ;
        RECT 58.400 195.840 58.660 196.100 ;
        RECT 58.860 195.840 59.120 196.100 ;
        RECT 63.000 195.840 63.260 196.100 ;
        RECT 65.760 195.840 66.020 196.100 ;
        RECT 74.960 195.840 75.220 196.100 ;
        RECT 80.480 195.840 80.740 196.100 ;
        RECT 85.080 195.840 85.340 196.100 ;
        RECT 86.460 195.840 86.720 196.100 ;
        RECT 26.765 195.330 27.025 195.590 ;
        RECT 27.085 195.330 27.345 195.590 ;
        RECT 27.405 195.330 27.665 195.590 ;
        RECT 27.725 195.330 27.985 195.590 ;
        RECT 28.045 195.330 28.305 195.590 ;
        RECT 45.275 195.330 45.535 195.590 ;
        RECT 45.595 195.330 45.855 195.590 ;
        RECT 45.915 195.330 46.175 195.590 ;
        RECT 46.235 195.330 46.495 195.590 ;
        RECT 46.555 195.330 46.815 195.590 ;
        RECT 63.785 195.330 64.045 195.590 ;
        RECT 64.105 195.330 64.365 195.590 ;
        RECT 64.425 195.330 64.685 195.590 ;
        RECT 64.745 195.330 65.005 195.590 ;
        RECT 65.065 195.330 65.325 195.590 ;
        RECT 82.295 195.330 82.555 195.590 ;
        RECT 82.615 195.330 82.875 195.590 ;
        RECT 82.935 195.330 83.195 195.590 ;
        RECT 83.255 195.330 83.515 195.590 ;
        RECT 83.575 195.330 83.835 195.590 ;
        RECT 43.680 194.820 43.940 195.080 ;
        RECT 44.140 194.820 44.400 195.080 ;
        RECT 80.480 194.820 80.740 195.080 ;
        RECT 84.160 194.820 84.420 195.080 ;
        RECT 62.080 194.480 62.340 194.740 ;
        RECT 78.640 194.480 78.900 194.740 ;
        RECT 32.180 193.800 32.440 194.060 ;
        RECT 34.480 193.460 34.740 193.720 ;
        RECT 39.080 193.120 39.340 193.380 ;
        RECT 53.800 193.800 54.060 194.060 ;
        RECT 67.140 194.140 67.400 194.400 ;
        RECT 44.140 193.120 44.400 193.380 ;
        RECT 45.060 193.120 45.320 193.380 ;
        RECT 53.340 193.120 53.600 193.380 ;
        RECT 59.320 193.120 59.580 193.380 ;
        RECT 76.340 193.800 76.600 194.060 ;
        RECT 80.480 193.800 80.740 194.060 ;
        RECT 65.760 193.460 66.020 193.720 ;
        RECT 74.960 193.460 75.220 193.720 ;
        RECT 80.940 193.460 81.200 193.720 ;
        RECT 84.160 193.800 84.420 194.060 ;
        RECT 86.460 193.850 86.720 194.110 ;
        RECT 82.780 193.460 83.040 193.720 ;
        RECT 86.920 193.800 87.180 194.060 ;
        RECT 87.840 193.800 88.100 194.060 ;
        RECT 60.700 193.120 60.960 193.380 ;
        RECT 68.520 193.120 68.780 193.380 ;
        RECT 83.240 193.120 83.500 193.380 ;
        RECT 90.600 193.460 90.860 193.720 ;
        RECT 85.540 193.120 85.800 193.380 ;
        RECT 87.840 193.120 88.100 193.380 ;
        RECT 36.020 192.610 36.280 192.870 ;
        RECT 36.340 192.610 36.600 192.870 ;
        RECT 36.660 192.610 36.920 192.870 ;
        RECT 36.980 192.610 37.240 192.870 ;
        RECT 37.300 192.610 37.560 192.870 ;
        RECT 54.530 192.610 54.790 192.870 ;
        RECT 54.850 192.610 55.110 192.870 ;
        RECT 55.170 192.610 55.430 192.870 ;
        RECT 55.490 192.610 55.750 192.870 ;
        RECT 55.810 192.610 56.070 192.870 ;
        RECT 73.040 192.610 73.300 192.870 ;
        RECT 73.360 192.610 73.620 192.870 ;
        RECT 73.680 192.610 73.940 192.870 ;
        RECT 74.000 192.610 74.260 192.870 ;
        RECT 74.320 192.610 74.580 192.870 ;
        RECT 91.550 192.610 91.810 192.870 ;
        RECT 91.870 192.610 92.130 192.870 ;
        RECT 92.190 192.610 92.450 192.870 ;
        RECT 92.510 192.610 92.770 192.870 ;
        RECT 92.830 192.610 93.090 192.870 ;
        RECT 19.760 192.100 20.020 192.360 ;
        RECT 51.960 192.100 52.220 192.360 ;
        RECT 66.220 192.100 66.480 192.360 ;
        RECT 71.740 192.100 72.000 192.360 ;
        RECT 80.940 192.100 81.200 192.360 ;
        RECT 86.920 192.100 87.180 192.360 ;
        RECT 28.500 191.760 28.760 192.020 ;
        RECT 34.480 191.760 34.740 192.020 ;
        RECT 44.140 191.760 44.400 192.020 ;
        RECT 33.560 191.420 33.820 191.680 ;
        RECT 34.940 191.420 35.200 191.680 ;
        RECT 26.200 191.080 26.460 191.340 ;
        RECT 45.060 191.420 45.320 191.680 ;
        RECT 39.080 191.080 39.340 191.340 ;
        RECT 43.680 191.080 43.940 191.340 ;
        RECT 46.900 191.420 47.160 191.680 ;
        RECT 90.600 191.760 90.860 192.020 ;
        RECT 33.100 190.740 33.360 191.000 ;
        RECT 37.240 190.740 37.500 191.000 ;
        RECT 52.880 191.420 53.140 191.680 ;
        RECT 53.340 191.420 53.600 191.680 ;
        RECT 59.780 191.420 60.040 191.680 ;
        RECT 63.000 191.420 63.260 191.680 ;
        RECT 66.680 191.420 66.940 191.680 ;
        RECT 68.520 191.420 68.780 191.680 ;
        RECT 76.340 191.420 76.600 191.680 ;
        RECT 81.860 191.420 82.120 191.680 ;
        RECT 85.080 191.420 85.340 191.680 ;
        RECT 57.940 191.080 58.200 191.340 ;
        RECT 86.000 191.080 86.260 191.340 ;
        RECT 87.840 191.080 88.100 191.340 ;
        RECT 53.800 190.740 54.060 191.000 ;
        RECT 56.100 190.740 56.360 191.000 ;
        RECT 62.540 190.740 62.800 191.000 ;
        RECT 43.220 190.400 43.480 190.660 ;
        RECT 51.500 190.400 51.760 190.660 ;
        RECT 52.420 190.400 52.680 190.660 ;
        RECT 56.560 190.400 56.820 190.660 ;
        RECT 59.320 190.400 59.580 190.660 ;
        RECT 63.000 190.400 63.260 190.660 ;
        RECT 72.660 190.400 72.920 190.660 ;
        RECT 26.765 189.890 27.025 190.150 ;
        RECT 27.085 189.890 27.345 190.150 ;
        RECT 27.405 189.890 27.665 190.150 ;
        RECT 27.725 189.890 27.985 190.150 ;
        RECT 28.045 189.890 28.305 190.150 ;
        RECT 45.275 189.890 45.535 190.150 ;
        RECT 45.595 189.890 45.855 190.150 ;
        RECT 45.915 189.890 46.175 190.150 ;
        RECT 46.235 189.890 46.495 190.150 ;
        RECT 46.555 189.890 46.815 190.150 ;
        RECT 63.785 189.890 64.045 190.150 ;
        RECT 64.105 189.890 64.365 190.150 ;
        RECT 64.425 189.890 64.685 190.150 ;
        RECT 64.745 189.890 65.005 190.150 ;
        RECT 65.065 189.890 65.325 190.150 ;
        RECT 82.295 189.890 82.555 190.150 ;
        RECT 82.615 189.890 82.875 190.150 ;
        RECT 82.935 189.890 83.195 190.150 ;
        RECT 83.255 189.890 83.515 190.150 ;
        RECT 83.575 189.890 83.835 190.150 ;
        RECT 28.500 189.380 28.760 189.640 ;
        RECT 33.100 189.380 33.360 189.640 ;
        RECT 34.020 189.040 34.280 189.300 ;
        RECT 35.400 189.040 35.660 189.300 ;
        RECT 43.680 189.380 43.940 189.640 ;
        RECT 46.900 189.380 47.160 189.640 ;
        RECT 52.880 189.380 53.140 189.640 ;
        RECT 60.700 189.380 60.960 189.640 ;
        RECT 40.000 189.040 40.260 189.300 ;
        RECT 44.140 189.040 44.400 189.300 ;
        RECT 74.960 189.380 75.220 189.640 ;
        RECT 75.880 189.380 76.140 189.640 ;
        RECT 68.520 189.040 68.780 189.300 ;
        RECT 35.860 188.700 36.120 188.960 ;
        RECT 33.560 188.360 33.820 188.620 ;
        RECT 34.480 188.020 34.740 188.280 ;
        RECT 35.400 188.360 35.660 188.620 ;
        RECT 37.240 188.360 37.500 188.620 ;
        RECT 39.540 188.360 39.800 188.620 ;
        RECT 48.280 188.360 48.540 188.620 ;
        RECT 51.500 188.360 51.760 188.620 ;
        RECT 52.420 188.360 52.680 188.620 ;
        RECT 53.800 188.360 54.060 188.620 ;
        RECT 56.100 188.360 56.360 188.620 ;
        RECT 56.560 188.360 56.820 188.620 ;
        RECT 58.860 188.360 59.120 188.620 ;
        RECT 62.540 188.700 62.800 188.960 ;
        RECT 63.460 188.700 63.720 188.960 ;
        RECT 38.160 187.680 38.420 187.940 ;
        RECT 38.620 187.680 38.880 187.940 ;
        RECT 39.080 187.680 39.340 187.940 ;
        RECT 42.760 188.020 43.020 188.280 ;
        RECT 47.360 187.680 47.620 187.940 ;
        RECT 57.020 188.020 57.280 188.280 ;
        RECT 61.160 187.680 61.420 187.940 ;
        RECT 63.920 188.360 64.180 188.620 ;
        RECT 63.460 188.020 63.720 188.280 ;
        RECT 68.980 188.020 69.240 188.280 ;
        RECT 65.300 187.680 65.560 187.940 ;
        RECT 71.280 187.680 71.540 187.940 ;
        RECT 72.200 187.680 72.460 187.940 ;
        RECT 72.660 187.680 72.920 187.940 ;
        RECT 75.420 187.680 75.680 187.940 ;
        RECT 36.020 187.170 36.280 187.430 ;
        RECT 36.340 187.170 36.600 187.430 ;
        RECT 36.660 187.170 36.920 187.430 ;
        RECT 36.980 187.170 37.240 187.430 ;
        RECT 37.300 187.170 37.560 187.430 ;
        RECT 54.530 187.170 54.790 187.430 ;
        RECT 54.850 187.170 55.110 187.430 ;
        RECT 55.170 187.170 55.430 187.430 ;
        RECT 55.490 187.170 55.750 187.430 ;
        RECT 55.810 187.170 56.070 187.430 ;
        RECT 73.040 187.170 73.300 187.430 ;
        RECT 73.360 187.170 73.620 187.430 ;
        RECT 73.680 187.170 73.940 187.430 ;
        RECT 74.000 187.170 74.260 187.430 ;
        RECT 74.320 187.170 74.580 187.430 ;
        RECT 91.550 187.170 91.810 187.430 ;
        RECT 91.870 187.170 92.130 187.430 ;
        RECT 92.190 187.170 92.450 187.430 ;
        RECT 92.510 187.170 92.770 187.430 ;
        RECT 92.830 187.170 93.090 187.430 ;
        RECT 26.200 186.660 26.460 186.920 ;
        RECT 26.200 185.980 26.460 186.240 ;
        RECT 34.940 186.660 35.200 186.920 ;
        RECT 32.180 185.980 32.440 186.240 ;
        RECT 33.100 185.980 33.360 186.240 ;
        RECT 28.960 184.960 29.220 185.220 ;
        RECT 31.720 184.960 31.980 185.220 ;
        RECT 34.480 185.980 34.740 186.240 ;
        RECT 35.400 186.320 35.660 186.580 ;
        RECT 41.840 186.660 42.100 186.920 ;
        RECT 58.860 186.660 59.120 186.920 ;
        RECT 35.860 185.980 36.120 186.240 ;
        RECT 40.000 186.150 40.260 186.410 ;
        RECT 47.360 186.320 47.620 186.580 ;
        RECT 35.400 184.960 35.660 185.220 ;
        RECT 38.160 185.640 38.420 185.900 ;
        RECT 38.620 185.640 38.880 185.900 ;
        RECT 36.780 185.300 37.040 185.560 ;
        RECT 37.700 185.300 37.960 185.560 ;
        RECT 40.460 185.640 40.720 185.900 ;
        RECT 43.220 185.980 43.480 186.240 ;
        RECT 57.020 185.980 57.280 186.240 ;
        RECT 60.240 185.980 60.500 186.240 ;
        RECT 63.920 186.320 64.180 186.580 ;
        RECT 62.540 185.980 62.800 186.240 ;
        RECT 79.100 186.660 79.360 186.920 ;
        RECT 68.980 186.320 69.240 186.580 ;
        RECT 65.300 185.980 65.560 186.240 ;
        RECT 65.760 185.980 66.020 186.240 ;
        RECT 71.280 185.980 71.540 186.240 ;
        RECT 44.140 185.640 44.400 185.900 ;
        RECT 60.700 185.640 60.960 185.900 ;
        RECT 69.900 185.640 70.160 185.900 ;
        RECT 75.420 185.980 75.680 186.240 ;
        RECT 74.960 185.640 75.220 185.900 ;
        RECT 77.720 185.640 77.980 185.900 ;
        RECT 78.640 185.980 78.900 186.240 ;
        RECT 80.020 185.980 80.280 186.240 ;
        RECT 80.480 185.980 80.740 186.240 ;
        RECT 81.860 185.980 82.120 186.240 ;
        RECT 86.920 185.980 87.180 186.240 ;
        RECT 83.700 185.640 83.960 185.900 ;
        RECT 42.300 184.960 42.560 185.220 ;
        RECT 44.600 184.960 44.860 185.220 ;
        RECT 50.120 184.960 50.380 185.220 ;
        RECT 62.080 184.960 62.340 185.220 ;
        RECT 68.520 184.960 68.780 185.220 ;
        RECT 70.820 184.960 71.080 185.220 ;
        RECT 85.540 184.960 85.800 185.220 ;
        RECT 90.140 184.960 90.400 185.220 ;
        RECT 26.765 184.450 27.025 184.710 ;
        RECT 27.085 184.450 27.345 184.710 ;
        RECT 27.405 184.450 27.665 184.710 ;
        RECT 27.725 184.450 27.985 184.710 ;
        RECT 28.045 184.450 28.305 184.710 ;
        RECT 45.275 184.450 45.535 184.710 ;
        RECT 45.595 184.450 45.855 184.710 ;
        RECT 45.915 184.450 46.175 184.710 ;
        RECT 46.235 184.450 46.495 184.710 ;
        RECT 46.555 184.450 46.815 184.710 ;
        RECT 63.785 184.450 64.045 184.710 ;
        RECT 64.105 184.450 64.365 184.710 ;
        RECT 64.425 184.450 64.685 184.710 ;
        RECT 64.745 184.450 65.005 184.710 ;
        RECT 65.065 184.450 65.325 184.710 ;
        RECT 82.295 184.450 82.555 184.710 ;
        RECT 82.615 184.450 82.875 184.710 ;
        RECT 82.935 184.450 83.195 184.710 ;
        RECT 83.255 184.450 83.515 184.710 ;
        RECT 83.575 184.450 83.835 184.710 ;
        RECT 26.200 183.940 26.460 184.200 ;
        RECT 31.720 183.940 31.980 184.200 ;
        RECT 32.180 183.940 32.440 184.200 ;
        RECT 34.480 183.600 34.740 183.860 ;
        RECT 36.780 183.600 37.040 183.860 ;
        RECT 37.700 183.940 37.960 184.200 ;
        RECT 44.140 183.940 44.400 184.200 ;
        RECT 48.280 183.940 48.540 184.200 ;
        RECT 41.840 183.600 42.100 183.860 ;
        RECT 42.760 183.600 43.020 183.860 ;
        RECT 44.600 183.600 44.860 183.860 ;
        RECT 34.020 183.260 34.280 183.520 ;
        RECT 38.620 183.260 38.880 183.520 ;
        RECT 28.960 182.920 29.220 183.180 ;
        RECT 29.420 182.920 29.680 183.180 ;
        RECT 40.460 182.920 40.720 183.180 ;
        RECT 31.260 182.580 31.520 182.840 ;
        RECT 42.300 182.920 42.560 183.180 ;
        RECT 42.760 182.580 43.020 182.840 ;
        RECT 44.600 182.920 44.860 183.180 ;
        RECT 47.360 183.260 47.620 183.520 ;
        RECT 57.020 183.940 57.280 184.200 ;
        RECT 67.140 183.940 67.400 184.200 ;
        RECT 80.020 183.940 80.280 184.200 ;
        RECT 84.160 183.940 84.420 184.200 ;
        RECT 86.920 183.940 87.180 184.200 ;
        RECT 65.760 183.600 66.020 183.860 ;
        RECT 59.780 183.260 60.040 183.520 ;
        RECT 86.000 183.600 86.260 183.860 ;
        RECT 48.740 182.920 49.000 183.180 ;
        RECT 50.120 182.920 50.380 183.180 ;
        RECT 52.880 182.920 53.140 183.180 ;
        RECT 49.660 182.580 49.920 182.840 ;
        RECT 57.480 182.920 57.740 183.180 ;
        RECT 70.820 183.260 71.080 183.520 ;
        RECT 88.300 183.940 88.560 184.200 ;
        RECT 69.900 182.920 70.160 183.180 ;
        RECT 72.660 182.920 72.920 183.180 ;
        RECT 72.200 182.580 72.460 182.840 ;
        RECT 84.160 182.920 84.420 183.180 ;
        RECT 85.080 182.920 85.340 183.180 ;
        RECT 85.540 182.920 85.800 183.180 ;
        RECT 86.460 182.920 86.720 183.180 ;
        RECT 90.140 182.580 90.400 182.840 ;
        RECT 42.300 182.240 42.560 182.500 ;
        RECT 56.560 182.240 56.820 182.500 ;
        RECT 84.160 182.240 84.420 182.500 ;
        RECT 86.920 182.240 87.180 182.500 ;
        RECT 36.020 181.730 36.280 181.990 ;
        RECT 36.340 181.730 36.600 181.990 ;
        RECT 36.660 181.730 36.920 181.990 ;
        RECT 36.980 181.730 37.240 181.990 ;
        RECT 37.300 181.730 37.560 181.990 ;
        RECT 54.530 181.730 54.790 181.990 ;
        RECT 54.850 181.730 55.110 181.990 ;
        RECT 55.170 181.730 55.430 181.990 ;
        RECT 55.490 181.730 55.750 181.990 ;
        RECT 55.810 181.730 56.070 181.990 ;
        RECT 73.040 181.730 73.300 181.990 ;
        RECT 73.360 181.730 73.620 181.990 ;
        RECT 73.680 181.730 73.940 181.990 ;
        RECT 74.000 181.730 74.260 181.990 ;
        RECT 74.320 181.730 74.580 181.990 ;
        RECT 91.550 181.730 91.810 181.990 ;
        RECT 91.870 181.730 92.130 181.990 ;
        RECT 92.190 181.730 92.450 181.990 ;
        RECT 92.510 181.730 92.770 181.990 ;
        RECT 92.830 181.730 93.090 181.990 ;
        RECT 35.400 181.220 35.660 181.480 ;
        RECT 41.840 181.220 42.100 181.480 ;
        RECT 42.300 181.220 42.560 181.480 ;
        RECT 48.740 181.220 49.000 181.480 ;
        RECT 61.160 181.220 61.420 181.480 ;
        RECT 62.080 181.220 62.340 181.480 ;
        RECT 39.080 180.880 39.340 181.140 ;
        RECT 40.920 180.540 41.180 180.800 ;
        RECT 42.760 180.540 43.020 180.800 ;
        RECT 38.620 180.200 38.880 180.460 ;
        RECT 68.980 180.540 69.240 180.800 ;
        RECT 75.420 180.540 75.680 180.800 ;
        RECT 77.720 180.540 77.980 180.800 ;
        RECT 78.640 180.540 78.900 180.800 ;
        RECT 49.660 179.860 49.920 180.120 ;
        RECT 73.120 180.200 73.380 180.460 ;
        RECT 40.920 179.520 41.180 179.780 ;
        RECT 41.840 179.520 42.100 179.780 ;
        RECT 43.680 179.520 43.940 179.780 ;
        RECT 61.160 179.520 61.420 179.780 ;
        RECT 62.080 179.520 62.340 179.780 ;
        RECT 75.420 179.520 75.680 179.780 ;
        RECT 26.765 179.010 27.025 179.270 ;
        RECT 27.085 179.010 27.345 179.270 ;
        RECT 27.405 179.010 27.665 179.270 ;
        RECT 27.725 179.010 27.985 179.270 ;
        RECT 28.045 179.010 28.305 179.270 ;
        RECT 45.275 179.010 45.535 179.270 ;
        RECT 45.595 179.010 45.855 179.270 ;
        RECT 45.915 179.010 46.175 179.270 ;
        RECT 46.235 179.010 46.495 179.270 ;
        RECT 46.555 179.010 46.815 179.270 ;
        RECT 63.785 179.010 64.045 179.270 ;
        RECT 64.105 179.010 64.365 179.270 ;
        RECT 64.425 179.010 64.685 179.270 ;
        RECT 64.745 179.010 65.005 179.270 ;
        RECT 65.065 179.010 65.325 179.270 ;
        RECT 82.295 179.010 82.555 179.270 ;
        RECT 82.615 179.010 82.875 179.270 ;
        RECT 82.935 179.010 83.195 179.270 ;
        RECT 83.255 179.010 83.515 179.270 ;
        RECT 83.575 179.010 83.835 179.270 ;
        RECT 37.700 178.500 37.960 178.760 ;
        RECT 33.100 178.160 33.360 178.420 ;
        RECT 22.980 177.480 23.240 177.740 ;
        RECT 32.180 177.140 32.440 177.400 ;
        RECT 31.720 176.800 31.980 177.060 ;
        RECT 38.620 178.160 38.880 178.420 ;
        RECT 55.180 178.500 55.440 178.760 ;
        RECT 56.560 178.500 56.820 178.760 ;
        RECT 60.700 178.500 60.960 178.760 ;
        RECT 34.020 177.820 34.280 178.080 ;
        RECT 40.000 177.820 40.260 178.080 ;
        RECT 35.400 177.140 35.660 177.400 ;
        RECT 38.160 177.480 38.420 177.740 ;
        RECT 40.920 177.820 41.180 178.080 ;
        RECT 41.840 177.480 42.100 177.740 ;
        RECT 39.540 177.140 39.800 177.400 ;
        RECT 34.480 176.800 34.740 177.060 ;
        RECT 38.620 176.800 38.880 177.060 ;
        RECT 43.680 177.480 43.940 177.740 ;
        RECT 47.820 177.480 48.080 177.740 ;
        RECT 51.040 177.480 51.300 177.740 ;
        RECT 52.880 177.480 53.140 177.740 ;
        RECT 53.340 177.480 53.600 177.740 ;
        RECT 55.180 177.480 55.440 177.740 ;
        RECT 59.320 178.160 59.580 178.420 ;
        RECT 61.160 177.820 61.420 178.080 ;
        RECT 43.220 176.800 43.480 177.060 ;
        RECT 46.900 176.800 47.160 177.060 ;
        RECT 48.280 176.800 48.540 177.060 ;
        RECT 51.500 177.140 51.760 177.400 ;
        RECT 53.800 177.140 54.060 177.400 ;
        RECT 63.000 177.480 63.260 177.740 ;
        RECT 77.720 178.160 77.980 178.420 ;
        RECT 86.000 177.820 86.260 178.080 ;
        RECT 80.480 177.480 80.740 177.740 ;
        RECT 53.340 176.800 53.600 177.060 ;
        RECT 69.440 177.140 69.700 177.400 ;
        RECT 61.620 176.800 61.880 177.060 ;
        RECT 68.520 176.800 68.780 177.060 ;
        RECT 69.900 176.800 70.160 177.060 ;
        RECT 72.660 177.140 72.920 177.400 ;
        RECT 76.800 177.140 77.060 177.400 ;
        RECT 86.920 177.140 87.180 177.400 ;
        RECT 88.300 177.480 88.560 177.740 ;
        RECT 90.600 177.140 90.860 177.400 ;
        RECT 73.120 176.800 73.380 177.060 ;
        RECT 80.940 176.800 81.200 177.060 ;
        RECT 36.020 176.290 36.280 176.550 ;
        RECT 36.340 176.290 36.600 176.550 ;
        RECT 36.660 176.290 36.920 176.550 ;
        RECT 36.980 176.290 37.240 176.550 ;
        RECT 37.300 176.290 37.560 176.550 ;
        RECT 54.530 176.290 54.790 176.550 ;
        RECT 54.850 176.290 55.110 176.550 ;
        RECT 55.170 176.290 55.430 176.550 ;
        RECT 55.490 176.290 55.750 176.550 ;
        RECT 55.810 176.290 56.070 176.550 ;
        RECT 73.040 176.290 73.300 176.550 ;
        RECT 73.360 176.290 73.620 176.550 ;
        RECT 73.680 176.290 73.940 176.550 ;
        RECT 74.000 176.290 74.260 176.550 ;
        RECT 74.320 176.290 74.580 176.550 ;
        RECT 91.550 176.290 91.810 176.550 ;
        RECT 91.870 176.290 92.130 176.550 ;
        RECT 92.190 176.290 92.450 176.550 ;
        RECT 92.510 176.290 92.770 176.550 ;
        RECT 92.830 176.290 93.090 176.550 ;
        RECT 31.720 175.780 31.980 176.040 ;
        RECT 32.180 175.780 32.440 176.040 ;
        RECT 33.100 175.780 33.360 176.040 ;
        RECT 38.620 175.780 38.880 176.040 ;
        RECT 40.000 175.780 40.260 176.040 ;
        RECT 51.500 175.780 51.760 176.040 ;
        RECT 57.480 175.780 57.740 176.040 ;
        RECT 61.620 175.780 61.880 176.040 ;
        RECT 62.080 175.780 62.340 176.040 ;
        RECT 65.760 175.780 66.020 176.040 ;
        RECT 68.980 175.780 69.240 176.040 ;
        RECT 72.660 175.780 72.920 176.040 ;
        RECT 33.560 175.100 33.820 175.360 ;
        RECT 35.400 175.100 35.660 175.360 ;
        RECT 37.700 175.100 37.960 175.360 ;
        RECT 29.880 174.760 30.140 175.020 ;
        RECT 34.480 174.760 34.740 175.020 ;
        RECT 43.220 175.440 43.480 175.700 ;
        RECT 46.900 175.440 47.160 175.700 ;
        RECT 51.960 175.440 52.220 175.700 ;
        RECT 44.600 174.760 44.860 175.020 ;
        RECT 63.920 175.100 64.180 175.360 ;
        RECT 65.300 175.100 65.560 175.360 ;
        RECT 66.680 175.440 66.940 175.700 ;
        RECT 80.020 175.780 80.280 176.040 ;
        RECT 80.940 175.780 81.200 176.040 ;
        RECT 68.520 175.100 68.780 175.360 ;
        RECT 69.440 175.100 69.700 175.360 ;
        RECT 69.900 175.100 70.160 175.360 ;
        RECT 75.420 175.100 75.680 175.360 ;
        RECT 34.020 174.420 34.280 174.680 ;
        RECT 44.140 174.420 44.400 174.680 ;
        RECT 25.280 174.080 25.540 174.340 ;
        RECT 40.920 174.080 41.180 174.340 ;
        RECT 53.340 174.080 53.600 174.340 ;
        RECT 61.160 174.080 61.420 174.340 ;
        RECT 77.720 175.100 77.980 175.360 ;
        RECT 65.300 174.420 65.560 174.680 ;
        RECT 66.220 174.080 66.480 174.340 ;
        RECT 68.980 174.420 69.240 174.680 ;
        RECT 71.740 174.420 72.000 174.680 ;
        RECT 78.640 175.100 78.900 175.360 ;
        RECT 88.300 175.780 88.560 176.040 ;
        RECT 80.020 174.760 80.280 175.020 ;
        RECT 80.480 174.760 80.740 175.020 ;
        RECT 86.000 174.080 86.260 174.340 ;
        RECT 90.600 174.080 90.860 174.340 ;
        RECT 26.765 173.570 27.025 173.830 ;
        RECT 27.085 173.570 27.345 173.830 ;
        RECT 27.405 173.570 27.665 173.830 ;
        RECT 27.725 173.570 27.985 173.830 ;
        RECT 28.045 173.570 28.305 173.830 ;
        RECT 45.275 173.570 45.535 173.830 ;
        RECT 45.595 173.570 45.855 173.830 ;
        RECT 45.915 173.570 46.175 173.830 ;
        RECT 46.235 173.570 46.495 173.830 ;
        RECT 46.555 173.570 46.815 173.830 ;
        RECT 63.785 173.570 64.045 173.830 ;
        RECT 64.105 173.570 64.365 173.830 ;
        RECT 64.425 173.570 64.685 173.830 ;
        RECT 64.745 173.570 65.005 173.830 ;
        RECT 65.065 173.570 65.325 173.830 ;
        RECT 82.295 173.570 82.555 173.830 ;
        RECT 82.615 173.570 82.875 173.830 ;
        RECT 82.935 173.570 83.195 173.830 ;
        RECT 83.255 173.570 83.515 173.830 ;
        RECT 83.575 173.570 83.835 173.830 ;
        RECT 29.880 173.060 30.140 173.320 ;
        RECT 22.980 172.040 23.240 172.300 ;
        RECT 28.960 172.040 29.220 172.300 ;
        RECT 35.860 172.720 36.120 172.980 ;
        RECT 41.840 173.060 42.100 173.320 ;
        RECT 47.820 173.060 48.080 173.320 ;
        RECT 71.740 173.060 72.000 173.320 ;
        RECT 80.020 173.060 80.280 173.320 ;
        RECT 43.680 172.720 43.940 172.980 ;
        RECT 77.260 172.720 77.520 172.980 ;
        RECT 37.700 172.380 37.960 172.640 ;
        RECT 47.360 172.380 47.620 172.640 ;
        RECT 61.620 172.380 61.880 172.640 ;
        RECT 38.160 172.040 38.420 172.300 ;
        RECT 39.540 172.040 39.800 172.300 ;
        RECT 41.380 172.040 41.640 172.300 ;
        RECT 48.280 172.040 48.540 172.300 ;
        RECT 52.420 172.040 52.680 172.300 ;
        RECT 31.260 171.700 31.520 171.960 ;
        RECT 34.020 171.700 34.280 171.960 ;
        RECT 34.480 171.700 34.740 171.960 ;
        RECT 32.640 171.360 32.900 171.620 ;
        RECT 39.080 171.360 39.340 171.620 ;
        RECT 40.000 171.360 40.260 171.620 ;
        RECT 59.320 172.040 59.580 172.300 ;
        RECT 59.780 172.040 60.040 172.300 ;
        RECT 60.240 172.040 60.500 172.300 ;
        RECT 61.160 172.040 61.420 172.300 ;
        RECT 63.000 171.700 63.260 171.960 ;
        RECT 66.220 172.040 66.480 172.300 ;
        RECT 78.640 172.040 78.900 172.300 ;
        RECT 81.400 172.040 81.660 172.300 ;
        RECT 86.920 172.040 87.180 172.300 ;
        RECT 43.680 171.360 43.940 171.620 ;
        RECT 56.560 171.360 56.820 171.620 ;
        RECT 57.940 171.360 58.200 171.620 ;
        RECT 60.700 171.360 60.960 171.620 ;
        RECT 75.420 171.360 75.680 171.620 ;
        RECT 85.080 171.360 85.340 171.620 ;
        RECT 36.020 170.850 36.280 171.110 ;
        RECT 36.340 170.850 36.600 171.110 ;
        RECT 36.660 170.850 36.920 171.110 ;
        RECT 36.980 170.850 37.240 171.110 ;
        RECT 37.300 170.850 37.560 171.110 ;
        RECT 54.530 170.850 54.790 171.110 ;
        RECT 54.850 170.850 55.110 171.110 ;
        RECT 55.170 170.850 55.430 171.110 ;
        RECT 55.490 170.850 55.750 171.110 ;
        RECT 55.810 170.850 56.070 171.110 ;
        RECT 73.040 170.850 73.300 171.110 ;
        RECT 73.360 170.850 73.620 171.110 ;
        RECT 73.680 170.850 73.940 171.110 ;
        RECT 74.000 170.850 74.260 171.110 ;
        RECT 74.320 170.850 74.580 171.110 ;
        RECT 91.550 170.850 91.810 171.110 ;
        RECT 91.870 170.850 92.130 171.110 ;
        RECT 92.190 170.850 92.450 171.110 ;
        RECT 92.510 170.850 92.770 171.110 ;
        RECT 92.830 170.850 93.090 171.110 ;
        RECT 25.280 170.340 25.540 170.600 ;
        RECT 32.640 170.340 32.900 170.600 ;
        RECT 63.000 170.340 63.260 170.600 ;
        RECT 66.680 170.340 66.940 170.600 ;
        RECT 67.600 170.340 67.860 170.600 ;
        RECT 29.420 170.000 29.680 170.260 ;
        RECT 40.460 170.000 40.720 170.260 ;
        RECT 43.680 170.000 43.940 170.260 ;
        RECT 39.080 169.660 39.340 169.920 ;
        RECT 52.420 169.660 52.680 169.920 ;
        RECT 53.800 169.660 54.060 169.920 ;
        RECT 58.400 169.660 58.660 169.920 ;
        RECT 60.700 169.660 60.960 169.920 ;
        RECT 75.880 170.000 76.140 170.260 ;
        RECT 78.640 170.000 78.900 170.260 ;
        RECT 68.520 169.660 68.780 169.920 ;
        RECT 72.200 169.660 72.460 169.920 ;
        RECT 75.420 169.660 75.680 169.920 ;
        RECT 35.860 169.320 36.120 169.580 ;
        RECT 38.620 169.320 38.880 169.580 ;
        RECT 40.000 169.320 40.260 169.580 ;
        RECT 74.960 169.320 75.220 169.580 ;
        RECT 78.180 169.660 78.440 169.920 ;
        RECT 81.400 170.000 81.660 170.260 ;
        RECT 80.940 169.660 81.200 169.920 ;
        RECT 28.960 168.980 29.220 169.240 ;
        RECT 32.180 168.980 32.440 169.240 ;
        RECT 44.600 168.980 44.860 169.240 ;
        RECT 79.100 169.320 79.360 169.580 ;
        RECT 79.560 168.980 79.820 169.240 ;
        RECT 38.160 168.640 38.420 168.900 ;
        RECT 62.080 168.640 62.340 168.900 ;
        RECT 66.680 168.640 66.940 168.900 ;
        RECT 77.260 168.640 77.520 168.900 ;
        RECT 78.640 168.640 78.900 168.900 ;
        RECT 85.540 168.640 85.800 168.900 ;
        RECT 26.765 168.130 27.025 168.390 ;
        RECT 27.085 168.130 27.345 168.390 ;
        RECT 27.405 168.130 27.665 168.390 ;
        RECT 27.725 168.130 27.985 168.390 ;
        RECT 28.045 168.130 28.305 168.390 ;
        RECT 45.275 168.130 45.535 168.390 ;
        RECT 45.595 168.130 45.855 168.390 ;
        RECT 45.915 168.130 46.175 168.390 ;
        RECT 46.235 168.130 46.495 168.390 ;
        RECT 46.555 168.130 46.815 168.390 ;
        RECT 63.785 168.130 64.045 168.390 ;
        RECT 64.105 168.130 64.365 168.390 ;
        RECT 64.425 168.130 64.685 168.390 ;
        RECT 64.745 168.130 65.005 168.390 ;
        RECT 65.065 168.130 65.325 168.390 ;
        RECT 82.295 168.130 82.555 168.390 ;
        RECT 82.615 168.130 82.875 168.390 ;
        RECT 82.935 168.130 83.195 168.390 ;
        RECT 83.255 168.130 83.515 168.390 ;
        RECT 83.575 168.130 83.835 168.390 ;
        RECT 37.700 167.620 37.960 167.880 ;
        RECT 39.540 167.620 39.800 167.880 ;
        RECT 53.800 167.620 54.060 167.880 ;
        RECT 29.880 167.280 30.140 167.540 ;
        RECT 47.360 167.280 47.620 167.540 ;
        RECT 35.860 166.940 36.120 167.200 ;
        RECT 70.360 167.620 70.620 167.880 ;
        RECT 76.800 167.620 77.060 167.880 ;
        RECT 80.940 167.620 81.200 167.880 ;
        RECT 29.880 165.920 30.140 166.180 ;
        RECT 34.940 165.920 35.200 166.180 ;
        RECT 38.620 166.600 38.880 166.860 ;
        RECT 39.080 166.600 39.340 166.860 ;
        RECT 44.600 166.600 44.860 166.860 ;
        RECT 42.300 166.260 42.560 166.520 ;
        RECT 52.880 166.260 53.140 166.520 ;
        RECT 54.260 166.600 54.520 166.860 ;
        RECT 56.560 166.600 56.820 166.860 ;
        RECT 62.540 166.600 62.800 166.860 ;
        RECT 66.220 167.280 66.480 167.540 ;
        RECT 66.680 167.280 66.940 167.540 ;
        RECT 38.160 165.920 38.420 166.180 ;
        RECT 40.000 165.920 40.260 166.180 ;
        RECT 53.340 165.920 53.600 166.180 ;
        RECT 63.000 165.920 63.260 166.180 ;
        RECT 68.060 166.600 68.320 166.860 ;
        RECT 72.660 166.600 72.920 166.860 ;
        RECT 68.520 166.260 68.780 166.520 ;
        RECT 70.820 166.260 71.080 166.520 ;
        RECT 71.740 165.920 72.000 166.180 ;
        RECT 76.800 165.920 77.060 166.180 ;
        RECT 77.720 166.600 77.980 166.860 ;
        RECT 85.080 166.600 85.340 166.860 ;
        RECT 85.540 166.600 85.800 166.860 ;
        RECT 86.460 166.600 86.720 166.860 ;
        RECT 90.600 166.600 90.860 166.860 ;
        RECT 78.180 166.260 78.440 166.520 ;
        RECT 79.100 165.920 79.360 166.180 ;
        RECT 83.700 165.920 83.960 166.180 ;
        RECT 36.020 165.410 36.280 165.670 ;
        RECT 36.340 165.410 36.600 165.670 ;
        RECT 36.660 165.410 36.920 165.670 ;
        RECT 36.980 165.410 37.240 165.670 ;
        RECT 37.300 165.410 37.560 165.670 ;
        RECT 54.530 165.410 54.790 165.670 ;
        RECT 54.850 165.410 55.110 165.670 ;
        RECT 55.170 165.410 55.430 165.670 ;
        RECT 55.490 165.410 55.750 165.670 ;
        RECT 55.810 165.410 56.070 165.670 ;
        RECT 73.040 165.410 73.300 165.670 ;
        RECT 73.360 165.410 73.620 165.670 ;
        RECT 73.680 165.410 73.940 165.670 ;
        RECT 74.000 165.410 74.260 165.670 ;
        RECT 74.320 165.410 74.580 165.670 ;
        RECT 91.550 165.410 91.810 165.670 ;
        RECT 91.870 165.410 92.130 165.670 ;
        RECT 92.190 165.410 92.450 165.670 ;
        RECT 92.510 165.410 92.770 165.670 ;
        RECT 92.830 165.410 93.090 165.670 ;
        RECT 33.560 164.900 33.820 165.160 ;
        RECT 29.880 164.560 30.140 164.820 ;
        RECT 29.420 164.220 29.680 164.480 ;
        RECT 34.480 164.220 34.740 164.480 ;
        RECT 34.940 164.220 35.200 164.480 ;
        RECT 39.080 164.560 39.340 164.820 ;
        RECT 42.300 164.900 42.560 165.160 ;
        RECT 53.340 164.900 53.600 165.160 ;
        RECT 53.800 164.900 54.060 165.160 ;
        RECT 63.000 164.900 63.260 165.160 ;
        RECT 70.820 164.900 71.080 165.160 ;
        RECT 77.720 164.900 77.980 165.160 ;
        RECT 78.180 164.900 78.440 165.160 ;
        RECT 29.420 163.200 29.680 163.460 ;
        RECT 36.320 163.200 36.580 163.460 ;
        RECT 38.160 163.880 38.420 164.140 ;
        RECT 44.600 164.220 44.860 164.480 ;
        RECT 47.360 164.220 47.620 164.480 ;
        RECT 48.740 164.220 49.000 164.480 ;
        RECT 72.660 164.560 72.920 164.820 ;
        RECT 57.940 164.220 58.200 164.480 ;
        RECT 87.840 164.560 88.100 164.820 ;
        RECT 80.480 164.220 80.740 164.480 ;
        RECT 83.700 164.220 83.960 164.480 ;
        RECT 90.600 164.220 90.860 164.480 ;
        RECT 49.200 163.540 49.460 163.800 ;
        RECT 37.700 163.200 37.960 163.460 ;
        RECT 44.140 163.200 44.400 163.460 ;
        RECT 46.900 163.200 47.160 163.460 ;
        RECT 59.780 163.540 60.040 163.800 ;
        RECT 78.640 163.540 78.900 163.800 ;
        RECT 79.100 163.200 79.360 163.460 ;
        RECT 79.560 163.200 79.820 163.460 ;
        RECT 26.765 162.690 27.025 162.950 ;
        RECT 27.085 162.690 27.345 162.950 ;
        RECT 27.405 162.690 27.665 162.950 ;
        RECT 27.725 162.690 27.985 162.950 ;
        RECT 28.045 162.690 28.305 162.950 ;
        RECT 45.275 162.690 45.535 162.950 ;
        RECT 45.595 162.690 45.855 162.950 ;
        RECT 45.915 162.690 46.175 162.950 ;
        RECT 46.235 162.690 46.495 162.950 ;
        RECT 46.555 162.690 46.815 162.950 ;
        RECT 63.785 162.690 64.045 162.950 ;
        RECT 64.105 162.690 64.365 162.950 ;
        RECT 64.425 162.690 64.685 162.950 ;
        RECT 64.745 162.690 65.005 162.950 ;
        RECT 65.065 162.690 65.325 162.950 ;
        RECT 82.295 162.690 82.555 162.950 ;
        RECT 82.615 162.690 82.875 162.950 ;
        RECT 82.935 162.690 83.195 162.950 ;
        RECT 83.255 162.690 83.515 162.950 ;
        RECT 83.575 162.690 83.835 162.950 ;
        RECT 29.420 162.180 29.680 162.440 ;
        RECT 36.320 162.180 36.580 162.440 ;
        RECT 22.520 161.500 22.780 161.760 ;
        RECT 38.160 162.180 38.420 162.440 ;
        RECT 49.200 162.180 49.460 162.440 ;
        RECT 65.760 162.180 66.020 162.440 ;
        RECT 70.360 162.180 70.620 162.440 ;
        RECT 86.920 162.180 87.180 162.440 ;
        RECT 43.220 161.840 43.480 162.100 ;
        RECT 47.360 161.840 47.620 162.100 ;
        RECT 48.740 161.840 49.000 162.100 ;
        RECT 64.380 161.840 64.640 162.100 ;
        RECT 33.560 161.160 33.820 161.420 ;
        RECT 37.700 161.160 37.960 161.420 ;
        RECT 38.160 161.160 38.420 161.420 ;
        RECT 39.080 161.160 39.340 161.420 ;
        RECT 54.720 161.500 54.980 161.760 ;
        RECT 66.680 161.840 66.940 162.100 ;
        RECT 75.880 161.840 76.140 162.100 ;
        RECT 77.720 161.840 77.980 162.100 ;
        RECT 90.600 161.840 90.860 162.100 ;
        RECT 45.520 161.160 45.780 161.420 ;
        RECT 45.980 161.160 46.240 161.420 ;
        RECT 46.900 161.160 47.160 161.420 ;
        RECT 52.420 161.160 52.680 161.420 ;
        RECT 49.200 160.820 49.460 161.080 ;
        RECT 57.940 161.160 58.200 161.420 ;
        RECT 60.700 161.160 60.960 161.420 ;
        RECT 29.880 160.480 30.140 160.740 ;
        RECT 34.940 160.480 35.200 160.740 ;
        RECT 44.140 160.480 44.400 160.740 ;
        RECT 48.740 160.480 49.000 160.740 ;
        RECT 49.660 160.480 49.920 160.740 ;
        RECT 54.720 160.480 54.980 160.740 ;
        RECT 60.700 160.480 60.960 160.740 ;
        RECT 61.160 160.480 61.420 160.740 ;
        RECT 63.920 161.160 64.180 161.420 ;
        RECT 64.380 161.160 64.640 161.420 ;
        RECT 65.760 161.160 66.020 161.420 ;
        RECT 66.680 160.820 66.940 161.080 ;
        RECT 71.740 161.160 72.000 161.420 ;
        RECT 72.660 161.160 72.920 161.420 ;
        RECT 77.260 161.160 77.520 161.420 ;
        RECT 87.840 161.160 88.100 161.420 ;
        RECT 67.140 160.480 67.400 160.740 ;
        RECT 71.280 160.480 71.540 160.740 ;
        RECT 72.200 160.480 72.460 160.740 ;
        RECT 78.180 160.480 78.440 160.740 ;
        RECT 79.560 160.480 79.820 160.740 ;
        RECT 88.300 160.480 88.560 160.740 ;
        RECT 36.020 159.970 36.280 160.230 ;
        RECT 36.340 159.970 36.600 160.230 ;
        RECT 36.660 159.970 36.920 160.230 ;
        RECT 36.980 159.970 37.240 160.230 ;
        RECT 37.300 159.970 37.560 160.230 ;
        RECT 54.530 159.970 54.790 160.230 ;
        RECT 54.850 159.970 55.110 160.230 ;
        RECT 55.170 159.970 55.430 160.230 ;
        RECT 55.490 159.970 55.750 160.230 ;
        RECT 55.810 159.970 56.070 160.230 ;
        RECT 73.040 159.970 73.300 160.230 ;
        RECT 73.360 159.970 73.620 160.230 ;
        RECT 73.680 159.970 73.940 160.230 ;
        RECT 74.000 159.970 74.260 160.230 ;
        RECT 74.320 159.970 74.580 160.230 ;
        RECT 91.550 159.970 91.810 160.230 ;
        RECT 91.870 159.970 92.130 160.230 ;
        RECT 92.190 159.970 92.450 160.230 ;
        RECT 92.510 159.970 92.770 160.230 ;
        RECT 92.830 159.970 93.090 160.230 ;
        RECT 34.940 159.460 35.200 159.720 ;
        RECT 35.400 159.460 35.660 159.720 ;
        RECT 34.020 159.120 34.280 159.380 ;
        RECT 33.560 158.780 33.820 159.040 ;
        RECT 45.520 159.460 45.780 159.720 ;
        RECT 48.280 159.460 48.540 159.720 ;
        RECT 49.660 159.460 49.920 159.720 ;
        RECT 52.420 159.460 52.680 159.720 ;
        RECT 61.620 159.460 61.880 159.720 ;
        RECT 64.380 159.460 64.640 159.720 ;
        RECT 72.200 159.460 72.460 159.720 ;
        RECT 76.340 159.460 76.600 159.720 ;
        RECT 39.080 158.780 39.340 159.040 ;
        RECT 44.140 158.780 44.400 159.040 ;
        RECT 45.520 158.780 45.780 159.040 ;
        RECT 45.980 158.440 46.240 158.700 ;
        RECT 47.360 158.780 47.620 159.040 ;
        RECT 48.740 158.780 49.000 159.040 ;
        RECT 57.480 159.120 57.740 159.380 ;
        RECT 52.880 158.780 53.140 159.040 ;
        RECT 60.700 158.780 60.960 159.040 ;
        RECT 49.200 158.440 49.460 158.700 ;
        RECT 67.140 158.440 67.400 158.700 ;
        RECT 71.280 158.440 71.540 158.700 ;
        RECT 75.880 158.780 76.140 159.040 ;
        RECT 78.180 158.780 78.440 159.040 ;
        RECT 80.480 158.440 80.740 158.700 ;
        RECT 34.020 157.760 34.280 158.020 ;
        RECT 41.840 157.760 42.100 158.020 ;
        RECT 49.200 157.760 49.460 158.020 ;
        RECT 54.260 157.760 54.520 158.020 ;
        RECT 73.580 157.760 73.840 158.020 ;
        RECT 87.840 157.760 88.100 158.020 ;
        RECT 26.765 157.250 27.025 157.510 ;
        RECT 27.085 157.250 27.345 157.510 ;
        RECT 27.405 157.250 27.665 157.510 ;
        RECT 27.725 157.250 27.985 157.510 ;
        RECT 28.045 157.250 28.305 157.510 ;
        RECT 45.275 157.250 45.535 157.510 ;
        RECT 45.595 157.250 45.855 157.510 ;
        RECT 45.915 157.250 46.175 157.510 ;
        RECT 46.235 157.250 46.495 157.510 ;
        RECT 46.555 157.250 46.815 157.510 ;
        RECT 63.785 157.250 64.045 157.510 ;
        RECT 64.105 157.250 64.365 157.510 ;
        RECT 64.425 157.250 64.685 157.510 ;
        RECT 64.745 157.250 65.005 157.510 ;
        RECT 65.065 157.250 65.325 157.510 ;
        RECT 82.295 157.250 82.555 157.510 ;
        RECT 82.615 157.250 82.875 157.510 ;
        RECT 82.935 157.250 83.195 157.510 ;
        RECT 83.255 157.250 83.515 157.510 ;
        RECT 83.575 157.250 83.835 157.510 ;
        RECT 39.080 156.740 39.340 157.000 ;
        RECT 46.900 156.740 47.160 157.000 ;
        RECT 49.200 156.740 49.460 157.000 ;
        RECT 67.140 156.740 67.400 157.000 ;
        RECT 79.100 156.740 79.360 157.000 ;
        RECT 88.300 156.740 88.560 157.000 ;
        RECT 32.180 156.060 32.440 156.320 ;
        RECT 41.840 155.720 42.100 155.980 ;
        RECT 55.180 155.720 55.440 155.980 ;
        RECT 63.000 155.720 63.260 155.980 ;
        RECT 80.480 156.060 80.740 156.320 ;
        RECT 73.580 155.720 73.840 155.980 ;
        RECT 34.020 155.380 34.280 155.640 ;
        RECT 62.080 155.380 62.340 155.640 ;
        RECT 117.400 155.300 118.000 155.900 ;
        RECT 36.020 154.530 36.280 154.790 ;
        RECT 36.340 154.530 36.600 154.790 ;
        RECT 36.660 154.530 36.920 154.790 ;
        RECT 36.980 154.530 37.240 154.790 ;
        RECT 37.300 154.530 37.560 154.790 ;
        RECT 54.530 154.530 54.790 154.790 ;
        RECT 54.850 154.530 55.110 154.790 ;
        RECT 55.170 154.530 55.430 154.790 ;
        RECT 55.490 154.530 55.750 154.790 ;
        RECT 55.810 154.530 56.070 154.790 ;
        RECT 73.040 154.530 73.300 154.790 ;
        RECT 73.360 154.530 73.620 154.790 ;
        RECT 73.680 154.530 73.940 154.790 ;
        RECT 74.000 154.530 74.260 154.790 ;
        RECT 74.320 154.530 74.580 154.790 ;
        RECT 91.550 154.530 91.810 154.790 ;
        RECT 91.870 154.530 92.130 154.790 ;
        RECT 92.190 154.530 92.450 154.790 ;
        RECT 92.510 154.530 92.770 154.790 ;
        RECT 92.830 154.530 93.090 154.790 ;
        RECT 26.765 151.810 27.025 152.070 ;
        RECT 27.085 151.810 27.345 152.070 ;
        RECT 27.405 151.810 27.665 152.070 ;
        RECT 27.725 151.810 27.985 152.070 ;
        RECT 28.045 151.810 28.305 152.070 ;
        RECT 45.275 151.810 45.535 152.070 ;
        RECT 45.595 151.810 45.855 152.070 ;
        RECT 45.915 151.810 46.175 152.070 ;
        RECT 46.235 151.810 46.495 152.070 ;
        RECT 46.555 151.810 46.815 152.070 ;
        RECT 63.785 151.810 64.045 152.070 ;
        RECT 64.105 151.810 64.365 152.070 ;
        RECT 64.425 151.810 64.685 152.070 ;
        RECT 64.745 151.810 65.005 152.070 ;
        RECT 65.065 151.810 65.325 152.070 ;
        RECT 82.295 151.810 82.555 152.070 ;
        RECT 82.615 151.810 82.875 152.070 ;
        RECT 82.935 151.810 83.195 152.070 ;
        RECT 83.255 151.810 83.515 152.070 ;
        RECT 83.575 151.810 83.835 152.070 ;
        RECT 77.260 151.300 77.520 151.560 ;
        RECT 79.560 151.300 79.820 151.560 ;
        RECT 63.000 150.620 63.260 150.880 ;
        RECT 65.300 150.620 65.560 150.880 ;
        RECT 36.020 149.090 36.280 149.350 ;
        RECT 36.340 149.090 36.600 149.350 ;
        RECT 36.660 149.090 36.920 149.350 ;
        RECT 36.980 149.090 37.240 149.350 ;
        RECT 37.300 149.090 37.560 149.350 ;
        RECT 54.530 149.090 54.790 149.350 ;
        RECT 54.850 149.090 55.110 149.350 ;
        RECT 55.170 149.090 55.430 149.350 ;
        RECT 55.490 149.090 55.750 149.350 ;
        RECT 55.810 149.090 56.070 149.350 ;
        RECT 73.040 149.090 73.300 149.350 ;
        RECT 73.360 149.090 73.620 149.350 ;
        RECT 73.680 149.090 73.940 149.350 ;
        RECT 74.000 149.090 74.260 149.350 ;
        RECT 74.320 149.090 74.580 149.350 ;
        RECT 91.550 149.090 91.810 149.350 ;
        RECT 91.870 149.090 92.130 149.350 ;
        RECT 92.190 149.090 92.450 149.350 ;
        RECT 92.510 149.090 92.770 149.350 ;
        RECT 92.830 149.090 93.090 149.350 ;
        RECT 115.900 152.500 116.500 153.100 ;
        RECT 118.900 155.200 119.500 155.800 ;
        RECT 120.400 155.100 121.000 155.700 ;
        RECT 121.800 154.100 122.400 154.700 ;
        RECT 26.765 146.370 27.025 146.630 ;
        RECT 27.085 146.370 27.345 146.630 ;
        RECT 27.405 146.370 27.665 146.630 ;
        RECT 27.725 146.370 27.985 146.630 ;
        RECT 28.045 146.370 28.305 146.630 ;
        RECT 45.275 146.370 45.535 146.630 ;
        RECT 45.595 146.370 45.855 146.630 ;
        RECT 45.915 146.370 46.175 146.630 ;
        RECT 46.235 146.370 46.495 146.630 ;
        RECT 46.555 146.370 46.815 146.630 ;
        RECT 63.785 146.370 64.045 146.630 ;
        RECT 64.105 146.370 64.365 146.630 ;
        RECT 64.425 146.370 64.685 146.630 ;
        RECT 64.745 146.370 65.005 146.630 ;
        RECT 65.065 146.370 65.325 146.630 ;
        RECT 82.295 146.370 82.555 146.630 ;
        RECT 82.615 146.370 82.875 146.630 ;
        RECT 82.935 146.370 83.195 146.630 ;
        RECT 83.255 146.370 83.515 146.630 ;
        RECT 83.575 146.370 83.835 146.630 ;
        RECT 36.020 143.650 36.280 143.910 ;
        RECT 36.340 143.650 36.600 143.910 ;
        RECT 36.660 143.650 36.920 143.910 ;
        RECT 36.980 143.650 37.240 143.910 ;
        RECT 37.300 143.650 37.560 143.910 ;
        RECT 54.530 143.650 54.790 143.910 ;
        RECT 54.850 143.650 55.110 143.910 ;
        RECT 55.170 143.650 55.430 143.910 ;
        RECT 55.490 143.650 55.750 143.910 ;
        RECT 55.810 143.650 56.070 143.910 ;
        RECT 73.040 143.650 73.300 143.910 ;
        RECT 73.360 143.650 73.620 143.910 ;
        RECT 73.680 143.650 73.940 143.910 ;
        RECT 74.000 143.650 74.260 143.910 ;
        RECT 74.320 143.650 74.580 143.910 ;
        RECT 91.550 143.650 91.810 143.910 ;
        RECT 91.870 143.650 92.130 143.910 ;
        RECT 92.190 143.650 92.450 143.910 ;
        RECT 92.510 143.650 92.770 143.910 ;
        RECT 92.830 143.650 93.090 143.910 ;
        RECT 26.765 140.930 27.025 141.190 ;
        RECT 27.085 140.930 27.345 141.190 ;
        RECT 27.405 140.930 27.665 141.190 ;
        RECT 27.725 140.930 27.985 141.190 ;
        RECT 28.045 140.930 28.305 141.190 ;
        RECT 45.275 140.930 45.535 141.190 ;
        RECT 45.595 140.930 45.855 141.190 ;
        RECT 45.915 140.930 46.175 141.190 ;
        RECT 46.235 140.930 46.495 141.190 ;
        RECT 46.555 140.930 46.815 141.190 ;
        RECT 63.785 140.930 64.045 141.190 ;
        RECT 64.105 140.930 64.365 141.190 ;
        RECT 64.425 140.930 64.685 141.190 ;
        RECT 64.745 140.930 65.005 141.190 ;
        RECT 65.065 140.930 65.325 141.190 ;
        RECT 82.295 140.930 82.555 141.190 ;
        RECT 82.615 140.930 82.875 141.190 ;
        RECT 82.935 140.930 83.195 141.190 ;
        RECT 83.255 140.930 83.515 141.190 ;
        RECT 83.575 140.930 83.835 141.190 ;
        RECT 36.020 138.210 36.280 138.470 ;
        RECT 36.340 138.210 36.600 138.470 ;
        RECT 36.660 138.210 36.920 138.470 ;
        RECT 36.980 138.210 37.240 138.470 ;
        RECT 37.300 138.210 37.560 138.470 ;
        RECT 54.530 138.210 54.790 138.470 ;
        RECT 54.850 138.210 55.110 138.470 ;
        RECT 55.170 138.210 55.430 138.470 ;
        RECT 55.490 138.210 55.750 138.470 ;
        RECT 55.810 138.210 56.070 138.470 ;
        RECT 73.040 138.210 73.300 138.470 ;
        RECT 73.360 138.210 73.620 138.470 ;
        RECT 73.680 138.210 73.940 138.470 ;
        RECT 74.000 138.210 74.260 138.470 ;
        RECT 74.320 138.210 74.580 138.470 ;
        RECT 91.550 138.210 91.810 138.470 ;
        RECT 91.870 138.210 92.130 138.470 ;
        RECT 92.190 138.210 92.450 138.470 ;
        RECT 92.510 138.210 92.770 138.470 ;
        RECT 92.830 138.210 93.090 138.470 ;
        RECT 26.765 135.490 27.025 135.750 ;
        RECT 27.085 135.490 27.345 135.750 ;
        RECT 27.405 135.490 27.665 135.750 ;
        RECT 27.725 135.490 27.985 135.750 ;
        RECT 28.045 135.490 28.305 135.750 ;
        RECT 45.275 135.490 45.535 135.750 ;
        RECT 45.595 135.490 45.855 135.750 ;
        RECT 45.915 135.490 46.175 135.750 ;
        RECT 46.235 135.490 46.495 135.750 ;
        RECT 46.555 135.490 46.815 135.750 ;
        RECT 63.785 135.490 64.045 135.750 ;
        RECT 64.105 135.490 64.365 135.750 ;
        RECT 64.425 135.490 64.685 135.750 ;
        RECT 64.745 135.490 65.005 135.750 ;
        RECT 65.065 135.490 65.325 135.750 ;
        RECT 82.295 135.490 82.555 135.750 ;
        RECT 82.615 135.490 82.875 135.750 ;
        RECT 82.935 135.490 83.195 135.750 ;
        RECT 83.255 135.490 83.515 135.750 ;
        RECT 83.575 135.490 83.835 135.750 ;
        RECT 36.020 132.770 36.280 133.030 ;
        RECT 36.340 132.770 36.600 133.030 ;
        RECT 36.660 132.770 36.920 133.030 ;
        RECT 36.980 132.770 37.240 133.030 ;
        RECT 37.300 132.770 37.560 133.030 ;
        RECT 54.530 132.770 54.790 133.030 ;
        RECT 54.850 132.770 55.110 133.030 ;
        RECT 55.170 132.770 55.430 133.030 ;
        RECT 55.490 132.770 55.750 133.030 ;
        RECT 55.810 132.770 56.070 133.030 ;
        RECT 73.040 132.770 73.300 133.030 ;
        RECT 73.360 132.770 73.620 133.030 ;
        RECT 73.680 132.770 73.940 133.030 ;
        RECT 74.000 132.770 74.260 133.030 ;
        RECT 74.320 132.770 74.580 133.030 ;
        RECT 91.550 132.770 91.810 133.030 ;
        RECT 91.870 132.770 92.130 133.030 ;
        RECT 92.190 132.770 92.450 133.030 ;
        RECT 92.510 132.770 92.770 133.030 ;
        RECT 92.830 132.770 93.090 133.030 ;
        RECT 130.300 25.800 130.900 26.400 ;
      LAYER met2 ;
        RECT 19.750 208.180 20.030 210.180 ;
        RECT 26.190 208.180 26.470 210.180 ;
        RECT 32.630 208.180 32.910 210.180 ;
        RECT 39.070 208.180 39.350 210.180 ;
        RECT 45.510 208.180 45.790 210.180 ;
        RECT 51.950 208.180 52.230 210.180 ;
        RECT 58.390 208.180 58.670 210.180 ;
        RECT 64.830 208.180 65.110 210.180 ;
        RECT 71.270 208.180 71.550 210.180 ;
        RECT 77.710 208.180 77.990 210.180 ;
        RECT 84.150 208.180 84.430 210.180 ;
        RECT 90.590 208.180 90.870 210.180 ;
        RECT 19.820 192.390 19.960 208.180 ;
        RECT 26.260 204.970 26.400 208.180 ;
        RECT 26.765 206.155 28.305 206.525 ;
        RECT 32.700 204.970 32.840 208.180 ;
        RECT 39.140 204.970 39.280 208.180 ;
        RECT 45.580 207.430 45.720 208.180 ;
        RECT 45.580 207.290 47.100 207.430 ;
        RECT 40.460 206.690 40.720 207.010 ;
        RECT 26.200 204.650 26.460 204.970 ;
        RECT 32.640 204.650 32.900 204.970 ;
        RECT 39.080 204.650 39.340 204.970 ;
        RECT 40.520 204.630 40.660 206.690 ;
        RECT 45.275 206.155 46.815 206.525 ;
        RECT 46.960 205.990 47.100 207.290 ;
        RECT 45.980 205.670 46.240 205.990 ;
        RECT 46.900 205.670 47.160 205.990 ;
        RECT 47.820 205.670 48.080 205.990 ;
        RECT 45.520 204.650 45.780 204.970 ;
        RECT 40.460 204.310 40.720 204.630 ;
        RECT 26.200 203.970 26.460 204.290 ;
        RECT 28.500 203.970 28.760 204.290 ;
        RECT 26.260 203.270 26.400 203.970 ;
        RECT 26.200 202.950 26.460 203.270 ;
        RECT 26.765 200.715 28.305 201.085 ;
        RECT 28.560 200.550 28.700 203.970 ;
        RECT 36.020 203.435 37.560 203.805 ;
        RECT 28.960 202.610 29.220 202.930 ;
        RECT 29.020 200.550 29.160 202.610 ;
        RECT 32.180 201.930 32.440 202.250 ;
        RECT 31.260 201.250 31.520 201.570 ;
        RECT 28.500 200.230 28.760 200.550 ;
        RECT 28.960 200.230 29.220 200.550 ;
        RECT 26.765 195.275 28.305 195.645 ;
        RECT 19.760 192.070 20.020 192.390 ;
        RECT 28.500 191.730 28.760 192.050 ;
        RECT 26.200 191.050 26.460 191.370 ;
        RECT 26.260 186.950 26.400 191.050 ;
        RECT 26.765 189.835 28.305 190.205 ;
        RECT 28.560 189.670 28.700 191.730 ;
        RECT 28.500 189.350 28.760 189.670 ;
        RECT 26.200 186.630 26.460 186.950 ;
        RECT 26.200 185.950 26.460 186.270 ;
        RECT 26.260 184.230 26.400 185.950 ;
        RECT 28.960 184.930 29.220 185.250 ;
        RECT 26.765 184.395 28.305 184.765 ;
        RECT 26.200 183.910 26.460 184.230 ;
        RECT 29.020 183.210 29.160 184.930 ;
        RECT 28.960 182.890 29.220 183.210 ;
        RECT 29.420 182.890 29.680 183.210 ;
        RECT 26.765 178.955 28.305 179.325 ;
        RECT 22.980 177.450 23.240 177.770 ;
        RECT 23.040 172.330 23.180 177.450 ;
        RECT 25.280 174.050 25.540 174.370 ;
        RECT 22.980 172.010 23.240 172.330 ;
        RECT 23.040 164.750 23.180 172.010 ;
        RECT 25.340 170.630 25.480 174.050 ;
        RECT 26.765 173.515 28.305 173.885 ;
        RECT 28.960 172.010 29.220 172.330 ;
        RECT 25.280 170.310 25.540 170.630 ;
        RECT 29.020 169.270 29.160 172.010 ;
        RECT 29.480 170.290 29.620 182.890 ;
        RECT 31.320 182.870 31.460 201.250 ;
        RECT 32.240 199.530 32.380 201.930 ;
        RECT 34.940 201.590 35.200 201.910 ;
        RECT 35.000 200.550 35.140 201.590 ;
        RECT 34.940 200.230 35.200 200.550 ;
        RECT 32.180 199.210 32.440 199.530 ;
        RECT 32.240 194.090 32.380 199.210 ;
        RECT 36.020 197.995 37.560 198.365 ;
        RECT 32.180 193.770 32.440 194.090 ;
        RECT 32.240 186.270 32.380 193.770 ;
        RECT 34.480 193.430 34.740 193.750 ;
        RECT 34.540 192.050 34.680 193.430 ;
        RECT 39.080 193.090 39.340 193.410 ;
        RECT 36.020 192.555 37.560 192.925 ;
        RECT 34.480 191.730 34.740 192.050 ;
        RECT 33.560 191.390 33.820 191.710 ;
        RECT 34.940 191.390 35.200 191.710 ;
        RECT 33.100 190.710 33.360 191.030 ;
        RECT 33.160 189.670 33.300 190.710 ;
        RECT 33.100 189.350 33.360 189.670 ;
        RECT 33.620 188.650 33.760 191.390 ;
        RECT 34.020 189.010 34.280 189.330 ;
        RECT 33.560 188.330 33.820 188.650 ;
        RECT 32.180 185.950 32.440 186.270 ;
        RECT 33.090 186.095 33.370 186.465 ;
        RECT 33.100 185.950 33.360 186.095 ;
        RECT 31.720 184.930 31.980 185.250 ;
        RECT 31.780 184.230 31.920 184.930 ;
        RECT 32.240 184.230 32.380 185.950 ;
        RECT 31.720 183.910 31.980 184.230 ;
        RECT 32.180 183.910 32.440 184.230 ;
        RECT 31.260 182.550 31.520 182.870 ;
        RECT 29.880 174.730 30.140 175.050 ;
        RECT 29.940 173.350 30.080 174.730 ;
        RECT 29.880 173.030 30.140 173.350 ;
        RECT 29.420 169.970 29.680 170.290 ;
        RECT 28.960 168.950 29.220 169.270 ;
        RECT 26.765 168.075 28.305 168.445 ;
        RECT 22.580 164.610 23.180 164.750 ;
        RECT 22.580 161.790 22.720 164.610 ;
        RECT 29.480 164.510 29.620 169.970 ;
        RECT 29.940 167.570 30.080 173.030 ;
        RECT 31.320 171.990 31.460 182.550 ;
        RECT 33.100 178.130 33.360 178.450 ;
        RECT 32.180 177.110 32.440 177.430 ;
        RECT 31.720 176.770 31.980 177.090 ;
        RECT 31.780 176.070 31.920 176.770 ;
        RECT 32.240 176.070 32.380 177.110 ;
        RECT 33.160 176.070 33.300 178.130 ;
        RECT 31.720 175.750 31.980 176.070 ;
        RECT 32.180 175.750 32.440 176.070 ;
        RECT 33.100 175.750 33.360 176.070 ;
        RECT 33.620 175.390 33.760 188.330 ;
        RECT 34.080 183.550 34.220 189.010 ;
        RECT 34.480 187.990 34.740 188.310 ;
        RECT 34.540 186.270 34.680 187.990 ;
        RECT 35.000 186.950 35.140 191.390 ;
        RECT 39.140 191.370 39.280 193.090 ;
        RECT 40.520 192.350 40.660 204.310 ;
        RECT 44.140 203.970 44.400 204.290 ;
        RECT 44.600 203.970 44.860 204.290 ;
        RECT 43.220 202.270 43.480 202.590 ;
        RECT 43.280 199.530 43.420 202.270 ;
        RECT 43.680 199.890 43.940 200.210 ;
        RECT 43.220 199.210 43.480 199.530 ;
        RECT 43.740 195.110 43.880 199.890 ;
        RECT 44.200 199.530 44.340 203.970 ;
        RECT 44.660 203.270 44.800 203.970 ;
        RECT 44.600 202.950 44.860 203.270 ;
        RECT 45.580 202.590 45.720 204.650 ;
        RECT 45.520 202.270 45.780 202.590 ;
        RECT 46.040 201.570 46.180 205.670 ;
        RECT 46.900 204.650 47.160 204.970 ;
        RECT 47.360 204.650 47.620 204.970 ;
        RECT 46.960 202.250 47.100 204.650 ;
        RECT 46.900 201.930 47.160 202.250 ;
        RECT 44.600 201.250 44.860 201.570 ;
        RECT 45.980 201.250 46.240 201.570 ;
        RECT 46.900 201.250 47.160 201.570 ;
        RECT 44.140 199.210 44.400 199.530 ;
        RECT 44.200 195.110 44.340 199.210 ;
        RECT 44.660 198.850 44.800 201.250 ;
        RECT 45.275 200.715 46.815 201.085 ;
        RECT 46.960 200.550 47.100 201.250 ;
        RECT 46.900 200.230 47.160 200.550 ;
        RECT 47.420 200.210 47.560 204.650 ;
        RECT 47.880 202.930 48.020 205.670 ;
        RECT 52.020 204.970 52.160 208.180 ;
        RECT 58.460 204.970 58.600 208.180 ;
        RECT 64.900 207.430 65.040 208.180 ;
        RECT 64.900 207.290 65.960 207.430 ;
        RECT 63.785 206.155 65.325 206.525 ;
        RECT 65.820 205.650 65.960 207.290 ;
        RECT 71.340 205.650 71.480 208.180 ;
        RECT 76.340 206.690 76.600 207.010 ;
        RECT 72.660 205.670 72.920 205.990 ;
        RECT 65.760 205.330 66.020 205.650 ;
        RECT 71.280 205.330 71.540 205.650 ;
        RECT 51.960 204.650 52.220 204.970 ;
        RECT 57.480 204.650 57.740 204.970 ;
        RECT 58.400 204.650 58.660 204.970 ;
        RECT 66.220 204.650 66.480 204.970 ;
        RECT 53.340 203.970 53.600 204.290 ;
        RECT 52.420 202.950 52.680 203.270 ;
        RECT 47.820 202.610 48.080 202.930 ;
        RECT 47.360 199.890 47.620 200.210 ;
        RECT 44.600 198.530 44.860 198.850 ;
        RECT 43.680 194.790 43.940 195.110 ;
        RECT 44.140 194.790 44.400 195.110 ;
        RECT 44.140 193.090 44.400 193.410 ;
        RECT 40.520 192.210 41.580 192.350 ;
        RECT 39.080 191.050 39.340 191.370 ;
        RECT 37.240 190.710 37.500 191.030 ;
        RECT 35.400 189.010 35.660 189.330 ;
        RECT 35.460 188.650 35.600 189.010 ;
        RECT 35.860 188.670 36.120 188.990 ;
        RECT 35.400 188.330 35.660 188.650 ;
        RECT 35.920 187.880 36.060 188.670 ;
        RECT 37.300 188.650 37.440 190.710 ;
        RECT 37.240 188.330 37.500 188.650 ;
        RECT 39.140 187.970 39.280 191.050 ;
        RECT 40.000 189.010 40.260 189.330 ;
        RECT 39.540 188.330 39.800 188.650 ;
        RECT 35.460 187.740 36.060 187.880 ;
        RECT 34.940 186.630 35.200 186.950 ;
        RECT 35.460 186.610 35.600 187.740 ;
        RECT 38.160 187.650 38.420 187.970 ;
        RECT 38.620 187.650 38.880 187.970 ;
        RECT 39.080 187.650 39.340 187.970 ;
        RECT 36.020 187.115 37.560 187.485 ;
        RECT 35.400 186.290 35.660 186.610 ;
        RECT 38.220 186.520 38.360 187.650 ;
        RECT 34.480 185.950 34.740 186.270 ;
        RECT 35.850 186.095 36.130 186.465 ;
        RECT 37.300 186.380 38.360 186.520 ;
        RECT 38.680 186.465 38.820 187.650 ;
        RECT 35.860 185.950 36.120 186.095 ;
        RECT 34.540 183.890 34.680 185.950 ;
        RECT 36.780 185.270 37.040 185.590 ;
        RECT 35.400 184.930 35.660 185.250 ;
        RECT 34.480 183.570 34.740 183.890 ;
        RECT 34.020 183.230 34.280 183.550 ;
        RECT 34.080 178.110 34.220 183.230 ;
        RECT 34.020 177.790 34.280 178.110 ;
        RECT 33.560 175.070 33.820 175.390 ;
        RECT 31.260 171.670 31.520 171.990 ;
        RECT 32.640 171.330 32.900 171.650 ;
        RECT 32.700 170.630 32.840 171.330 ;
        RECT 32.640 170.310 32.900 170.630 ;
        RECT 32.180 168.950 32.440 169.270 ;
        RECT 29.880 167.250 30.140 167.570 ;
        RECT 29.880 165.890 30.140 166.210 ;
        RECT 29.940 164.850 30.080 165.890 ;
        RECT 29.880 164.530 30.140 164.850 ;
        RECT 29.420 164.190 29.680 164.510 ;
        RECT 29.420 163.170 29.680 163.490 ;
        RECT 26.765 162.635 28.305 163.005 ;
        RECT 29.480 162.470 29.620 163.170 ;
        RECT 29.420 162.150 29.680 162.470 ;
        RECT 22.520 161.470 22.780 161.790 ;
        RECT 29.940 160.770 30.080 164.530 ;
        RECT 29.880 160.450 30.140 160.770 ;
        RECT 26.765 157.195 28.305 157.565 ;
        RECT 32.240 156.350 32.380 168.950 ;
        RECT 33.620 165.190 33.760 175.070 ;
        RECT 34.080 174.710 34.220 177.790 ;
        RECT 34.540 177.090 34.680 183.570 ;
        RECT 35.460 181.510 35.600 184.930 ;
        RECT 36.840 183.890 36.980 185.270 ;
        RECT 36.780 183.570 37.040 183.890 ;
        RECT 37.300 182.950 37.440 186.380 ;
        RECT 38.610 186.095 38.890 186.465 ;
        RECT 38.160 185.785 38.420 185.930 ;
        RECT 37.700 185.270 37.960 185.590 ;
        RECT 38.150 185.415 38.430 185.785 ;
        RECT 38.620 185.610 38.880 185.930 ;
        RECT 37.760 184.230 37.900 185.270 ;
        RECT 37.700 183.910 37.960 184.230 ;
        RECT 38.680 183.550 38.820 185.610 ;
        RECT 38.620 183.230 38.880 183.550 ;
        RECT 37.300 182.810 38.360 182.950 ;
        RECT 36.020 181.675 37.560 182.045 ;
        RECT 35.400 181.190 35.660 181.510 ;
        RECT 37.700 178.470 37.960 178.790 ;
        RECT 35.400 177.110 35.660 177.430 ;
        RECT 34.480 176.770 34.740 177.090 ;
        RECT 34.540 175.050 34.680 176.770 ;
        RECT 35.460 175.390 35.600 177.110 ;
        RECT 36.020 176.235 37.560 176.605 ;
        RECT 37.760 175.390 37.900 178.470 ;
        RECT 38.220 177.770 38.360 182.810 ;
        RECT 39.140 181.170 39.280 187.650 ;
        RECT 39.080 180.850 39.340 181.170 ;
        RECT 38.620 180.170 38.880 180.490 ;
        RECT 38.680 178.450 38.820 180.170 ;
        RECT 38.620 178.130 38.880 178.450 ;
        RECT 38.160 177.450 38.420 177.770 ;
        RECT 39.600 177.430 39.740 188.330 ;
        RECT 40.060 186.440 40.200 189.010 ;
        RECT 40.000 186.120 40.260 186.440 ;
        RECT 40.460 185.785 40.720 185.930 ;
        RECT 40.450 185.415 40.730 185.785 ;
        RECT 40.460 182.890 40.720 183.210 ;
        RECT 40.000 177.790 40.260 178.110 ;
        RECT 39.540 177.110 39.800 177.430 ;
        RECT 38.620 176.770 38.880 177.090 ;
        RECT 38.680 176.070 38.820 176.770 ;
        RECT 40.060 176.070 40.200 177.790 ;
        RECT 38.620 175.750 38.880 176.070 ;
        RECT 40.000 175.750 40.260 176.070 ;
        RECT 35.400 175.070 35.660 175.390 ;
        RECT 37.700 175.070 37.960 175.390 ;
        RECT 34.480 174.730 34.740 175.050 ;
        RECT 34.020 174.390 34.280 174.710 ;
        RECT 35.460 172.920 35.600 175.070 ;
        RECT 35.860 172.920 36.120 173.010 ;
        RECT 35.460 172.780 36.120 172.920 ;
        RECT 35.860 172.690 36.120 172.780 ;
        RECT 37.760 172.670 37.900 175.070 ;
        RECT 37.700 172.350 37.960 172.670 ;
        RECT 34.020 171.670 34.280 171.990 ;
        RECT 34.480 171.670 34.740 171.990 ;
        RECT 33.560 164.870 33.820 165.190 ;
        RECT 33.620 161.450 33.760 164.870 ;
        RECT 33.560 161.130 33.820 161.450 ;
        RECT 33.620 159.070 33.760 161.130 ;
        RECT 34.080 159.410 34.220 171.670 ;
        RECT 34.540 164.510 34.680 171.670 ;
        RECT 36.020 170.795 37.560 171.165 ;
        RECT 35.860 169.290 36.120 169.610 ;
        RECT 35.920 167.230 36.060 169.290 ;
        RECT 37.760 167.910 37.900 172.350 ;
        RECT 38.160 172.010 38.420 172.330 ;
        RECT 39.540 172.010 39.800 172.330 ;
        RECT 38.220 168.930 38.360 172.010 ;
        RECT 39.080 171.330 39.340 171.650 ;
        RECT 39.140 169.950 39.280 171.330 ;
        RECT 39.080 169.630 39.340 169.950 ;
        RECT 38.620 169.290 38.880 169.610 ;
        RECT 38.160 168.610 38.420 168.930 ;
        RECT 37.700 167.590 37.960 167.910 ;
        RECT 35.860 166.910 36.120 167.230 ;
        RECT 38.680 166.890 38.820 169.290 ;
        RECT 39.140 166.890 39.280 169.630 ;
        RECT 39.600 167.910 39.740 172.010 ;
        RECT 40.000 171.330 40.260 171.650 ;
        RECT 40.060 169.610 40.200 171.330 ;
        RECT 40.520 170.290 40.660 182.890 ;
        RECT 40.920 180.510 41.180 180.830 ;
        RECT 40.980 179.810 41.120 180.510 ;
        RECT 40.920 179.490 41.180 179.810 ;
        RECT 40.920 177.790 41.180 178.110 ;
        RECT 40.980 174.370 41.120 177.790 ;
        RECT 40.920 174.050 41.180 174.370 ;
        RECT 41.440 172.330 41.580 192.210 ;
        RECT 44.200 192.050 44.340 193.090 ;
        RECT 44.140 191.730 44.400 192.050 ;
        RECT 43.680 191.050 43.940 191.370 ;
        RECT 44.660 191.110 44.800 198.530 ;
        RECT 47.880 197.150 48.020 202.610 ;
        RECT 48.280 201.250 48.540 201.570 ;
        RECT 50.120 201.250 50.380 201.570 ;
        RECT 48.340 200.210 48.480 201.250 ;
        RECT 48.280 199.890 48.540 200.210 ;
        RECT 50.180 199.870 50.320 201.250 ;
        RECT 50.120 199.550 50.380 199.870 ;
        RECT 47.820 196.830 48.080 197.150 ;
        RECT 47.820 195.810 48.080 196.130 ;
        RECT 45.275 195.275 46.815 195.645 ;
        RECT 45.060 193.090 45.320 193.410 ;
        RECT 45.120 191.710 45.260 193.090 ;
        RECT 45.060 191.390 45.320 191.710 ;
        RECT 46.900 191.390 47.160 191.710 ;
        RECT 43.220 190.370 43.480 190.690 ;
        RECT 42.760 187.990 43.020 188.310 ;
        RECT 41.840 186.630 42.100 186.950 ;
        RECT 41.900 186.465 42.040 186.630 ;
        RECT 41.830 186.095 42.110 186.465 ;
        RECT 42.300 184.930 42.560 185.250 ;
        RECT 41.840 183.570 42.100 183.890 ;
        RECT 41.900 181.510 42.040 183.570 ;
        RECT 42.360 183.210 42.500 184.930 ;
        RECT 42.820 183.890 42.960 187.990 ;
        RECT 43.280 186.270 43.420 190.370 ;
        RECT 43.740 189.670 43.880 191.050 ;
        RECT 44.200 190.970 44.800 191.110 ;
        RECT 43.680 189.350 43.940 189.670 ;
        RECT 44.200 189.330 44.340 190.970 ;
        RECT 45.275 189.835 46.815 190.205 ;
        RECT 46.960 189.670 47.100 191.390 ;
        RECT 46.900 189.350 47.160 189.670 ;
        RECT 44.140 189.010 44.400 189.330 ;
        RECT 47.360 187.650 47.620 187.970 ;
        RECT 47.420 186.610 47.560 187.650 ;
        RECT 47.360 186.290 47.620 186.610 ;
        RECT 43.220 185.950 43.480 186.270 ;
        RECT 44.140 185.610 44.400 185.930 ;
        RECT 44.200 184.230 44.340 185.610 ;
        RECT 44.600 184.930 44.860 185.250 ;
        RECT 44.140 183.910 44.400 184.230 ;
        RECT 44.660 183.890 44.800 184.930 ;
        RECT 45.275 184.395 46.815 184.765 ;
        RECT 42.760 183.570 43.020 183.890 ;
        RECT 44.600 183.570 44.860 183.890 ;
        RECT 47.880 183.630 48.020 195.810 ;
        RECT 51.960 192.070 52.220 192.390 ;
        RECT 51.500 190.370 51.760 190.690 ;
        RECT 51.560 188.650 51.700 190.370 ;
        RECT 48.280 188.330 48.540 188.650 ;
        RECT 51.500 188.330 51.760 188.650 ;
        RECT 48.340 184.230 48.480 188.330 ;
        RECT 50.120 184.930 50.380 185.250 ;
        RECT 48.280 183.910 48.540 184.230 ;
        RECT 44.660 183.210 44.800 183.570 ;
        RECT 47.420 183.550 48.020 183.630 ;
        RECT 47.360 183.490 48.020 183.550 ;
        RECT 47.360 183.230 47.620 183.490 ;
        RECT 42.300 182.890 42.560 183.210 ;
        RECT 44.600 182.890 44.860 183.210 ;
        RECT 42.760 182.550 43.020 182.870 ;
        RECT 42.300 182.210 42.560 182.530 ;
        RECT 42.360 181.510 42.500 182.210 ;
        RECT 41.840 181.190 42.100 181.510 ;
        RECT 42.300 181.190 42.560 181.510 ;
        RECT 42.820 180.830 42.960 182.550 ;
        RECT 42.760 180.510 43.020 180.830 ;
        RECT 41.840 179.490 42.100 179.810 ;
        RECT 43.680 179.490 43.940 179.810 ;
        RECT 41.900 177.770 42.040 179.490 ;
        RECT 43.740 177.770 43.880 179.490 ;
        RECT 45.275 178.955 46.815 179.325 ;
        RECT 41.840 177.450 42.100 177.770 ;
        RECT 43.680 177.450 43.940 177.770 ;
        RECT 41.900 173.350 42.040 177.450 ;
        RECT 43.220 176.770 43.480 177.090 ;
        RECT 43.280 175.730 43.420 176.770 ;
        RECT 43.220 175.410 43.480 175.730 ;
        RECT 41.840 173.030 42.100 173.350 ;
        RECT 41.380 172.010 41.640 172.330 ;
        RECT 40.460 169.970 40.720 170.290 ;
        RECT 40.000 169.290 40.260 169.610 ;
        RECT 39.540 167.590 39.800 167.910 ;
        RECT 38.620 166.570 38.880 166.890 ;
        RECT 39.080 166.570 39.340 166.890 ;
        RECT 34.940 165.890 35.200 166.210 ;
        RECT 38.160 165.890 38.420 166.210 ;
        RECT 35.000 164.510 35.140 165.890 ;
        RECT 36.020 165.355 37.560 165.725 ;
        RECT 34.480 164.190 34.740 164.510 ;
        RECT 34.940 164.190 35.200 164.510 ;
        RECT 34.540 161.190 34.680 164.190 ;
        RECT 38.220 164.170 38.360 165.890 ;
        RECT 39.140 164.850 39.280 166.570 ;
        RECT 40.060 166.210 40.200 169.290 ;
        RECT 42.300 166.230 42.560 166.550 ;
        RECT 40.000 165.890 40.260 166.210 ;
        RECT 42.360 165.190 42.500 166.230 ;
        RECT 42.300 164.870 42.560 165.190 ;
        RECT 39.080 164.530 39.340 164.850 ;
        RECT 38.160 163.850 38.420 164.170 ;
        RECT 36.320 163.170 36.580 163.490 ;
        RECT 37.700 163.170 37.960 163.490 ;
        RECT 36.380 162.470 36.520 163.170 ;
        RECT 36.320 162.150 36.580 162.470 ;
        RECT 37.760 161.450 37.900 163.170 ;
        RECT 38.220 162.470 38.360 163.850 ;
        RECT 38.160 162.150 38.420 162.470 ;
        RECT 38.220 161.450 38.360 162.150 ;
        RECT 39.140 161.450 39.280 164.530 ;
        RECT 43.280 162.130 43.420 175.410 ;
        RECT 43.740 173.010 43.880 177.450 ;
        RECT 46.900 176.770 47.160 177.090 ;
        RECT 46.960 175.730 47.100 176.770 ;
        RECT 46.900 175.410 47.160 175.730 ;
        RECT 47.420 175.585 47.560 183.230 ;
        RECT 50.180 183.210 50.320 184.930 ;
        RECT 48.740 182.890 49.000 183.210 ;
        RECT 50.120 182.890 50.380 183.210 ;
        RECT 48.800 181.510 48.940 182.890 ;
        RECT 49.660 182.550 49.920 182.870 ;
        RECT 48.740 181.190 49.000 181.510 ;
        RECT 49.720 180.150 49.860 182.550 ;
        RECT 49.660 179.830 49.920 180.150 ;
        RECT 47.820 177.450 48.080 177.770 ;
        RECT 49.720 177.680 49.860 179.830 ;
        RECT 51.040 177.680 51.300 177.770 ;
        RECT 49.720 177.540 51.300 177.680 ;
        RECT 51.040 177.450 51.300 177.540 ;
        RECT 47.350 175.215 47.630 175.585 ;
        RECT 44.600 174.730 44.860 175.050 ;
        RECT 44.140 174.390 44.400 174.710 ;
        RECT 43.680 172.690 43.940 173.010 ;
        RECT 43.680 171.330 43.940 171.650 ;
        RECT 43.740 170.290 43.880 171.330 ;
        RECT 43.680 169.970 43.940 170.290 ;
        RECT 44.200 163.490 44.340 174.390 ;
        RECT 44.660 169.270 44.800 174.730 ;
        RECT 45.275 173.515 46.815 173.885 ;
        RECT 47.420 172.670 47.560 175.215 ;
        RECT 47.880 173.350 48.020 177.450 ;
        RECT 51.500 177.110 51.760 177.430 ;
        RECT 48.280 176.770 48.540 177.090 ;
        RECT 47.820 173.030 48.080 173.350 ;
        RECT 47.360 172.350 47.620 172.670 ;
        RECT 48.340 172.330 48.480 176.770 ;
        RECT 51.560 176.070 51.700 177.110 ;
        RECT 51.500 175.750 51.760 176.070 ;
        RECT 52.020 175.730 52.160 192.070 ;
        RECT 52.480 190.690 52.620 202.950 ;
        RECT 53.400 202.590 53.540 203.970 ;
        RECT 54.530 203.435 56.070 203.805 ;
        RECT 57.540 203.270 57.680 204.650 ;
        RECT 57.940 204.310 58.200 204.630 ;
        RECT 57.480 202.950 57.740 203.270 ;
        RECT 53.340 202.270 53.600 202.590 ;
        RECT 57.020 202.270 57.280 202.590 ;
        RECT 53.400 198.850 53.540 202.270 ;
        RECT 57.080 200.550 57.220 202.270 ;
        RECT 57.020 200.230 57.280 200.550 ;
        RECT 53.340 198.530 53.600 198.850 ;
        RECT 54.530 197.995 56.070 198.365 ;
        RECT 58.000 196.810 58.140 204.310 ;
        RECT 60.240 203.970 60.500 204.290 ;
        RECT 60.700 203.970 60.960 204.290 ;
        RECT 63.000 203.970 63.260 204.290 ;
        RECT 58.400 200.230 58.660 200.550 ;
        RECT 57.940 196.490 58.200 196.810 ;
        RECT 58.460 196.550 58.600 200.230 ;
        RECT 60.300 199.870 60.440 203.970 ;
        RECT 60.240 199.550 60.500 199.870 ;
        RECT 58.860 199.210 59.120 199.530 ;
        RECT 58.920 197.150 59.060 199.210 ;
        RECT 58.860 196.830 59.120 197.150 ;
        RECT 59.780 196.830 60.040 197.150 ;
        RECT 53.800 195.810 54.060 196.130 ;
        RECT 53.860 194.090 54.000 195.810 ;
        RECT 53.800 193.770 54.060 194.090 ;
        RECT 53.340 193.090 53.600 193.410 ;
        RECT 53.400 191.710 53.540 193.090 ;
        RECT 54.530 192.555 56.070 192.925 ;
        RECT 52.880 191.390 53.140 191.710 ;
        RECT 53.340 191.390 53.600 191.710 ;
        RECT 52.420 190.370 52.680 190.690 ;
        RECT 52.480 188.650 52.620 190.370 ;
        RECT 52.940 189.670 53.080 191.390 ;
        RECT 58.000 191.370 58.140 196.490 ;
        RECT 58.460 196.410 59.060 196.550 ;
        RECT 58.920 196.130 59.060 196.410 ;
        RECT 58.400 195.810 58.660 196.130 ;
        RECT 58.860 195.810 59.120 196.130 ;
        RECT 57.940 191.050 58.200 191.370 ;
        RECT 53.800 190.710 54.060 191.030 ;
        RECT 56.100 190.710 56.360 191.030 ;
        RECT 52.880 189.350 53.140 189.670 ;
        RECT 53.860 188.650 54.000 190.710 ;
        RECT 56.160 188.650 56.300 190.710 ;
        RECT 56.560 190.370 56.820 190.690 ;
        RECT 56.620 188.650 56.760 190.370 ;
        RECT 52.420 188.330 52.680 188.650 ;
        RECT 53.800 188.330 54.060 188.650 ;
        RECT 56.100 188.330 56.360 188.650 ;
        RECT 56.560 188.330 56.820 188.650 ;
        RECT 57.020 187.990 57.280 188.310 ;
        RECT 54.530 187.115 56.070 187.485 ;
        RECT 57.080 186.270 57.220 187.990 ;
        RECT 57.020 185.950 57.280 186.270 ;
        RECT 57.080 184.230 57.220 185.950 ;
        RECT 57.020 183.910 57.280 184.230 ;
        RECT 52.880 182.890 53.140 183.210 ;
        RECT 57.480 182.890 57.740 183.210 ;
        RECT 52.940 177.770 53.080 182.890 ;
        RECT 56.560 182.210 56.820 182.530 ;
        RECT 54.530 181.675 56.070 182.045 ;
        RECT 56.620 178.790 56.760 182.210 ;
        RECT 55.180 178.470 55.440 178.790 ;
        RECT 56.560 178.470 56.820 178.790 ;
        RECT 55.240 177.770 55.380 178.470 ;
        RECT 52.880 177.450 53.140 177.770 ;
        RECT 53.340 177.450 53.600 177.770 ;
        RECT 55.180 177.510 55.440 177.770 ;
        RECT 53.860 177.450 55.440 177.510 ;
        RECT 51.960 175.410 52.220 175.730 ;
        RECT 48.280 172.010 48.540 172.330 ;
        RECT 52.420 172.010 52.680 172.330 ;
        RECT 52.480 169.950 52.620 172.010 ;
        RECT 52.420 169.630 52.680 169.950 ;
        RECT 44.600 168.950 44.860 169.270 ;
        RECT 44.660 166.890 44.800 168.950 ;
        RECT 45.275 168.075 46.815 168.445 ;
        RECT 47.360 167.250 47.620 167.570 ;
        RECT 52.940 167.310 53.080 177.450 ;
        RECT 53.400 177.090 53.540 177.450 ;
        RECT 53.860 177.430 55.380 177.450 ;
        RECT 53.800 177.370 55.380 177.430 ;
        RECT 53.800 177.110 54.060 177.370 ;
        RECT 53.340 176.770 53.600 177.090 ;
        RECT 53.400 174.370 53.540 176.770 ;
        RECT 54.530 176.235 56.070 176.605 ;
        RECT 57.540 176.070 57.680 182.890 ;
        RECT 57.480 175.750 57.740 176.070 ;
        RECT 53.340 174.050 53.600 174.370 ;
        RECT 56.560 171.330 56.820 171.650 ;
        RECT 54.530 170.795 56.070 171.165 ;
        RECT 53.800 169.630 54.060 169.950 ;
        RECT 53.860 167.910 54.000 169.630 ;
        RECT 53.800 167.590 54.060 167.910 ;
        RECT 44.600 166.570 44.860 166.890 ;
        RECT 47.420 164.510 47.560 167.250 ;
        RECT 52.940 167.170 54.000 167.310 ;
        RECT 52.880 166.230 53.140 166.550 ;
        RECT 44.600 164.190 44.860 164.510 ;
        RECT 47.360 164.190 47.620 164.510 ;
        RECT 48.740 164.190 49.000 164.510 ;
        RECT 44.140 163.170 44.400 163.490 ;
        RECT 43.220 161.810 43.480 162.130 ;
        RECT 44.660 161.870 44.800 164.190 ;
        RECT 46.900 163.170 47.160 163.490 ;
        RECT 45.275 162.635 46.815 163.005 ;
        RECT 44.660 161.730 45.720 161.870 ;
        RECT 45.580 161.450 45.720 161.730 ;
        RECT 46.960 161.450 47.100 163.170 ;
        RECT 47.420 162.130 47.560 164.190 ;
        RECT 48.800 162.130 48.940 164.190 ;
        RECT 49.200 163.510 49.460 163.830 ;
        RECT 49.260 162.470 49.400 163.510 ;
        RECT 49.200 162.150 49.460 162.470 ;
        RECT 47.360 161.810 47.620 162.130 ;
        RECT 48.740 161.810 49.000 162.130 ;
        RECT 34.540 161.050 35.600 161.190 ;
        RECT 37.700 161.130 37.960 161.450 ;
        RECT 38.160 161.130 38.420 161.450 ;
        RECT 39.080 161.130 39.340 161.450 ;
        RECT 45.520 161.130 45.780 161.450 ;
        RECT 45.980 161.130 46.240 161.450 ;
        RECT 46.900 161.130 47.160 161.450 ;
        RECT 52.420 161.130 52.680 161.450 ;
        RECT 34.940 160.450 35.200 160.770 ;
        RECT 35.000 159.750 35.140 160.450 ;
        RECT 35.460 159.750 35.600 161.050 ;
        RECT 36.020 159.915 37.560 160.285 ;
        RECT 34.940 159.430 35.200 159.750 ;
        RECT 35.400 159.430 35.660 159.750 ;
        RECT 34.020 159.090 34.280 159.410 ;
        RECT 39.140 159.070 39.280 161.130 ;
        RECT 44.140 160.450 44.400 160.770 ;
        RECT 44.200 159.070 44.340 160.450 ;
        RECT 45.580 159.750 45.720 161.130 ;
        RECT 45.520 159.430 45.780 159.750 ;
        RECT 33.560 158.750 33.820 159.070 ;
        RECT 39.080 158.750 39.340 159.070 ;
        RECT 44.140 158.750 44.400 159.070 ;
        RECT 45.520 158.750 45.780 159.070 ;
        RECT 34.020 157.730 34.280 158.050 ;
        RECT 32.180 156.030 32.440 156.350 ;
        RECT 34.080 155.670 34.220 157.730 ;
        RECT 39.140 157.030 39.280 158.750 ;
        RECT 41.840 157.730 42.100 158.050 ;
        RECT 45.580 157.850 45.720 158.750 ;
        RECT 46.040 158.730 46.180 161.130 ;
        RECT 49.200 160.790 49.460 161.110 ;
        RECT 48.740 160.450 49.000 160.770 ;
        RECT 48.280 159.430 48.540 159.750 ;
        RECT 48.340 159.150 48.480 159.430 ;
        RECT 47.420 159.070 48.480 159.150 ;
        RECT 48.800 159.070 48.940 160.450 ;
        RECT 47.360 159.010 48.480 159.070 ;
        RECT 47.360 158.750 47.620 159.010 ;
        RECT 48.740 158.750 49.000 159.070 ;
        RECT 49.260 158.730 49.400 160.790 ;
        RECT 49.660 160.450 49.920 160.770 ;
        RECT 49.720 159.750 49.860 160.450 ;
        RECT 52.480 159.750 52.620 161.130 ;
        RECT 49.660 159.430 49.920 159.750 ;
        RECT 52.420 159.430 52.680 159.750 ;
        RECT 52.940 159.070 53.080 166.230 ;
        RECT 53.340 165.890 53.600 166.210 ;
        RECT 53.400 165.190 53.540 165.890 ;
        RECT 53.860 165.190 54.000 167.170 ;
        RECT 56.620 166.890 56.760 171.330 ;
        RECT 54.260 166.630 54.520 166.890 ;
        RECT 54.710 166.630 54.990 166.745 ;
        RECT 54.260 166.570 54.990 166.630 ;
        RECT 56.560 166.570 56.820 166.890 ;
        RECT 54.320 166.490 54.990 166.570 ;
        RECT 54.710 166.375 54.990 166.490 ;
        RECT 54.530 165.355 56.070 165.725 ;
        RECT 53.340 164.870 53.600 165.190 ;
        RECT 53.800 164.870 54.060 165.190 ;
        RECT 54.720 161.470 54.980 161.790 ;
        RECT 54.780 160.770 54.920 161.470 ;
        RECT 54.720 160.450 54.980 160.770 ;
        RECT 54.530 159.915 56.070 160.285 ;
        RECT 57.540 159.410 57.680 175.750 ;
        RECT 57.940 171.330 58.200 171.650 ;
        RECT 58.000 164.510 58.140 171.330 ;
        RECT 58.460 169.950 58.600 195.810 ;
        RECT 59.320 193.090 59.580 193.410 ;
        RECT 59.380 190.690 59.520 193.090 ;
        RECT 59.840 191.710 59.980 196.830 ;
        RECT 60.760 196.470 60.900 203.970 ;
        RECT 62.540 202.950 62.800 203.270 ;
        RECT 60.700 196.150 60.960 196.470 ;
        RECT 62.080 194.450 62.340 194.770 ;
        RECT 60.700 193.090 60.960 193.410 ;
        RECT 59.780 191.390 60.040 191.710 ;
        RECT 59.320 190.370 59.580 190.690 ;
        RECT 60.760 189.670 60.900 193.090 ;
        RECT 60.700 189.350 60.960 189.670 ;
        RECT 58.860 188.330 59.120 188.650 ;
        RECT 58.920 186.950 59.060 188.330 ;
        RECT 58.860 186.630 59.120 186.950 ;
        RECT 60.240 185.950 60.500 186.270 ;
        RECT 59.780 183.230 60.040 183.550 ;
        RECT 59.320 178.130 59.580 178.450 ;
        RECT 59.380 172.330 59.520 178.130 ;
        RECT 59.840 172.330 59.980 183.230 ;
        RECT 60.300 172.330 60.440 185.950 ;
        RECT 60.760 185.930 60.900 189.350 ;
        RECT 61.160 187.650 61.420 187.970 ;
        RECT 60.700 185.610 60.960 185.930 ;
        RECT 61.220 181.510 61.360 187.650 ;
        RECT 62.140 185.670 62.280 194.450 ;
        RECT 62.600 191.030 62.740 202.950 ;
        RECT 63.060 199.870 63.200 203.970 ;
        RECT 66.280 203.270 66.420 204.650 ;
        RECT 67.600 203.970 67.860 204.290 ;
        RECT 72.200 203.970 72.460 204.290 ;
        RECT 66.220 202.950 66.480 203.270 ;
        RECT 66.680 202.270 66.940 202.590 ;
        RECT 67.140 202.270 67.400 202.590 ;
        RECT 63.785 200.715 65.325 201.085 ;
        RECT 66.740 200.550 66.880 202.270 ;
        RECT 66.680 200.230 66.940 200.550 ;
        RECT 63.000 199.550 63.260 199.870 ;
        RECT 65.300 199.210 65.560 199.530 ;
        RECT 65.360 197.150 65.500 199.210 ;
        RECT 65.300 196.830 65.560 197.150 ;
        RECT 66.220 196.490 66.480 196.810 ;
        RECT 63.000 195.810 63.260 196.130 ;
        RECT 65.760 195.810 66.020 196.130 ;
        RECT 63.060 191.710 63.200 195.810 ;
        RECT 63.785 195.275 65.325 195.645 ;
        RECT 65.820 193.750 65.960 195.810 ;
        RECT 65.760 193.430 66.020 193.750 ;
        RECT 66.280 192.390 66.420 196.490 ;
        RECT 67.200 194.430 67.340 202.270 ;
        RECT 67.660 199.530 67.800 203.970 ;
        RECT 72.260 199.870 72.400 203.970 ;
        RECT 72.200 199.550 72.460 199.870 ;
        RECT 67.600 199.210 67.860 199.530 ;
        RECT 67.140 194.110 67.400 194.430 ;
        RECT 66.220 192.070 66.480 192.390 ;
        RECT 63.000 191.390 63.260 191.710 ;
        RECT 66.680 191.390 66.940 191.710 ;
        RECT 62.540 190.710 62.800 191.030 ;
        RECT 62.600 188.990 62.740 190.710 ;
        RECT 63.000 190.370 63.260 190.690 ;
        RECT 63.060 189.070 63.200 190.370 ;
        RECT 63.785 189.835 65.325 190.205 ;
        RECT 63.060 188.990 63.660 189.070 ;
        RECT 62.540 188.670 62.800 188.990 ;
        RECT 63.060 188.930 63.720 188.990 ;
        RECT 63.460 188.670 63.720 188.930 ;
        RECT 62.600 186.270 62.740 188.670 ;
        RECT 63.920 188.330 64.180 188.650 ;
        RECT 63.460 188.220 63.720 188.310 ;
        RECT 63.060 188.080 63.720 188.220 ;
        RECT 62.540 185.950 62.800 186.270 ;
        RECT 62.140 185.530 62.740 185.670 ;
        RECT 62.080 184.930 62.340 185.250 ;
        RECT 62.140 181.510 62.280 184.930 ;
        RECT 61.160 181.190 61.420 181.510 ;
        RECT 62.080 181.190 62.340 181.510 ;
        RECT 61.160 179.490 61.420 179.810 ;
        RECT 62.080 179.490 62.340 179.810 ;
        RECT 60.700 178.470 60.960 178.790 ;
        RECT 59.320 172.010 59.580 172.330 ;
        RECT 59.780 172.010 60.040 172.330 ;
        RECT 60.240 172.010 60.500 172.330 ;
        RECT 58.400 169.630 58.660 169.950 ;
        RECT 57.940 164.190 58.200 164.510 ;
        RECT 58.000 161.450 58.140 164.190 ;
        RECT 59.840 163.830 59.980 172.010 ;
        RECT 60.760 171.650 60.900 178.470 ;
        RECT 61.220 178.110 61.360 179.490 ;
        RECT 61.160 177.790 61.420 178.110 ;
        RECT 61.620 176.770 61.880 177.090 ;
        RECT 61.680 176.070 61.820 176.770 ;
        RECT 62.140 176.070 62.280 179.490 ;
        RECT 61.620 175.750 61.880 176.070 ;
        RECT 62.080 175.750 62.340 176.070 ;
        RECT 62.070 175.215 62.350 175.585 ;
        RECT 61.160 174.050 61.420 174.370 ;
        RECT 61.220 172.330 61.360 174.050 ;
        RECT 61.620 172.350 61.880 172.670 ;
        RECT 61.160 172.010 61.420 172.330 ;
        RECT 60.700 171.330 60.960 171.650 ;
        RECT 60.700 169.630 60.960 169.950 ;
        RECT 59.780 163.510 60.040 163.830 ;
        RECT 59.840 161.985 59.980 163.510 ;
        RECT 59.770 161.615 60.050 161.985 ;
        RECT 60.760 161.450 60.900 169.630 ;
        RECT 57.940 161.130 58.200 161.450 ;
        RECT 60.700 161.130 60.960 161.450 ;
        RECT 60.700 160.450 60.960 160.770 ;
        RECT 61.160 160.450 61.420 160.770 ;
        RECT 57.480 159.090 57.740 159.410 ;
        RECT 60.760 159.070 60.900 160.450 ;
        RECT 52.880 158.750 53.140 159.070 ;
        RECT 60.700 158.750 60.960 159.070 ;
        RECT 45.980 158.410 46.240 158.730 ;
        RECT 49.200 158.410 49.460 158.730 ;
        RECT 49.260 158.050 49.400 158.410 ;
        RECT 39.080 156.710 39.340 157.030 ;
        RECT 41.900 156.010 42.040 157.730 ;
        RECT 45.580 157.710 47.100 157.850 ;
        RECT 49.200 157.730 49.460 158.050 ;
        RECT 54.260 157.850 54.520 158.050 ;
        RECT 61.220 157.850 61.360 160.450 ;
        RECT 61.680 159.750 61.820 172.350 ;
        RECT 62.140 168.930 62.280 175.215 ;
        RECT 62.080 168.610 62.340 168.930 ;
        RECT 62.600 166.890 62.740 185.530 ;
        RECT 63.060 177.770 63.200 188.080 ;
        RECT 63.460 187.990 63.720 188.080 ;
        RECT 63.980 186.610 64.120 188.330 ;
        RECT 65.300 187.650 65.560 187.970 ;
        RECT 63.920 186.290 64.180 186.610 ;
        RECT 65.360 186.270 65.500 187.650 ;
        RECT 65.300 185.950 65.560 186.270 ;
        RECT 65.760 185.950 66.020 186.270 ;
        RECT 63.785 184.395 65.325 184.765 ;
        RECT 65.820 183.890 65.960 185.950 ;
        RECT 65.760 183.570 66.020 183.890 ;
        RECT 66.740 183.630 66.880 191.390 ;
        RECT 67.200 184.230 67.340 194.110 ;
        RECT 67.140 183.910 67.400 184.230 ;
        RECT 66.740 183.490 67.340 183.630 ;
        RECT 63.785 178.955 65.325 179.325 ;
        RECT 63.000 177.450 63.260 177.770 ;
        RECT 63.060 171.990 63.200 177.450 ;
        RECT 65.760 175.750 66.020 176.070 ;
        RECT 63.450 175.470 63.730 175.585 ;
        RECT 63.450 175.390 64.120 175.470 ;
        RECT 63.450 175.330 64.180 175.390 ;
        RECT 63.450 175.215 63.730 175.330 ;
        RECT 63.920 175.070 64.180 175.330 ;
        RECT 65.300 175.070 65.560 175.390 ;
        RECT 65.360 174.710 65.500 175.070 ;
        RECT 65.300 174.390 65.560 174.710 ;
        RECT 63.785 173.515 65.325 173.885 ;
        RECT 63.000 171.670 63.260 171.990 ;
        RECT 63.060 170.630 63.200 171.670 ;
        RECT 63.000 170.310 63.260 170.630 ;
        RECT 63.785 168.075 65.325 168.445 ;
        RECT 62.540 166.570 62.800 166.890 ;
        RECT 63.000 165.890 63.260 166.210 ;
        RECT 63.060 165.190 63.200 165.890 ;
        RECT 63.000 164.870 63.260 165.190 ;
        RECT 63.785 162.635 65.325 163.005 ;
        RECT 65.820 162.470 65.960 175.750 ;
        RECT 66.680 175.410 66.940 175.730 ;
        RECT 66.220 174.050 66.480 174.370 ;
        RECT 66.280 172.330 66.420 174.050 ;
        RECT 66.220 172.010 66.480 172.330 ;
        RECT 66.740 170.630 66.880 175.410 ;
        RECT 66.680 170.310 66.940 170.630 ;
        RECT 66.680 168.610 66.940 168.930 ;
        RECT 66.740 167.570 66.880 168.610 ;
        RECT 66.220 167.250 66.480 167.570 ;
        RECT 66.680 167.250 66.940 167.570 ;
        RECT 65.760 162.150 66.020 162.470 ;
        RECT 64.380 161.870 64.640 162.130 ;
        RECT 63.980 161.810 64.640 161.870 ;
        RECT 63.980 161.730 64.580 161.810 ;
        RECT 63.980 161.450 64.120 161.730 ;
        RECT 65.750 161.615 66.030 161.985 ;
        RECT 65.820 161.450 65.960 161.615 ;
        RECT 63.920 161.130 64.180 161.450 ;
        RECT 64.380 161.130 64.640 161.450 ;
        RECT 65.760 161.130 66.020 161.450 ;
        RECT 64.440 159.750 64.580 161.130 ;
        RECT 61.620 159.430 61.880 159.750 ;
        RECT 64.380 159.430 64.640 159.750 ;
        RECT 61.680 159.150 61.820 159.430 ;
        RECT 61.680 159.010 63.200 159.150 ;
        RECT 54.260 157.730 55.380 157.850 ;
        RECT 45.275 157.195 46.815 157.565 ;
        RECT 46.960 157.030 47.100 157.710 ;
        RECT 49.260 157.030 49.400 157.730 ;
        RECT 54.320 157.710 55.380 157.730 ;
        RECT 61.220 157.710 62.280 157.850 ;
        RECT 46.900 156.710 47.160 157.030 ;
        RECT 49.200 156.710 49.460 157.030 ;
        RECT 55.240 156.010 55.380 157.710 ;
        RECT 41.840 155.690 42.100 156.010 ;
        RECT 55.180 155.690 55.440 156.010 ;
        RECT 62.140 155.670 62.280 157.710 ;
        RECT 63.060 156.010 63.200 159.010 ;
        RECT 63.785 157.195 65.325 157.565 ;
        RECT 63.000 155.690 63.260 156.010 ;
        RECT 34.020 155.350 34.280 155.670 ;
        RECT 62.080 155.350 62.340 155.670 ;
        RECT 36.020 154.475 37.560 154.845 ;
        RECT 54.530 154.475 56.070 154.845 ;
        RECT 26.765 151.755 28.305 152.125 ;
        RECT 45.275 151.755 46.815 152.125 ;
        RECT 63.060 150.910 63.200 155.690 ;
        RECT 63.785 151.755 65.325 152.125 ;
        RECT 66.280 150.990 66.420 167.250 ;
        RECT 67.200 166.630 67.340 183.490 ;
        RECT 67.660 170.630 67.800 199.210 ;
        RECT 68.060 198.530 68.320 198.850 ;
        RECT 67.600 170.310 67.860 170.630 ;
        RECT 68.120 166.890 68.260 198.530 ;
        RECT 71.740 196.490 72.000 196.810 ;
        RECT 68.520 193.090 68.780 193.410 ;
        RECT 68.580 191.710 68.720 193.090 ;
        RECT 71.800 192.390 71.940 196.490 ;
        RECT 71.740 192.070 72.000 192.390 ;
        RECT 68.520 191.390 68.780 191.710 ;
        RECT 68.580 189.330 68.720 191.390 ;
        RECT 72.720 190.690 72.860 205.670 ;
        RECT 75.420 203.970 75.680 204.290 ;
        RECT 73.040 203.435 74.580 203.805 ;
        RECT 75.480 203.270 75.620 203.970 ;
        RECT 75.420 202.950 75.680 203.270 ;
        RECT 74.960 199.210 75.220 199.530 ;
        RECT 73.040 197.995 74.580 198.365 ;
        RECT 75.020 197.150 75.160 199.210 ;
        RECT 74.960 196.830 75.220 197.150 ;
        RECT 74.960 195.810 75.220 196.130 ;
        RECT 75.020 193.750 75.160 195.810 ;
        RECT 74.960 193.430 75.220 193.750 ;
        RECT 75.480 193.150 75.620 202.950 ;
        RECT 75.880 202.270 76.140 202.590 ;
        RECT 75.940 200.550 76.080 202.270 ;
        RECT 75.880 200.230 76.140 200.550 ;
        RECT 76.400 199.530 76.540 206.690 ;
        RECT 77.780 204.970 77.920 208.180 ;
        RECT 82.295 206.155 83.835 206.525 ;
        RECT 79.560 205.330 79.820 205.650 ;
        RECT 77.720 204.650 77.980 204.970 ;
        RECT 76.800 203.970 77.060 204.290 ;
        RECT 79.100 203.970 79.360 204.290 ;
        RECT 76.860 200.210 77.000 203.970 ;
        RECT 77.720 201.250 77.980 201.570 ;
        RECT 76.800 199.890 77.060 200.210 ;
        RECT 76.340 199.210 76.600 199.530 ;
        RECT 76.400 194.510 76.540 199.210 ;
        RECT 75.020 193.010 75.620 193.150 ;
        RECT 75.940 194.370 76.540 194.510 ;
        RECT 73.040 192.555 74.580 192.925 ;
        RECT 72.660 190.370 72.920 190.690 ;
        RECT 75.020 189.670 75.160 193.010 ;
        RECT 75.940 189.670 76.080 194.370 ;
        RECT 76.340 193.770 76.600 194.090 ;
        RECT 76.400 191.710 76.540 193.770 ;
        RECT 76.340 191.390 76.600 191.710 ;
        RECT 74.960 189.350 75.220 189.670 ;
        RECT 75.880 189.350 76.140 189.670 ;
        RECT 68.520 189.010 68.780 189.330 ;
        RECT 68.580 185.250 68.720 189.010 ;
        RECT 68.980 187.990 69.240 188.310 ;
        RECT 69.040 186.610 69.180 187.990 ;
        RECT 71.280 187.650 71.540 187.970 ;
        RECT 72.200 187.650 72.460 187.970 ;
        RECT 72.660 187.650 72.920 187.970 ;
        RECT 68.980 186.290 69.240 186.610 ;
        RECT 68.520 184.930 68.780 185.250 ;
        RECT 69.040 180.830 69.180 186.290 ;
        RECT 71.340 186.270 71.480 187.650 ;
        RECT 71.280 185.950 71.540 186.270 ;
        RECT 69.900 185.610 70.160 185.930 ;
        RECT 69.960 183.210 70.100 185.610 ;
        RECT 70.820 184.930 71.080 185.250 ;
        RECT 70.880 183.550 71.020 184.930 ;
        RECT 70.820 183.230 71.080 183.550 ;
        RECT 69.900 182.890 70.160 183.210 ;
        RECT 72.260 182.870 72.400 187.650 ;
        RECT 72.720 183.210 72.860 187.650 ;
        RECT 73.040 187.115 74.580 187.485 ;
        RECT 75.020 185.930 75.160 189.350 ;
        RECT 75.420 187.650 75.680 187.970 ;
        RECT 75.480 186.270 75.620 187.650 ;
        RECT 75.420 185.950 75.680 186.270 ;
        RECT 74.960 185.610 75.220 185.930 ;
        RECT 72.660 182.890 72.920 183.210 ;
        RECT 72.200 182.550 72.460 182.870 ;
        RECT 73.040 181.675 74.580 182.045 ;
        RECT 75.480 180.830 75.620 185.950 ;
        RECT 68.980 180.510 69.240 180.830 ;
        RECT 75.420 180.510 75.680 180.830 ;
        RECT 68.520 176.770 68.780 177.090 ;
        RECT 68.580 175.390 68.720 176.770 ;
        RECT 69.040 176.070 69.180 180.510 ;
        RECT 73.120 180.170 73.380 180.490 ;
        RECT 69.440 177.110 69.700 177.430 ;
        RECT 72.660 177.110 72.920 177.430 ;
        RECT 68.980 175.750 69.240 176.070 ;
        RECT 68.520 175.070 68.780 175.390 ;
        RECT 68.580 169.950 68.720 175.070 ;
        RECT 69.040 174.710 69.180 175.750 ;
        RECT 69.500 175.390 69.640 177.110 ;
        RECT 69.900 176.770 70.160 177.090 ;
        RECT 69.960 175.390 70.100 176.770 ;
        RECT 72.720 176.070 72.860 177.110 ;
        RECT 73.180 177.090 73.320 180.170 ;
        RECT 75.420 179.490 75.680 179.810 ;
        RECT 73.120 176.770 73.380 177.090 ;
        RECT 73.040 176.235 74.580 176.605 ;
        RECT 72.660 175.750 72.920 176.070 ;
        RECT 75.480 175.390 75.620 179.490 ;
        RECT 69.440 175.070 69.700 175.390 ;
        RECT 69.900 175.070 70.160 175.390 ;
        RECT 75.420 175.070 75.680 175.390 ;
        RECT 68.980 174.390 69.240 174.710 ;
        RECT 71.740 174.390 72.000 174.710 ;
        RECT 71.800 173.350 71.940 174.390 ;
        RECT 71.740 173.030 72.000 173.350 ;
        RECT 75.420 171.330 75.680 171.650 ;
        RECT 73.040 170.795 74.580 171.165 ;
        RECT 75.480 169.950 75.620 171.330 ;
        RECT 75.940 170.290 76.080 189.350 ;
        RECT 76.860 177.430 77.000 199.890 ;
        RECT 77.260 196.490 77.520 196.810 ;
        RECT 77.320 183.745 77.460 196.490 ;
        RECT 77.780 185.930 77.920 201.250 ;
        RECT 79.160 197.830 79.300 203.970 ;
        RECT 79.620 202.590 79.760 205.330 ;
        RECT 84.220 204.970 84.360 208.180 ;
        RECT 90.660 204.970 90.800 208.180 ;
        RECT 81.400 204.650 81.660 204.970 ;
        RECT 84.160 204.650 84.420 204.970 ;
        RECT 90.600 204.650 90.860 204.970 ;
        RECT 81.460 203.270 81.600 204.650 ;
        RECT 81.860 203.970 82.120 204.290 ;
        RECT 84.620 203.970 84.880 204.290 ;
        RECT 86.460 203.970 86.720 204.290 ;
        RECT 81.400 202.950 81.660 203.270 ;
        RECT 79.560 202.270 79.820 202.590 ;
        RECT 80.020 202.270 80.280 202.590 ;
        RECT 80.480 202.270 80.740 202.590 ;
        RECT 80.940 202.270 81.200 202.590 ;
        RECT 79.620 199.870 79.760 202.270 ;
        RECT 79.560 199.550 79.820 199.870 ;
        RECT 79.100 197.510 79.360 197.830 ;
        RECT 78.640 196.830 78.900 197.150 ;
        RECT 78.700 194.770 78.840 196.830 ;
        RECT 78.640 194.450 78.900 194.770 ;
        RECT 78.700 186.270 78.840 194.450 ;
        RECT 79.160 186.950 79.300 197.510 ;
        RECT 80.080 194.000 80.220 202.270 ;
        RECT 80.540 196.550 80.680 202.270 ;
        RECT 81.000 200.550 81.140 202.270 ;
        RECT 80.940 200.230 81.200 200.550 ;
        RECT 81.920 199.530 82.060 203.970 ;
        RECT 84.160 201.930 84.420 202.250 ;
        RECT 82.295 200.715 83.835 201.085 ;
        RECT 84.220 200.550 84.360 201.930 ;
        RECT 84.160 200.230 84.420 200.550 ;
        RECT 84.680 199.950 84.820 203.970 ;
        RECT 85.540 201.250 85.800 201.570 ;
        RECT 84.220 199.810 84.820 199.950 ;
        RECT 81.860 199.210 82.120 199.530 ;
        RECT 81.860 198.530 82.120 198.850 ;
        RECT 82.320 198.530 82.580 198.850 ;
        RECT 80.540 196.410 81.140 196.550 ;
        RECT 80.480 195.810 80.740 196.130 ;
        RECT 80.540 195.110 80.680 195.810 ;
        RECT 80.480 194.790 80.740 195.110 ;
        RECT 80.480 194.000 80.740 194.090 ;
        RECT 80.080 193.945 80.740 194.000 ;
        RECT 80.080 193.860 80.750 193.945 ;
        RECT 80.470 193.575 80.750 193.860 ;
        RECT 81.000 193.750 81.140 196.410 ;
        RECT 80.940 193.430 81.200 193.750 ;
        RECT 81.000 192.390 81.140 193.430 ;
        RECT 81.920 192.470 82.060 198.530 ;
        RECT 82.380 196.810 82.520 198.530 ;
        RECT 84.220 197.490 84.360 199.810 ;
        RECT 84.620 199.210 84.880 199.530 ;
        RECT 84.680 197.830 84.820 199.210 ;
        RECT 84.620 197.510 84.880 197.830 ;
        RECT 84.160 197.230 84.420 197.490 ;
        RECT 84.160 197.170 84.820 197.230 ;
        RECT 84.220 197.090 84.820 197.170 ;
        RECT 85.600 197.150 85.740 201.250 ;
        RECT 86.520 197.150 86.660 203.970 ;
        RECT 91.550 203.435 93.090 203.805 ;
        RECT 90.590 202.415 90.870 202.785 ;
        RECT 90.600 202.270 90.860 202.415 ;
        RECT 90.660 199.870 90.800 202.270 ;
        RECT 90.600 199.550 90.860 199.870 ;
        RECT 91.550 197.995 93.090 198.365 ;
        RECT 82.320 196.490 82.580 196.810 ;
        RECT 84.160 196.490 84.420 196.810 ;
        RECT 82.295 195.275 83.835 195.645 ;
        RECT 84.220 195.110 84.360 196.490 ;
        RECT 84.160 194.790 84.420 195.110 ;
        RECT 84.160 193.770 84.420 194.090 ;
        RECT 82.780 193.430 83.040 193.750 ;
        RECT 82.840 193.265 82.980 193.430 ;
        RECT 83.240 193.320 83.500 193.410 ;
        RECT 84.220 193.320 84.360 193.770 ;
        RECT 82.770 192.895 83.050 193.265 ;
        RECT 83.240 193.180 84.360 193.320 ;
        RECT 83.240 193.090 83.500 193.180 ;
        RECT 80.940 192.070 81.200 192.390 ;
        RECT 81.460 192.330 82.060 192.470 ;
        RECT 79.100 186.630 79.360 186.950 ;
        RECT 78.640 185.950 78.900 186.270 ;
        RECT 80.020 185.950 80.280 186.270 ;
        RECT 80.480 185.950 80.740 186.270 ;
        RECT 77.720 185.610 77.980 185.930 ;
        RECT 77.250 183.375 77.530 183.745 ;
        RECT 77.780 181.590 77.920 185.610 ;
        RECT 77.320 181.450 77.920 181.590 ;
        RECT 76.800 177.110 77.060 177.430 ;
        RECT 77.320 173.010 77.460 181.450 ;
        RECT 78.700 180.830 78.840 185.950 ;
        RECT 80.080 184.230 80.220 185.950 ;
        RECT 80.020 183.910 80.280 184.230 ;
        RECT 77.720 180.510 77.980 180.830 ;
        RECT 78.640 180.510 78.900 180.830 ;
        RECT 77.780 178.450 77.920 180.510 ;
        RECT 77.720 178.130 77.980 178.450 ;
        RECT 77.710 175.215 77.990 175.585 ;
        RECT 78.700 175.390 78.840 180.510 ;
        RECT 80.540 178.190 80.680 185.950 ;
        RECT 81.460 185.450 81.600 192.330 ;
        RECT 81.860 191.390 82.120 191.710 ;
        RECT 81.920 186.270 82.060 191.390 ;
        RECT 82.295 189.835 83.835 190.205 ;
        RECT 81.860 185.950 82.120 186.270 ;
        RECT 83.700 185.610 83.960 185.930 ;
        RECT 83.760 185.450 83.900 185.610 ;
        RECT 84.680 185.450 84.820 197.090 ;
        RECT 85.540 196.830 85.800 197.150 ;
        RECT 86.460 196.830 86.720 197.150 ;
        RECT 87.840 196.830 88.100 197.150 ;
        RECT 85.080 195.810 85.340 196.130 ;
        RECT 86.460 195.810 86.720 196.130 ;
        RECT 85.140 191.710 85.280 195.810 ;
        RECT 86.520 194.140 86.660 195.810 ;
        RECT 86.460 193.820 86.720 194.140 ;
        RECT 87.900 194.090 88.040 196.830 ;
        RECT 86.920 193.770 87.180 194.090 ;
        RECT 87.840 193.945 88.100 194.090 ;
        RECT 85.540 193.265 85.800 193.410 ;
        RECT 85.530 192.895 85.810 193.265 ;
        RECT 86.980 192.390 87.120 193.770 ;
        RECT 87.830 193.575 88.110 193.945 ;
        RECT 90.600 193.430 90.860 193.750 ;
        RECT 87.840 193.090 88.100 193.410 ;
        RECT 86.920 192.070 87.180 192.390 ;
        RECT 85.080 191.390 85.340 191.710 ;
        RECT 86.000 191.050 86.260 191.370 ;
        RECT 81.460 185.310 82.060 185.450 ;
        RECT 83.760 185.310 84.360 185.450 ;
        RECT 84.680 185.310 85.280 185.450 ;
        RECT 80.080 178.050 80.680 178.190 ;
        RECT 80.080 176.070 80.220 178.050 ;
        RECT 80.480 177.450 80.740 177.770 ;
        RECT 80.020 175.980 80.280 176.070 ;
        RECT 79.620 175.840 80.280 175.980 ;
        RECT 77.720 175.070 77.980 175.215 ;
        RECT 78.640 175.070 78.900 175.390 ;
        RECT 77.260 172.690 77.520 173.010 ;
        RECT 75.880 169.970 76.140 170.290 ;
        RECT 68.520 169.630 68.780 169.950 ;
        RECT 72.200 169.630 72.460 169.950 ;
        RECT 75.420 169.630 75.680 169.950 ;
        RECT 66.740 166.490 67.340 166.630 ;
        RECT 68.060 166.570 68.320 166.890 ;
        RECT 68.580 166.550 68.720 169.630 ;
        RECT 70.360 167.590 70.620 167.910 ;
        RECT 66.740 162.130 66.880 166.490 ;
        RECT 68.520 166.230 68.780 166.550 ;
        RECT 70.420 162.470 70.560 167.590 ;
        RECT 70.820 166.230 71.080 166.550 ;
        RECT 70.880 165.190 71.020 166.230 ;
        RECT 71.740 165.890 72.000 166.210 ;
        RECT 70.820 164.870 71.080 165.190 ;
        RECT 70.360 162.150 70.620 162.470 ;
        RECT 66.680 161.810 66.940 162.130 ;
        RECT 66.740 161.110 66.880 161.810 ;
        RECT 71.800 161.450 71.940 165.890 ;
        RECT 72.260 162.550 72.400 169.630 ;
        RECT 74.960 169.290 75.220 169.610 ;
        RECT 77.320 169.350 77.460 172.690 ;
        RECT 78.700 172.330 78.840 175.070 ;
        RECT 78.640 172.010 78.900 172.330 ;
        RECT 78.700 170.290 78.840 172.010 ;
        RECT 78.640 169.970 78.900 170.290 ;
        RECT 78.180 169.630 78.440 169.950 ;
        RECT 72.660 166.570 72.920 166.890 ;
        RECT 72.720 164.850 72.860 166.570 ;
        RECT 73.040 165.355 74.580 165.725 ;
        RECT 72.660 164.530 72.920 164.850 ;
        RECT 75.020 164.750 75.160 169.290 ;
        RECT 76.860 169.210 77.460 169.350 ;
        RECT 76.860 167.910 77.000 169.210 ;
        RECT 77.260 168.610 77.520 168.930 ;
        RECT 76.800 167.590 77.060 167.910 ;
        RECT 76.330 166.375 76.610 166.745 ;
        RECT 75.020 164.610 76.080 164.750 ;
        RECT 72.260 162.410 72.860 162.550 ;
        RECT 72.720 161.450 72.860 162.410 ;
        RECT 75.940 162.130 76.080 164.610 ;
        RECT 75.880 161.810 76.140 162.130 ;
        RECT 71.740 161.130 72.000 161.450 ;
        RECT 72.660 161.130 72.920 161.450 ;
        RECT 66.680 160.790 66.940 161.110 ;
        RECT 67.140 160.450 67.400 160.770 ;
        RECT 71.280 160.450 71.540 160.770 ;
        RECT 72.200 160.450 72.460 160.770 ;
        RECT 67.200 158.730 67.340 160.450 ;
        RECT 71.340 158.730 71.480 160.450 ;
        RECT 72.260 159.750 72.400 160.450 ;
        RECT 73.040 159.915 74.580 160.285 ;
        RECT 72.200 159.430 72.460 159.750 ;
        RECT 75.940 159.070 76.080 161.810 ;
        RECT 76.400 159.750 76.540 166.375 ;
        RECT 76.860 166.210 77.000 167.590 ;
        RECT 76.800 165.890 77.060 166.210 ;
        RECT 77.320 161.450 77.460 168.610 ;
        RECT 77.720 166.570 77.980 166.890 ;
        RECT 77.780 165.190 77.920 166.570 ;
        RECT 78.240 166.550 78.380 169.630 ;
        RECT 79.100 169.290 79.360 169.610 ;
        RECT 78.640 168.610 78.900 168.930 ;
        RECT 78.180 166.230 78.440 166.550 ;
        RECT 78.240 165.190 78.380 166.230 ;
        RECT 77.720 164.870 77.980 165.190 ;
        RECT 78.180 164.870 78.440 165.190 ;
        RECT 77.780 163.230 77.920 164.870 ;
        RECT 78.700 163.830 78.840 168.610 ;
        RECT 79.160 166.210 79.300 169.290 ;
        RECT 79.620 169.270 79.760 175.840 ;
        RECT 80.020 175.750 80.280 175.840 ;
        RECT 80.540 175.050 80.680 177.450 ;
        RECT 80.940 176.770 81.200 177.090 ;
        RECT 81.000 176.070 81.140 176.770 ;
        RECT 80.940 175.750 81.200 176.070 ;
        RECT 80.020 174.730 80.280 175.050 ;
        RECT 80.480 174.730 80.740 175.050 ;
        RECT 80.080 173.350 80.220 174.730 ;
        RECT 80.020 173.030 80.280 173.350 ;
        RECT 79.560 168.950 79.820 169.270 ;
        RECT 79.100 165.890 79.360 166.210 ;
        RECT 80.540 164.510 80.680 174.730 ;
        RECT 81.400 172.010 81.660 172.330 ;
        RECT 81.460 170.290 81.600 172.010 ;
        RECT 81.400 169.970 81.660 170.290 ;
        RECT 80.940 169.630 81.200 169.950 ;
        RECT 81.000 167.910 81.140 169.630 ;
        RECT 80.940 167.590 81.200 167.910 ;
        RECT 81.920 166.745 82.060 185.310 ;
        RECT 82.295 184.395 83.835 184.765 ;
        RECT 84.220 184.230 84.360 185.310 ;
        RECT 84.160 183.910 84.420 184.230 ;
        RECT 85.140 183.210 85.280 185.310 ;
        RECT 85.540 184.930 85.800 185.250 ;
        RECT 85.600 183.210 85.740 184.930 ;
        RECT 86.060 183.890 86.200 191.050 ;
        RECT 86.980 186.270 87.120 192.070 ;
        RECT 87.900 191.370 88.040 193.090 ;
        RECT 90.660 192.050 90.800 193.430 ;
        RECT 91.550 192.555 93.090 192.925 ;
        RECT 90.600 191.905 90.860 192.050 ;
        RECT 90.590 191.535 90.870 191.905 ;
        RECT 87.840 191.050 88.100 191.370 ;
        RECT 91.550 187.115 93.090 187.485 ;
        RECT 86.920 185.950 87.180 186.270 ;
        RECT 86.980 184.230 87.120 185.950 ;
        RECT 90.140 184.930 90.400 185.250 ;
        RECT 86.920 183.910 87.180 184.230 ;
        RECT 88.300 183.910 88.560 184.230 ;
        RECT 86.000 183.570 86.260 183.890 ;
        RECT 84.160 182.890 84.420 183.210 ;
        RECT 85.080 182.890 85.340 183.210 ;
        RECT 85.540 182.890 85.800 183.210 ;
        RECT 84.220 182.530 84.360 182.890 ;
        RECT 84.160 182.210 84.420 182.530 ;
        RECT 82.295 178.955 83.835 179.325 ;
        RECT 82.295 173.515 83.835 173.885 ;
        RECT 85.140 171.650 85.280 182.890 ;
        RECT 86.060 178.110 86.200 183.570 ;
        RECT 86.450 183.375 86.730 183.745 ;
        RECT 86.520 183.210 86.660 183.375 ;
        RECT 86.460 182.890 86.720 183.210 ;
        RECT 86.000 177.790 86.260 178.110 ;
        RECT 86.000 174.110 86.260 174.370 ;
        RECT 86.520 174.110 86.660 182.890 ;
        RECT 86.920 182.210 87.180 182.530 ;
        RECT 86.980 177.430 87.120 182.210 ;
        RECT 88.360 177.770 88.500 183.910 ;
        RECT 90.200 183.745 90.340 184.930 ;
        RECT 90.130 183.375 90.410 183.745 ;
        RECT 90.200 182.870 90.340 183.375 ;
        RECT 90.140 182.550 90.400 182.870 ;
        RECT 91.550 181.675 93.090 182.045 ;
        RECT 88.300 177.450 88.560 177.770 ;
        RECT 86.920 177.110 87.180 177.430 ;
        RECT 86.000 174.050 86.660 174.110 ;
        RECT 86.060 173.970 86.660 174.050 ;
        RECT 85.080 171.330 85.340 171.650 ;
        RECT 82.295 168.075 83.835 168.445 ;
        RECT 85.140 166.890 85.280 171.330 ;
        RECT 85.540 168.610 85.800 168.930 ;
        RECT 85.600 166.890 85.740 168.610 ;
        RECT 86.520 166.890 86.660 173.970 ;
        RECT 86.980 172.330 87.120 177.110 ;
        RECT 88.360 176.070 88.500 177.450 ;
        RECT 90.600 177.110 90.860 177.430 ;
        RECT 88.300 175.750 88.560 176.070 ;
        RECT 90.660 174.370 90.800 177.110 ;
        RECT 91.550 176.235 93.090 176.605 ;
        RECT 90.600 174.225 90.860 174.370 ;
        RECT 90.590 173.855 90.870 174.225 ;
        RECT 86.920 172.010 87.180 172.330 ;
        RECT 81.850 166.375 82.130 166.745 ;
        RECT 85.080 166.570 85.340 166.890 ;
        RECT 85.540 166.570 85.800 166.890 ;
        RECT 86.460 166.570 86.720 166.890 ;
        RECT 83.700 165.890 83.960 166.210 ;
        RECT 83.760 164.510 83.900 165.890 ;
        RECT 80.480 164.190 80.740 164.510 ;
        RECT 83.700 164.190 83.960 164.510 ;
        RECT 78.640 163.510 78.900 163.830 ;
        RECT 79.100 163.230 79.360 163.490 ;
        RECT 77.780 163.170 79.360 163.230 ;
        RECT 79.560 163.170 79.820 163.490 ;
        RECT 77.780 163.090 79.300 163.170 ;
        RECT 77.780 162.130 77.920 163.090 ;
        RECT 77.720 161.810 77.980 162.130 ;
        RECT 77.260 161.130 77.520 161.450 ;
        RECT 78.180 160.450 78.440 160.770 ;
        RECT 76.340 159.430 76.600 159.750 ;
        RECT 78.240 159.070 78.380 160.450 ;
        RECT 75.880 158.750 76.140 159.070 ;
        RECT 78.180 158.750 78.440 159.070 ;
        RECT 67.140 158.410 67.400 158.730 ;
        RECT 71.280 158.410 71.540 158.730 ;
        RECT 67.200 157.030 67.340 158.410 ;
        RECT 73.580 157.730 73.840 158.050 ;
        RECT 67.140 156.710 67.400 157.030 ;
        RECT 73.640 156.010 73.780 157.730 ;
        RECT 79.160 157.030 79.300 163.090 ;
        RECT 79.620 160.770 79.760 163.170 ;
        RECT 79.560 160.450 79.820 160.770 ;
        RECT 79.100 156.710 79.360 157.030 ;
        RECT 73.580 155.690 73.840 156.010 ;
        RECT 73.040 154.475 74.580 154.845 ;
        RECT 79.620 151.590 79.760 160.450 ;
        RECT 80.540 158.730 80.680 164.190 ;
        RECT 82.295 162.635 83.835 163.005 ;
        RECT 86.980 162.470 87.120 172.010 ;
        RECT 91.550 170.795 93.090 171.165 ;
        RECT 90.600 166.570 90.860 166.890 ;
        RECT 87.840 164.530 88.100 164.850 ;
        RECT 90.660 164.705 90.800 166.570 ;
        RECT 91.550 165.355 93.090 165.725 ;
        RECT 86.920 162.150 87.180 162.470 ;
        RECT 87.900 161.450 88.040 164.530 ;
        RECT 90.590 164.335 90.870 164.705 ;
        RECT 90.600 164.190 90.860 164.335 ;
        RECT 90.660 162.130 90.800 164.190 ;
        RECT 90.600 161.810 90.860 162.130 ;
        RECT 117.400 161.675 118.000 161.700 ;
        RECT 87.840 161.130 88.100 161.450 ;
        RECT 80.480 158.410 80.740 158.730 ;
        RECT 80.540 156.350 80.680 158.410 ;
        RECT 87.900 158.050 88.040 161.130 ;
        RECT 117.380 161.125 118.020 161.675 ;
        RECT 88.300 160.450 88.560 160.770 ;
        RECT 87.840 157.905 88.100 158.050 ;
        RECT 82.295 157.195 83.835 157.565 ;
        RECT 87.830 157.535 88.110 157.905 ;
        RECT 88.360 157.030 88.500 160.450 ;
        RECT 91.550 159.915 93.090 160.285 ;
        RECT 115.900 157.375 116.500 157.400 ;
        RECT 88.300 156.710 88.560 157.030 ;
        RECT 115.880 156.825 116.520 157.375 ;
        RECT 80.480 156.030 80.740 156.350 ;
        RECT 82.295 151.755 83.835 152.125 ;
        RECT 77.260 151.270 77.520 151.590 ;
        RECT 79.560 151.270 79.820 151.590 ;
        RECT 65.360 150.910 66.420 150.990 ;
        RECT 63.000 150.590 63.260 150.910 ;
        RECT 65.300 150.850 66.420 150.910 ;
        RECT 65.300 150.590 65.560 150.850 ;
        RECT 36.020 149.035 37.560 149.405 ;
        RECT 54.530 149.035 56.070 149.405 ;
        RECT 73.040 149.035 74.580 149.405 ;
        RECT 26.765 146.315 28.305 146.685 ;
        RECT 45.275 146.315 46.815 146.685 ;
        RECT 63.785 146.315 65.325 146.685 ;
        RECT 36.020 143.595 37.560 143.965 ;
        RECT 54.530 143.595 56.070 143.965 ;
        RECT 73.040 143.595 74.580 143.965 ;
        RECT 26.765 140.875 28.305 141.245 ;
        RECT 45.275 140.875 46.815 141.245 ;
        RECT 63.785 140.875 65.325 141.245 ;
        RECT 36.020 138.155 37.560 138.525 ;
        RECT 54.530 138.155 56.070 138.525 ;
        RECT 73.040 138.155 74.580 138.525 ;
        RECT 77.320 136.825 77.460 151.270 ;
        RECT 82.295 146.315 83.835 146.685 ;
        RECT 88.360 145.665 88.500 156.710 ;
        RECT 106.425 155.300 106.975 155.320 ;
        RECT 91.550 154.475 93.090 154.845 ;
        RECT 106.400 154.700 113.030 155.300 ;
        RECT 106.425 154.680 106.975 154.700 ;
        RECT 115.900 152.470 116.500 156.825 ;
        RECT 117.400 155.270 118.000 161.125 ;
        RECT 118.900 160.175 119.500 160.200 ;
        RECT 118.880 159.625 119.520 160.175 ;
        RECT 118.900 155.170 119.500 159.625 ;
        RECT 120.400 159.075 121.000 159.100 ;
        RECT 120.380 158.525 121.020 159.075 ;
        RECT 121.800 158.975 122.400 159.000 ;
        RECT 120.400 155.070 121.000 158.525 ;
        RECT 121.780 158.425 122.420 158.975 ;
        RECT 121.800 154.070 122.400 158.425 ;
        RECT 91.550 149.035 93.090 149.405 ;
        RECT 104.725 149.000 105.275 149.020 ;
        RECT 104.700 148.400 107.630 149.000 ;
        RECT 104.725 148.380 105.275 148.400 ;
        RECT 104.725 146.700 105.275 146.720 ;
        RECT 104.700 146.100 107.330 146.700 ;
        RECT 104.725 146.080 105.275 146.100 ;
        RECT 88.290 145.295 88.570 145.665 ;
        RECT 91.550 143.595 93.090 143.965 ;
        RECT 82.295 140.875 83.835 141.245 ;
        RECT 91.550 138.155 93.090 138.525 ;
        RECT 77.250 136.455 77.530 136.825 ;
        RECT 26.765 135.435 28.305 135.805 ;
        RECT 45.275 135.435 46.815 135.805 ;
        RECT 63.785 135.435 65.325 135.805 ;
        RECT 82.295 135.435 83.835 135.805 ;
        RECT 36.020 132.715 37.560 133.085 ;
        RECT 54.530 132.715 56.070 133.085 ;
        RECT 73.040 132.715 74.580 133.085 ;
        RECT 91.550 132.715 93.090 133.085 ;
        RECT 147.325 26.400 147.875 26.420 ;
        RECT 130.270 25.800 147.900 26.400 ;
        RECT 147.325 25.780 147.875 25.800 ;
      LAYER via2 ;
        RECT 26.795 206.200 27.075 206.480 ;
        RECT 27.195 206.200 27.475 206.480 ;
        RECT 27.595 206.200 27.875 206.480 ;
        RECT 27.995 206.200 28.275 206.480 ;
        RECT 45.305 206.200 45.585 206.480 ;
        RECT 45.705 206.200 45.985 206.480 ;
        RECT 46.105 206.200 46.385 206.480 ;
        RECT 46.505 206.200 46.785 206.480 ;
        RECT 26.795 200.760 27.075 201.040 ;
        RECT 27.195 200.760 27.475 201.040 ;
        RECT 27.595 200.760 27.875 201.040 ;
        RECT 27.995 200.760 28.275 201.040 ;
        RECT 36.050 203.480 36.330 203.760 ;
        RECT 36.450 203.480 36.730 203.760 ;
        RECT 36.850 203.480 37.130 203.760 ;
        RECT 37.250 203.480 37.530 203.760 ;
        RECT 26.795 195.320 27.075 195.600 ;
        RECT 27.195 195.320 27.475 195.600 ;
        RECT 27.595 195.320 27.875 195.600 ;
        RECT 27.995 195.320 28.275 195.600 ;
        RECT 26.795 189.880 27.075 190.160 ;
        RECT 27.195 189.880 27.475 190.160 ;
        RECT 27.595 189.880 27.875 190.160 ;
        RECT 27.995 189.880 28.275 190.160 ;
        RECT 26.795 184.440 27.075 184.720 ;
        RECT 27.195 184.440 27.475 184.720 ;
        RECT 27.595 184.440 27.875 184.720 ;
        RECT 27.995 184.440 28.275 184.720 ;
        RECT 26.795 179.000 27.075 179.280 ;
        RECT 27.195 179.000 27.475 179.280 ;
        RECT 27.595 179.000 27.875 179.280 ;
        RECT 27.995 179.000 28.275 179.280 ;
        RECT 26.795 173.560 27.075 173.840 ;
        RECT 27.195 173.560 27.475 173.840 ;
        RECT 27.595 173.560 27.875 173.840 ;
        RECT 27.995 173.560 28.275 173.840 ;
        RECT 36.050 198.040 36.330 198.320 ;
        RECT 36.450 198.040 36.730 198.320 ;
        RECT 36.850 198.040 37.130 198.320 ;
        RECT 37.250 198.040 37.530 198.320 ;
        RECT 36.050 192.600 36.330 192.880 ;
        RECT 36.450 192.600 36.730 192.880 ;
        RECT 36.850 192.600 37.130 192.880 ;
        RECT 37.250 192.600 37.530 192.880 ;
        RECT 33.090 186.140 33.370 186.420 ;
        RECT 26.795 168.120 27.075 168.400 ;
        RECT 27.195 168.120 27.475 168.400 ;
        RECT 27.595 168.120 27.875 168.400 ;
        RECT 27.995 168.120 28.275 168.400 ;
        RECT 45.305 200.760 45.585 201.040 ;
        RECT 45.705 200.760 45.985 201.040 ;
        RECT 46.105 200.760 46.385 201.040 ;
        RECT 46.505 200.760 46.785 201.040 ;
        RECT 63.815 206.200 64.095 206.480 ;
        RECT 64.215 206.200 64.495 206.480 ;
        RECT 64.615 206.200 64.895 206.480 ;
        RECT 65.015 206.200 65.295 206.480 ;
        RECT 36.050 187.160 36.330 187.440 ;
        RECT 36.450 187.160 36.730 187.440 ;
        RECT 36.850 187.160 37.130 187.440 ;
        RECT 37.250 187.160 37.530 187.440 ;
        RECT 35.850 186.140 36.130 186.420 ;
        RECT 26.795 162.680 27.075 162.960 ;
        RECT 27.195 162.680 27.475 162.960 ;
        RECT 27.595 162.680 27.875 162.960 ;
        RECT 27.995 162.680 28.275 162.960 ;
        RECT 26.795 157.240 27.075 157.520 ;
        RECT 27.195 157.240 27.475 157.520 ;
        RECT 27.595 157.240 27.875 157.520 ;
        RECT 27.995 157.240 28.275 157.520 ;
        RECT 38.610 186.140 38.890 186.420 ;
        RECT 38.150 185.460 38.430 185.740 ;
        RECT 36.050 181.720 36.330 182.000 ;
        RECT 36.450 181.720 36.730 182.000 ;
        RECT 36.850 181.720 37.130 182.000 ;
        RECT 37.250 181.720 37.530 182.000 ;
        RECT 36.050 176.280 36.330 176.560 ;
        RECT 36.450 176.280 36.730 176.560 ;
        RECT 36.850 176.280 37.130 176.560 ;
        RECT 37.250 176.280 37.530 176.560 ;
        RECT 40.450 185.460 40.730 185.740 ;
        RECT 36.050 170.840 36.330 171.120 ;
        RECT 36.450 170.840 36.730 171.120 ;
        RECT 36.850 170.840 37.130 171.120 ;
        RECT 37.250 170.840 37.530 171.120 ;
        RECT 45.305 195.320 45.585 195.600 ;
        RECT 45.705 195.320 45.985 195.600 ;
        RECT 46.105 195.320 46.385 195.600 ;
        RECT 46.505 195.320 46.785 195.600 ;
        RECT 41.830 186.140 42.110 186.420 ;
        RECT 45.305 189.880 45.585 190.160 ;
        RECT 45.705 189.880 45.985 190.160 ;
        RECT 46.105 189.880 46.385 190.160 ;
        RECT 46.505 189.880 46.785 190.160 ;
        RECT 45.305 184.440 45.585 184.720 ;
        RECT 45.705 184.440 45.985 184.720 ;
        RECT 46.105 184.440 46.385 184.720 ;
        RECT 46.505 184.440 46.785 184.720 ;
        RECT 45.305 179.000 45.585 179.280 ;
        RECT 45.705 179.000 45.985 179.280 ;
        RECT 46.105 179.000 46.385 179.280 ;
        RECT 46.505 179.000 46.785 179.280 ;
        RECT 36.050 165.400 36.330 165.680 ;
        RECT 36.450 165.400 36.730 165.680 ;
        RECT 36.850 165.400 37.130 165.680 ;
        RECT 37.250 165.400 37.530 165.680 ;
        RECT 47.350 175.260 47.630 175.540 ;
        RECT 45.305 173.560 45.585 173.840 ;
        RECT 45.705 173.560 45.985 173.840 ;
        RECT 46.105 173.560 46.385 173.840 ;
        RECT 46.505 173.560 46.785 173.840 ;
        RECT 54.560 203.480 54.840 203.760 ;
        RECT 54.960 203.480 55.240 203.760 ;
        RECT 55.360 203.480 55.640 203.760 ;
        RECT 55.760 203.480 56.040 203.760 ;
        RECT 54.560 198.040 54.840 198.320 ;
        RECT 54.960 198.040 55.240 198.320 ;
        RECT 55.360 198.040 55.640 198.320 ;
        RECT 55.760 198.040 56.040 198.320 ;
        RECT 54.560 192.600 54.840 192.880 ;
        RECT 54.960 192.600 55.240 192.880 ;
        RECT 55.360 192.600 55.640 192.880 ;
        RECT 55.760 192.600 56.040 192.880 ;
        RECT 54.560 187.160 54.840 187.440 ;
        RECT 54.960 187.160 55.240 187.440 ;
        RECT 55.360 187.160 55.640 187.440 ;
        RECT 55.760 187.160 56.040 187.440 ;
        RECT 54.560 181.720 54.840 182.000 ;
        RECT 54.960 181.720 55.240 182.000 ;
        RECT 55.360 181.720 55.640 182.000 ;
        RECT 55.760 181.720 56.040 182.000 ;
        RECT 45.305 168.120 45.585 168.400 ;
        RECT 45.705 168.120 45.985 168.400 ;
        RECT 46.105 168.120 46.385 168.400 ;
        RECT 46.505 168.120 46.785 168.400 ;
        RECT 54.560 176.280 54.840 176.560 ;
        RECT 54.960 176.280 55.240 176.560 ;
        RECT 55.360 176.280 55.640 176.560 ;
        RECT 55.760 176.280 56.040 176.560 ;
        RECT 54.560 170.840 54.840 171.120 ;
        RECT 54.960 170.840 55.240 171.120 ;
        RECT 55.360 170.840 55.640 171.120 ;
        RECT 55.760 170.840 56.040 171.120 ;
        RECT 45.305 162.680 45.585 162.960 ;
        RECT 45.705 162.680 45.985 162.960 ;
        RECT 46.105 162.680 46.385 162.960 ;
        RECT 46.505 162.680 46.785 162.960 ;
        RECT 36.050 159.960 36.330 160.240 ;
        RECT 36.450 159.960 36.730 160.240 ;
        RECT 36.850 159.960 37.130 160.240 ;
        RECT 37.250 159.960 37.530 160.240 ;
        RECT 54.710 166.420 54.990 166.700 ;
        RECT 54.560 165.400 54.840 165.680 ;
        RECT 54.960 165.400 55.240 165.680 ;
        RECT 55.360 165.400 55.640 165.680 ;
        RECT 55.760 165.400 56.040 165.680 ;
        RECT 54.560 159.960 54.840 160.240 ;
        RECT 54.960 159.960 55.240 160.240 ;
        RECT 55.360 159.960 55.640 160.240 ;
        RECT 55.760 159.960 56.040 160.240 ;
        RECT 63.815 200.760 64.095 201.040 ;
        RECT 64.215 200.760 64.495 201.040 ;
        RECT 64.615 200.760 64.895 201.040 ;
        RECT 65.015 200.760 65.295 201.040 ;
        RECT 63.815 195.320 64.095 195.600 ;
        RECT 64.215 195.320 64.495 195.600 ;
        RECT 64.615 195.320 64.895 195.600 ;
        RECT 65.015 195.320 65.295 195.600 ;
        RECT 63.815 189.880 64.095 190.160 ;
        RECT 64.215 189.880 64.495 190.160 ;
        RECT 64.615 189.880 64.895 190.160 ;
        RECT 65.015 189.880 65.295 190.160 ;
        RECT 62.070 175.260 62.350 175.540 ;
        RECT 59.770 161.660 60.050 161.940 ;
        RECT 63.815 184.440 64.095 184.720 ;
        RECT 64.215 184.440 64.495 184.720 ;
        RECT 64.615 184.440 64.895 184.720 ;
        RECT 65.015 184.440 65.295 184.720 ;
        RECT 63.815 179.000 64.095 179.280 ;
        RECT 64.215 179.000 64.495 179.280 ;
        RECT 64.615 179.000 64.895 179.280 ;
        RECT 65.015 179.000 65.295 179.280 ;
        RECT 63.450 175.260 63.730 175.540 ;
        RECT 63.815 173.560 64.095 173.840 ;
        RECT 64.215 173.560 64.495 173.840 ;
        RECT 64.615 173.560 64.895 173.840 ;
        RECT 65.015 173.560 65.295 173.840 ;
        RECT 63.815 168.120 64.095 168.400 ;
        RECT 64.215 168.120 64.495 168.400 ;
        RECT 64.615 168.120 64.895 168.400 ;
        RECT 65.015 168.120 65.295 168.400 ;
        RECT 63.815 162.680 64.095 162.960 ;
        RECT 64.215 162.680 64.495 162.960 ;
        RECT 64.615 162.680 64.895 162.960 ;
        RECT 65.015 162.680 65.295 162.960 ;
        RECT 65.750 161.660 66.030 161.940 ;
        RECT 45.305 157.240 45.585 157.520 ;
        RECT 45.705 157.240 45.985 157.520 ;
        RECT 46.105 157.240 46.385 157.520 ;
        RECT 46.505 157.240 46.785 157.520 ;
        RECT 63.815 157.240 64.095 157.520 ;
        RECT 64.215 157.240 64.495 157.520 ;
        RECT 64.615 157.240 64.895 157.520 ;
        RECT 65.015 157.240 65.295 157.520 ;
        RECT 36.050 154.520 36.330 154.800 ;
        RECT 36.450 154.520 36.730 154.800 ;
        RECT 36.850 154.520 37.130 154.800 ;
        RECT 37.250 154.520 37.530 154.800 ;
        RECT 54.560 154.520 54.840 154.800 ;
        RECT 54.960 154.520 55.240 154.800 ;
        RECT 55.360 154.520 55.640 154.800 ;
        RECT 55.760 154.520 56.040 154.800 ;
        RECT 26.795 151.800 27.075 152.080 ;
        RECT 27.195 151.800 27.475 152.080 ;
        RECT 27.595 151.800 27.875 152.080 ;
        RECT 27.995 151.800 28.275 152.080 ;
        RECT 45.305 151.800 45.585 152.080 ;
        RECT 45.705 151.800 45.985 152.080 ;
        RECT 46.105 151.800 46.385 152.080 ;
        RECT 46.505 151.800 46.785 152.080 ;
        RECT 63.815 151.800 64.095 152.080 ;
        RECT 64.215 151.800 64.495 152.080 ;
        RECT 64.615 151.800 64.895 152.080 ;
        RECT 65.015 151.800 65.295 152.080 ;
        RECT 73.070 203.480 73.350 203.760 ;
        RECT 73.470 203.480 73.750 203.760 ;
        RECT 73.870 203.480 74.150 203.760 ;
        RECT 74.270 203.480 74.550 203.760 ;
        RECT 73.070 198.040 73.350 198.320 ;
        RECT 73.470 198.040 73.750 198.320 ;
        RECT 73.870 198.040 74.150 198.320 ;
        RECT 74.270 198.040 74.550 198.320 ;
        RECT 82.325 206.200 82.605 206.480 ;
        RECT 82.725 206.200 83.005 206.480 ;
        RECT 83.125 206.200 83.405 206.480 ;
        RECT 83.525 206.200 83.805 206.480 ;
        RECT 73.070 192.600 73.350 192.880 ;
        RECT 73.470 192.600 73.750 192.880 ;
        RECT 73.870 192.600 74.150 192.880 ;
        RECT 74.270 192.600 74.550 192.880 ;
        RECT 73.070 187.160 73.350 187.440 ;
        RECT 73.470 187.160 73.750 187.440 ;
        RECT 73.870 187.160 74.150 187.440 ;
        RECT 74.270 187.160 74.550 187.440 ;
        RECT 73.070 181.720 73.350 182.000 ;
        RECT 73.470 181.720 73.750 182.000 ;
        RECT 73.870 181.720 74.150 182.000 ;
        RECT 74.270 181.720 74.550 182.000 ;
        RECT 73.070 176.280 73.350 176.560 ;
        RECT 73.470 176.280 73.750 176.560 ;
        RECT 73.870 176.280 74.150 176.560 ;
        RECT 74.270 176.280 74.550 176.560 ;
        RECT 73.070 170.840 73.350 171.120 ;
        RECT 73.470 170.840 73.750 171.120 ;
        RECT 73.870 170.840 74.150 171.120 ;
        RECT 74.270 170.840 74.550 171.120 ;
        RECT 82.325 200.760 82.605 201.040 ;
        RECT 82.725 200.760 83.005 201.040 ;
        RECT 83.125 200.760 83.405 201.040 ;
        RECT 83.525 200.760 83.805 201.040 ;
        RECT 80.470 193.620 80.750 193.900 ;
        RECT 91.580 203.480 91.860 203.760 ;
        RECT 91.980 203.480 92.260 203.760 ;
        RECT 92.380 203.480 92.660 203.760 ;
        RECT 92.780 203.480 93.060 203.760 ;
        RECT 90.590 202.460 90.870 202.740 ;
        RECT 91.580 198.040 91.860 198.320 ;
        RECT 91.980 198.040 92.260 198.320 ;
        RECT 92.380 198.040 92.660 198.320 ;
        RECT 92.780 198.040 93.060 198.320 ;
        RECT 82.325 195.320 82.605 195.600 ;
        RECT 82.725 195.320 83.005 195.600 ;
        RECT 83.125 195.320 83.405 195.600 ;
        RECT 83.525 195.320 83.805 195.600 ;
        RECT 82.770 192.940 83.050 193.220 ;
        RECT 77.250 183.420 77.530 183.700 ;
        RECT 77.710 175.260 77.990 175.540 ;
        RECT 82.325 189.880 82.605 190.160 ;
        RECT 82.725 189.880 83.005 190.160 ;
        RECT 83.125 189.880 83.405 190.160 ;
        RECT 83.525 189.880 83.805 190.160 ;
        RECT 85.530 192.940 85.810 193.220 ;
        RECT 87.830 193.620 88.110 193.900 ;
        RECT 73.070 165.400 73.350 165.680 ;
        RECT 73.470 165.400 73.750 165.680 ;
        RECT 73.870 165.400 74.150 165.680 ;
        RECT 74.270 165.400 74.550 165.680 ;
        RECT 76.330 166.420 76.610 166.700 ;
        RECT 73.070 159.960 73.350 160.240 ;
        RECT 73.470 159.960 73.750 160.240 ;
        RECT 73.870 159.960 74.150 160.240 ;
        RECT 74.270 159.960 74.550 160.240 ;
        RECT 82.325 184.440 82.605 184.720 ;
        RECT 82.725 184.440 83.005 184.720 ;
        RECT 83.125 184.440 83.405 184.720 ;
        RECT 83.525 184.440 83.805 184.720 ;
        RECT 91.580 192.600 91.860 192.880 ;
        RECT 91.980 192.600 92.260 192.880 ;
        RECT 92.380 192.600 92.660 192.880 ;
        RECT 92.780 192.600 93.060 192.880 ;
        RECT 90.590 191.580 90.870 191.860 ;
        RECT 91.580 187.160 91.860 187.440 ;
        RECT 91.980 187.160 92.260 187.440 ;
        RECT 92.380 187.160 92.660 187.440 ;
        RECT 92.780 187.160 93.060 187.440 ;
        RECT 82.325 179.000 82.605 179.280 ;
        RECT 82.725 179.000 83.005 179.280 ;
        RECT 83.125 179.000 83.405 179.280 ;
        RECT 83.525 179.000 83.805 179.280 ;
        RECT 82.325 173.560 82.605 173.840 ;
        RECT 82.725 173.560 83.005 173.840 ;
        RECT 83.125 173.560 83.405 173.840 ;
        RECT 83.525 173.560 83.805 173.840 ;
        RECT 86.450 183.420 86.730 183.700 ;
        RECT 90.130 183.420 90.410 183.700 ;
        RECT 91.580 181.720 91.860 182.000 ;
        RECT 91.980 181.720 92.260 182.000 ;
        RECT 92.380 181.720 92.660 182.000 ;
        RECT 92.780 181.720 93.060 182.000 ;
        RECT 82.325 168.120 82.605 168.400 ;
        RECT 82.725 168.120 83.005 168.400 ;
        RECT 83.125 168.120 83.405 168.400 ;
        RECT 83.525 168.120 83.805 168.400 ;
        RECT 91.580 176.280 91.860 176.560 ;
        RECT 91.980 176.280 92.260 176.560 ;
        RECT 92.380 176.280 92.660 176.560 ;
        RECT 92.780 176.280 93.060 176.560 ;
        RECT 90.590 173.900 90.870 174.180 ;
        RECT 81.850 166.420 82.130 166.700 ;
        RECT 73.070 154.520 73.350 154.800 ;
        RECT 73.470 154.520 73.750 154.800 ;
        RECT 73.870 154.520 74.150 154.800 ;
        RECT 74.270 154.520 74.550 154.800 ;
        RECT 82.325 162.680 82.605 162.960 ;
        RECT 82.725 162.680 83.005 162.960 ;
        RECT 83.125 162.680 83.405 162.960 ;
        RECT 83.525 162.680 83.805 162.960 ;
        RECT 91.580 170.840 91.860 171.120 ;
        RECT 91.980 170.840 92.260 171.120 ;
        RECT 92.380 170.840 92.660 171.120 ;
        RECT 92.780 170.840 93.060 171.120 ;
        RECT 91.580 165.400 91.860 165.680 ;
        RECT 91.980 165.400 92.260 165.680 ;
        RECT 92.380 165.400 92.660 165.680 ;
        RECT 92.780 165.400 93.060 165.680 ;
        RECT 90.590 164.380 90.870 164.660 ;
        RECT 117.425 161.125 117.975 161.675 ;
        RECT 87.830 157.580 88.110 157.860 ;
        RECT 82.325 157.240 82.605 157.520 ;
        RECT 82.725 157.240 83.005 157.520 ;
        RECT 83.125 157.240 83.405 157.520 ;
        RECT 83.525 157.240 83.805 157.520 ;
        RECT 91.580 159.960 91.860 160.240 ;
        RECT 91.980 159.960 92.260 160.240 ;
        RECT 92.380 159.960 92.660 160.240 ;
        RECT 92.780 159.960 93.060 160.240 ;
        RECT 115.925 156.825 116.475 157.375 ;
        RECT 82.325 151.800 82.605 152.080 ;
        RECT 82.725 151.800 83.005 152.080 ;
        RECT 83.125 151.800 83.405 152.080 ;
        RECT 83.525 151.800 83.805 152.080 ;
        RECT 36.050 149.080 36.330 149.360 ;
        RECT 36.450 149.080 36.730 149.360 ;
        RECT 36.850 149.080 37.130 149.360 ;
        RECT 37.250 149.080 37.530 149.360 ;
        RECT 54.560 149.080 54.840 149.360 ;
        RECT 54.960 149.080 55.240 149.360 ;
        RECT 55.360 149.080 55.640 149.360 ;
        RECT 55.760 149.080 56.040 149.360 ;
        RECT 73.070 149.080 73.350 149.360 ;
        RECT 73.470 149.080 73.750 149.360 ;
        RECT 73.870 149.080 74.150 149.360 ;
        RECT 74.270 149.080 74.550 149.360 ;
        RECT 26.795 146.360 27.075 146.640 ;
        RECT 27.195 146.360 27.475 146.640 ;
        RECT 27.595 146.360 27.875 146.640 ;
        RECT 27.995 146.360 28.275 146.640 ;
        RECT 45.305 146.360 45.585 146.640 ;
        RECT 45.705 146.360 45.985 146.640 ;
        RECT 46.105 146.360 46.385 146.640 ;
        RECT 46.505 146.360 46.785 146.640 ;
        RECT 63.815 146.360 64.095 146.640 ;
        RECT 64.215 146.360 64.495 146.640 ;
        RECT 64.615 146.360 64.895 146.640 ;
        RECT 65.015 146.360 65.295 146.640 ;
        RECT 36.050 143.640 36.330 143.920 ;
        RECT 36.450 143.640 36.730 143.920 ;
        RECT 36.850 143.640 37.130 143.920 ;
        RECT 37.250 143.640 37.530 143.920 ;
        RECT 54.560 143.640 54.840 143.920 ;
        RECT 54.960 143.640 55.240 143.920 ;
        RECT 55.360 143.640 55.640 143.920 ;
        RECT 55.760 143.640 56.040 143.920 ;
        RECT 73.070 143.640 73.350 143.920 ;
        RECT 73.470 143.640 73.750 143.920 ;
        RECT 73.870 143.640 74.150 143.920 ;
        RECT 74.270 143.640 74.550 143.920 ;
        RECT 26.795 140.920 27.075 141.200 ;
        RECT 27.195 140.920 27.475 141.200 ;
        RECT 27.595 140.920 27.875 141.200 ;
        RECT 27.995 140.920 28.275 141.200 ;
        RECT 45.305 140.920 45.585 141.200 ;
        RECT 45.705 140.920 45.985 141.200 ;
        RECT 46.105 140.920 46.385 141.200 ;
        RECT 46.505 140.920 46.785 141.200 ;
        RECT 63.815 140.920 64.095 141.200 ;
        RECT 64.215 140.920 64.495 141.200 ;
        RECT 64.615 140.920 64.895 141.200 ;
        RECT 65.015 140.920 65.295 141.200 ;
        RECT 36.050 138.200 36.330 138.480 ;
        RECT 36.450 138.200 36.730 138.480 ;
        RECT 36.850 138.200 37.130 138.480 ;
        RECT 37.250 138.200 37.530 138.480 ;
        RECT 54.560 138.200 54.840 138.480 ;
        RECT 54.960 138.200 55.240 138.480 ;
        RECT 55.360 138.200 55.640 138.480 ;
        RECT 55.760 138.200 56.040 138.480 ;
        RECT 73.070 138.200 73.350 138.480 ;
        RECT 73.470 138.200 73.750 138.480 ;
        RECT 73.870 138.200 74.150 138.480 ;
        RECT 74.270 138.200 74.550 138.480 ;
        RECT 82.325 146.360 82.605 146.640 ;
        RECT 82.725 146.360 83.005 146.640 ;
        RECT 83.125 146.360 83.405 146.640 ;
        RECT 83.525 146.360 83.805 146.640 ;
        RECT 91.580 154.520 91.860 154.800 ;
        RECT 91.980 154.520 92.260 154.800 ;
        RECT 92.380 154.520 92.660 154.800 ;
        RECT 92.780 154.520 93.060 154.800 ;
        RECT 106.425 154.725 106.975 155.275 ;
        RECT 118.925 159.625 119.475 160.175 ;
        RECT 120.425 158.525 120.975 159.075 ;
        RECT 121.825 158.425 122.375 158.975 ;
        RECT 91.580 149.080 91.860 149.360 ;
        RECT 91.980 149.080 92.260 149.360 ;
        RECT 92.380 149.080 92.660 149.360 ;
        RECT 92.780 149.080 93.060 149.360 ;
        RECT 104.725 148.425 105.275 148.975 ;
        RECT 104.725 146.125 105.275 146.675 ;
        RECT 88.290 145.340 88.570 145.620 ;
        RECT 91.580 143.640 91.860 143.920 ;
        RECT 91.980 143.640 92.260 143.920 ;
        RECT 92.380 143.640 92.660 143.920 ;
        RECT 92.780 143.640 93.060 143.920 ;
        RECT 82.325 140.920 82.605 141.200 ;
        RECT 82.725 140.920 83.005 141.200 ;
        RECT 83.125 140.920 83.405 141.200 ;
        RECT 83.525 140.920 83.805 141.200 ;
        RECT 91.580 138.200 91.860 138.480 ;
        RECT 91.980 138.200 92.260 138.480 ;
        RECT 92.380 138.200 92.660 138.480 ;
        RECT 92.780 138.200 93.060 138.480 ;
        RECT 77.250 136.500 77.530 136.780 ;
        RECT 26.795 135.480 27.075 135.760 ;
        RECT 27.195 135.480 27.475 135.760 ;
        RECT 27.595 135.480 27.875 135.760 ;
        RECT 27.995 135.480 28.275 135.760 ;
        RECT 45.305 135.480 45.585 135.760 ;
        RECT 45.705 135.480 45.985 135.760 ;
        RECT 46.105 135.480 46.385 135.760 ;
        RECT 46.505 135.480 46.785 135.760 ;
        RECT 63.815 135.480 64.095 135.760 ;
        RECT 64.215 135.480 64.495 135.760 ;
        RECT 64.615 135.480 64.895 135.760 ;
        RECT 65.015 135.480 65.295 135.760 ;
        RECT 82.325 135.480 82.605 135.760 ;
        RECT 82.725 135.480 83.005 135.760 ;
        RECT 83.125 135.480 83.405 135.760 ;
        RECT 83.525 135.480 83.805 135.760 ;
        RECT 36.050 132.760 36.330 133.040 ;
        RECT 36.450 132.760 36.730 133.040 ;
        RECT 36.850 132.760 37.130 133.040 ;
        RECT 37.250 132.760 37.530 133.040 ;
        RECT 54.560 132.760 54.840 133.040 ;
        RECT 54.960 132.760 55.240 133.040 ;
        RECT 55.360 132.760 55.640 133.040 ;
        RECT 55.760 132.760 56.040 133.040 ;
        RECT 73.070 132.760 73.350 133.040 ;
        RECT 73.470 132.760 73.750 133.040 ;
        RECT 73.870 132.760 74.150 133.040 ;
        RECT 74.270 132.760 74.550 133.040 ;
        RECT 91.580 132.760 91.860 133.040 ;
        RECT 91.980 132.760 92.260 133.040 ;
        RECT 92.380 132.760 92.660 133.040 ;
        RECT 92.780 132.760 93.060 133.040 ;
        RECT 147.325 25.825 147.875 26.375 ;
      LAYER met3 ;
        RECT 26.745 206.175 28.325 206.505 ;
        RECT 45.255 206.175 46.835 206.505 ;
        RECT 63.765 206.175 65.345 206.505 ;
        RECT 82.275 206.175 83.855 206.505 ;
        RECT 36.000 203.455 37.580 203.785 ;
        RECT 54.510 203.455 56.090 203.785 ;
        RECT 73.020 203.455 74.600 203.785 ;
        RECT 91.530 203.455 93.110 203.785 ;
        RECT 90.565 202.750 90.895 202.765 ;
        RECT 93.520 202.750 122.400 202.900 ;
        RECT 90.565 202.450 122.400 202.750 ;
        RECT 90.565 202.435 90.895 202.450 ;
        RECT 93.520 202.300 122.400 202.450 ;
        RECT 26.745 200.735 28.325 201.065 ;
        RECT 45.255 200.735 46.835 201.065 ;
        RECT 63.765 200.735 65.345 201.065 ;
        RECT 82.275 200.735 83.855 201.065 ;
        RECT 36.000 198.015 37.580 198.345 ;
        RECT 54.510 198.015 56.090 198.345 ;
        RECT 73.020 198.015 74.600 198.345 ;
        RECT 91.530 198.015 93.110 198.345 ;
        RECT 26.745 195.295 28.325 195.625 ;
        RECT 45.255 195.295 46.835 195.625 ;
        RECT 63.765 195.295 65.345 195.625 ;
        RECT 82.275 195.295 83.855 195.625 ;
        RECT 80.445 193.910 80.775 193.925 ;
        RECT 87.805 193.910 88.135 193.925 ;
        RECT 80.445 193.610 88.135 193.910 ;
        RECT 80.445 193.595 80.775 193.610 ;
        RECT 87.805 193.595 88.135 193.610 ;
        RECT 82.745 193.230 83.075 193.245 ;
        RECT 85.505 193.230 85.835 193.245 ;
        RECT 82.745 192.930 85.835 193.230 ;
        RECT 82.745 192.915 83.075 192.930 ;
        RECT 85.505 192.915 85.835 192.930 ;
        RECT 36.000 192.575 37.580 192.905 ;
        RECT 54.510 192.575 56.090 192.905 ;
        RECT 73.020 192.575 74.600 192.905 ;
        RECT 91.530 192.575 93.110 192.905 ;
        RECT 93.520 192.780 121.000 193.380 ;
        RECT 90.565 191.870 90.895 191.885 ;
        RECT 94.030 191.870 94.330 192.780 ;
        RECT 90.565 191.570 94.330 191.870 ;
        RECT 90.565 191.555 90.895 191.570 ;
        RECT 26.745 189.855 28.325 190.185 ;
        RECT 45.255 189.855 46.835 190.185 ;
        RECT 63.765 189.855 65.345 190.185 ;
        RECT 82.275 189.855 83.855 190.185 ;
        RECT 36.000 187.135 37.580 187.465 ;
        RECT 54.510 187.135 56.090 187.465 ;
        RECT 73.020 187.135 74.600 187.465 ;
        RECT 91.530 187.135 93.110 187.465 ;
        RECT 33.065 186.430 33.395 186.445 ;
        RECT 35.825 186.430 36.155 186.445 ;
        RECT 38.585 186.430 38.915 186.445 ;
        RECT 41.805 186.430 42.135 186.445 ;
        RECT 33.065 186.130 42.135 186.430 ;
        RECT 33.065 186.115 33.395 186.130 ;
        RECT 35.825 186.115 36.155 186.130 ;
        RECT 38.585 186.115 38.915 186.130 ;
        RECT 41.805 186.115 42.135 186.130 ;
        RECT 38.125 185.750 38.455 185.765 ;
        RECT 40.425 185.750 40.755 185.765 ;
        RECT 38.125 185.450 40.755 185.750 ;
        RECT 38.125 185.435 38.455 185.450 ;
        RECT 40.425 185.435 40.755 185.450 ;
        RECT 26.745 184.415 28.325 184.745 ;
        RECT 45.255 184.415 46.835 184.745 ;
        RECT 63.765 184.415 65.345 184.745 ;
        RECT 82.275 184.415 83.855 184.745 ;
        RECT 77.225 183.710 77.555 183.725 ;
        RECT 86.425 183.710 86.755 183.725 ;
        RECT 77.225 183.410 86.755 183.710 ;
        RECT 77.225 183.395 77.555 183.410 ;
        RECT 86.425 183.395 86.755 183.410 ;
        RECT 90.105 183.710 90.435 183.725 ;
        RECT 93.520 183.710 119.500 183.860 ;
        RECT 90.105 183.410 119.500 183.710 ;
        RECT 90.105 183.395 90.435 183.410 ;
        RECT 93.520 183.260 119.500 183.410 ;
        RECT 36.000 181.695 37.580 182.025 ;
        RECT 54.510 181.695 56.090 182.025 ;
        RECT 73.020 181.695 74.600 182.025 ;
        RECT 91.530 181.695 93.110 182.025 ;
        RECT 26.745 178.975 28.325 179.305 ;
        RECT 45.255 178.975 46.835 179.305 ;
        RECT 63.765 178.975 65.345 179.305 ;
        RECT 82.275 178.975 83.855 179.305 ;
        RECT 36.000 176.255 37.580 176.585 ;
        RECT 54.510 176.255 56.090 176.585 ;
        RECT 73.020 176.255 74.600 176.585 ;
        RECT 91.530 176.255 93.110 176.585 ;
        RECT 47.325 175.550 47.655 175.565 ;
        RECT 62.045 175.550 62.375 175.565 ;
        RECT 63.425 175.550 63.755 175.565 ;
        RECT 77.685 175.550 78.015 175.565 ;
        RECT 47.325 175.250 78.015 175.550 ;
        RECT 47.325 175.235 47.655 175.250 ;
        RECT 62.045 175.235 62.375 175.250 ;
        RECT 63.425 175.235 63.755 175.250 ;
        RECT 77.685 175.235 78.015 175.250 ;
        RECT 90.565 174.190 90.895 174.205 ;
        RECT 93.520 174.190 118.000 174.340 ;
        RECT 90.565 173.890 118.000 174.190 ;
        RECT 90.565 173.875 90.895 173.890 ;
        RECT 26.745 173.535 28.325 173.865 ;
        RECT 45.255 173.535 46.835 173.865 ;
        RECT 63.765 173.535 65.345 173.865 ;
        RECT 82.275 173.535 83.855 173.865 ;
        RECT 93.520 173.740 118.000 173.890 ;
        RECT 36.000 170.815 37.580 171.145 ;
        RECT 54.510 170.815 56.090 171.145 ;
        RECT 73.020 170.815 74.600 171.145 ;
        RECT 91.530 170.815 93.110 171.145 ;
        RECT 26.745 168.095 28.325 168.425 ;
        RECT 45.255 168.095 46.835 168.425 ;
        RECT 63.765 168.095 65.345 168.425 ;
        RECT 82.275 168.095 83.855 168.425 ;
        RECT 54.685 166.710 55.015 166.725 ;
        RECT 76.305 166.710 76.635 166.725 ;
        RECT 81.825 166.710 82.155 166.725 ;
        RECT 54.685 166.410 82.155 166.710 ;
        RECT 54.685 166.395 55.015 166.410 ;
        RECT 76.305 166.395 76.635 166.410 ;
        RECT 81.825 166.395 82.155 166.410 ;
        RECT 36.000 165.375 37.580 165.705 ;
        RECT 54.510 165.375 56.090 165.705 ;
        RECT 73.020 165.375 74.600 165.705 ;
        RECT 91.530 165.375 93.110 165.705 ;
        RECT 90.565 164.670 90.895 164.685 ;
        RECT 93.520 164.670 116.500 164.820 ;
        RECT 90.565 164.370 116.500 164.670 ;
        RECT 90.565 164.355 90.895 164.370 ;
        RECT 93.520 164.220 116.500 164.370 ;
        RECT 26.745 162.655 28.325 162.985 ;
        RECT 45.255 162.655 46.835 162.985 ;
        RECT 63.765 162.655 65.345 162.985 ;
        RECT 82.275 162.655 83.855 162.985 ;
        RECT 59.745 161.950 60.075 161.965 ;
        RECT 65.725 161.950 66.055 161.965 ;
        RECT 59.745 161.650 66.055 161.950 ;
        RECT 59.745 161.635 60.075 161.650 ;
        RECT 65.725 161.635 66.055 161.650 ;
        RECT 36.000 159.935 37.580 160.265 ;
        RECT 54.510 159.935 56.090 160.265 ;
        RECT 73.020 159.935 74.600 160.265 ;
        RECT 91.530 159.935 93.110 160.265 ;
        RECT 87.805 157.870 88.135 157.885 ;
        RECT 87.805 157.570 94.330 157.870 ;
        RECT 87.805 157.555 88.135 157.570 ;
        RECT 26.745 157.215 28.325 157.545 ;
        RECT 45.255 157.215 46.835 157.545 ;
        RECT 63.765 157.215 65.345 157.545 ;
        RECT 82.275 157.215 83.855 157.545 ;
        RECT 94.030 155.300 94.330 157.570 ;
        RECT 115.900 156.800 116.500 164.220 ;
        RECT 117.400 161.100 118.000 173.740 ;
        RECT 118.900 159.600 119.500 183.260 ;
        RECT 120.400 158.500 121.000 192.780 ;
        RECT 121.800 158.400 122.400 202.300 ;
        RECT 36.000 154.495 37.580 154.825 ;
        RECT 54.510 154.495 56.090 154.825 ;
        RECT 73.020 154.495 74.600 154.825 ;
        RECT 91.530 154.495 93.110 154.825 ;
        RECT 93.520 154.700 107.000 155.300 ;
        RECT 26.745 151.775 28.325 152.105 ;
        RECT 45.255 151.775 46.835 152.105 ;
        RECT 63.765 151.775 65.345 152.105 ;
        RECT 82.275 151.775 83.855 152.105 ;
        RECT 36.000 149.055 37.580 149.385 ;
        RECT 54.510 149.055 56.090 149.385 ;
        RECT 73.020 149.055 74.600 149.385 ;
        RECT 91.530 149.055 93.110 149.385 ;
        RECT 99.100 148.400 105.300 149.000 ;
        RECT 26.745 146.335 28.325 146.665 ;
        RECT 45.255 146.335 46.835 146.665 ;
        RECT 63.765 146.335 65.345 146.665 ;
        RECT 82.275 146.335 83.855 146.665 ;
        RECT 99.100 145.780 99.700 148.400 ;
        RECT 88.265 145.630 88.595 145.645 ;
        RECT 93.520 145.630 99.700 145.780 ;
        RECT 88.265 145.330 99.700 145.630 ;
        RECT 88.265 145.315 88.595 145.330 ;
        RECT 93.520 145.180 99.700 145.330 ;
        RECT 36.000 143.615 37.580 143.945 ;
        RECT 54.510 143.615 56.090 143.945 ;
        RECT 73.020 143.615 74.600 143.945 ;
        RECT 91.530 143.615 93.110 143.945 ;
        RECT 26.745 140.895 28.325 141.225 ;
        RECT 45.255 140.895 46.835 141.225 ;
        RECT 63.765 140.895 65.345 141.225 ;
        RECT 82.275 140.895 83.855 141.225 ;
        RECT 36.000 138.175 37.580 138.505 ;
        RECT 54.510 138.175 56.090 138.505 ;
        RECT 73.020 138.175 74.600 138.505 ;
        RECT 91.530 138.175 93.110 138.505 ;
        RECT 77.225 136.790 77.555 136.805 ;
        RECT 77.225 136.490 85.130 136.790 ;
        RECT 77.225 136.475 77.555 136.490 ;
        RECT 84.830 136.110 85.130 136.490 ;
        RECT 104.700 136.260 105.300 146.700 ;
        RECT 93.520 136.110 105.300 136.260 ;
        RECT 84.830 135.810 105.300 136.110 ;
        RECT 26.745 135.455 28.325 135.785 ;
        RECT 45.255 135.455 46.835 135.785 ;
        RECT 63.765 135.455 65.345 135.785 ;
        RECT 82.275 135.455 83.855 135.785 ;
        RECT 93.520 135.660 105.300 135.810 ;
        RECT 36.000 132.735 37.580 133.065 ;
        RECT 54.510 132.735 56.090 133.065 ;
        RECT 73.020 132.735 74.600 133.065 ;
        RECT 91.530 132.735 93.110 133.065 ;
        RECT 156.565 26.400 157.155 26.425 ;
        RECT 147.300 25.800 157.160 26.400 ;
        RECT 156.565 25.775 157.155 25.800 ;
      LAYER via3 ;
        RECT 26.775 206.180 27.095 206.500 ;
        RECT 27.175 206.180 27.495 206.500 ;
        RECT 27.575 206.180 27.895 206.500 ;
        RECT 27.975 206.180 28.295 206.500 ;
        RECT 45.285 206.180 45.605 206.500 ;
        RECT 45.685 206.180 46.005 206.500 ;
        RECT 46.085 206.180 46.405 206.500 ;
        RECT 46.485 206.180 46.805 206.500 ;
        RECT 63.795 206.180 64.115 206.500 ;
        RECT 64.195 206.180 64.515 206.500 ;
        RECT 64.595 206.180 64.915 206.500 ;
        RECT 64.995 206.180 65.315 206.500 ;
        RECT 82.305 206.180 82.625 206.500 ;
        RECT 82.705 206.180 83.025 206.500 ;
        RECT 83.105 206.180 83.425 206.500 ;
        RECT 83.505 206.180 83.825 206.500 ;
        RECT 36.030 203.460 36.350 203.780 ;
        RECT 36.430 203.460 36.750 203.780 ;
        RECT 36.830 203.460 37.150 203.780 ;
        RECT 37.230 203.460 37.550 203.780 ;
        RECT 54.540 203.460 54.860 203.780 ;
        RECT 54.940 203.460 55.260 203.780 ;
        RECT 55.340 203.460 55.660 203.780 ;
        RECT 55.740 203.460 56.060 203.780 ;
        RECT 73.050 203.460 73.370 203.780 ;
        RECT 73.450 203.460 73.770 203.780 ;
        RECT 73.850 203.460 74.170 203.780 ;
        RECT 74.250 203.460 74.570 203.780 ;
        RECT 91.560 203.460 91.880 203.780 ;
        RECT 91.960 203.460 92.280 203.780 ;
        RECT 92.360 203.460 92.680 203.780 ;
        RECT 92.760 203.460 93.080 203.780 ;
        RECT 26.775 200.740 27.095 201.060 ;
        RECT 27.175 200.740 27.495 201.060 ;
        RECT 27.575 200.740 27.895 201.060 ;
        RECT 27.975 200.740 28.295 201.060 ;
        RECT 45.285 200.740 45.605 201.060 ;
        RECT 45.685 200.740 46.005 201.060 ;
        RECT 46.085 200.740 46.405 201.060 ;
        RECT 46.485 200.740 46.805 201.060 ;
        RECT 63.795 200.740 64.115 201.060 ;
        RECT 64.195 200.740 64.515 201.060 ;
        RECT 64.595 200.740 64.915 201.060 ;
        RECT 64.995 200.740 65.315 201.060 ;
        RECT 82.305 200.740 82.625 201.060 ;
        RECT 82.705 200.740 83.025 201.060 ;
        RECT 83.105 200.740 83.425 201.060 ;
        RECT 83.505 200.740 83.825 201.060 ;
        RECT 36.030 198.020 36.350 198.340 ;
        RECT 36.430 198.020 36.750 198.340 ;
        RECT 36.830 198.020 37.150 198.340 ;
        RECT 37.230 198.020 37.550 198.340 ;
        RECT 54.540 198.020 54.860 198.340 ;
        RECT 54.940 198.020 55.260 198.340 ;
        RECT 55.340 198.020 55.660 198.340 ;
        RECT 55.740 198.020 56.060 198.340 ;
        RECT 73.050 198.020 73.370 198.340 ;
        RECT 73.450 198.020 73.770 198.340 ;
        RECT 73.850 198.020 74.170 198.340 ;
        RECT 74.250 198.020 74.570 198.340 ;
        RECT 91.560 198.020 91.880 198.340 ;
        RECT 91.960 198.020 92.280 198.340 ;
        RECT 92.360 198.020 92.680 198.340 ;
        RECT 92.760 198.020 93.080 198.340 ;
        RECT 26.775 195.300 27.095 195.620 ;
        RECT 27.175 195.300 27.495 195.620 ;
        RECT 27.575 195.300 27.895 195.620 ;
        RECT 27.975 195.300 28.295 195.620 ;
        RECT 45.285 195.300 45.605 195.620 ;
        RECT 45.685 195.300 46.005 195.620 ;
        RECT 46.085 195.300 46.405 195.620 ;
        RECT 46.485 195.300 46.805 195.620 ;
        RECT 63.795 195.300 64.115 195.620 ;
        RECT 64.195 195.300 64.515 195.620 ;
        RECT 64.595 195.300 64.915 195.620 ;
        RECT 64.995 195.300 65.315 195.620 ;
        RECT 82.305 195.300 82.625 195.620 ;
        RECT 82.705 195.300 83.025 195.620 ;
        RECT 83.105 195.300 83.425 195.620 ;
        RECT 83.505 195.300 83.825 195.620 ;
        RECT 36.030 192.580 36.350 192.900 ;
        RECT 36.430 192.580 36.750 192.900 ;
        RECT 36.830 192.580 37.150 192.900 ;
        RECT 37.230 192.580 37.550 192.900 ;
        RECT 54.540 192.580 54.860 192.900 ;
        RECT 54.940 192.580 55.260 192.900 ;
        RECT 55.340 192.580 55.660 192.900 ;
        RECT 55.740 192.580 56.060 192.900 ;
        RECT 73.050 192.580 73.370 192.900 ;
        RECT 73.450 192.580 73.770 192.900 ;
        RECT 73.850 192.580 74.170 192.900 ;
        RECT 74.250 192.580 74.570 192.900 ;
        RECT 91.560 192.580 91.880 192.900 ;
        RECT 91.960 192.580 92.280 192.900 ;
        RECT 92.360 192.580 92.680 192.900 ;
        RECT 92.760 192.580 93.080 192.900 ;
        RECT 26.775 189.860 27.095 190.180 ;
        RECT 27.175 189.860 27.495 190.180 ;
        RECT 27.575 189.860 27.895 190.180 ;
        RECT 27.975 189.860 28.295 190.180 ;
        RECT 45.285 189.860 45.605 190.180 ;
        RECT 45.685 189.860 46.005 190.180 ;
        RECT 46.085 189.860 46.405 190.180 ;
        RECT 46.485 189.860 46.805 190.180 ;
        RECT 63.795 189.860 64.115 190.180 ;
        RECT 64.195 189.860 64.515 190.180 ;
        RECT 64.595 189.860 64.915 190.180 ;
        RECT 64.995 189.860 65.315 190.180 ;
        RECT 82.305 189.860 82.625 190.180 ;
        RECT 82.705 189.860 83.025 190.180 ;
        RECT 83.105 189.860 83.425 190.180 ;
        RECT 83.505 189.860 83.825 190.180 ;
        RECT 36.030 187.140 36.350 187.460 ;
        RECT 36.430 187.140 36.750 187.460 ;
        RECT 36.830 187.140 37.150 187.460 ;
        RECT 37.230 187.140 37.550 187.460 ;
        RECT 54.540 187.140 54.860 187.460 ;
        RECT 54.940 187.140 55.260 187.460 ;
        RECT 55.340 187.140 55.660 187.460 ;
        RECT 55.740 187.140 56.060 187.460 ;
        RECT 73.050 187.140 73.370 187.460 ;
        RECT 73.450 187.140 73.770 187.460 ;
        RECT 73.850 187.140 74.170 187.460 ;
        RECT 74.250 187.140 74.570 187.460 ;
        RECT 91.560 187.140 91.880 187.460 ;
        RECT 91.960 187.140 92.280 187.460 ;
        RECT 92.360 187.140 92.680 187.460 ;
        RECT 92.760 187.140 93.080 187.460 ;
        RECT 26.775 184.420 27.095 184.740 ;
        RECT 27.175 184.420 27.495 184.740 ;
        RECT 27.575 184.420 27.895 184.740 ;
        RECT 27.975 184.420 28.295 184.740 ;
        RECT 45.285 184.420 45.605 184.740 ;
        RECT 45.685 184.420 46.005 184.740 ;
        RECT 46.085 184.420 46.405 184.740 ;
        RECT 46.485 184.420 46.805 184.740 ;
        RECT 63.795 184.420 64.115 184.740 ;
        RECT 64.195 184.420 64.515 184.740 ;
        RECT 64.595 184.420 64.915 184.740 ;
        RECT 64.995 184.420 65.315 184.740 ;
        RECT 82.305 184.420 82.625 184.740 ;
        RECT 82.705 184.420 83.025 184.740 ;
        RECT 83.105 184.420 83.425 184.740 ;
        RECT 83.505 184.420 83.825 184.740 ;
        RECT 36.030 181.700 36.350 182.020 ;
        RECT 36.430 181.700 36.750 182.020 ;
        RECT 36.830 181.700 37.150 182.020 ;
        RECT 37.230 181.700 37.550 182.020 ;
        RECT 54.540 181.700 54.860 182.020 ;
        RECT 54.940 181.700 55.260 182.020 ;
        RECT 55.340 181.700 55.660 182.020 ;
        RECT 55.740 181.700 56.060 182.020 ;
        RECT 73.050 181.700 73.370 182.020 ;
        RECT 73.450 181.700 73.770 182.020 ;
        RECT 73.850 181.700 74.170 182.020 ;
        RECT 74.250 181.700 74.570 182.020 ;
        RECT 91.560 181.700 91.880 182.020 ;
        RECT 91.960 181.700 92.280 182.020 ;
        RECT 92.360 181.700 92.680 182.020 ;
        RECT 92.760 181.700 93.080 182.020 ;
        RECT 26.775 178.980 27.095 179.300 ;
        RECT 27.175 178.980 27.495 179.300 ;
        RECT 27.575 178.980 27.895 179.300 ;
        RECT 27.975 178.980 28.295 179.300 ;
        RECT 45.285 178.980 45.605 179.300 ;
        RECT 45.685 178.980 46.005 179.300 ;
        RECT 46.085 178.980 46.405 179.300 ;
        RECT 46.485 178.980 46.805 179.300 ;
        RECT 63.795 178.980 64.115 179.300 ;
        RECT 64.195 178.980 64.515 179.300 ;
        RECT 64.595 178.980 64.915 179.300 ;
        RECT 64.995 178.980 65.315 179.300 ;
        RECT 82.305 178.980 82.625 179.300 ;
        RECT 82.705 178.980 83.025 179.300 ;
        RECT 83.105 178.980 83.425 179.300 ;
        RECT 83.505 178.980 83.825 179.300 ;
        RECT 36.030 176.260 36.350 176.580 ;
        RECT 36.430 176.260 36.750 176.580 ;
        RECT 36.830 176.260 37.150 176.580 ;
        RECT 37.230 176.260 37.550 176.580 ;
        RECT 54.540 176.260 54.860 176.580 ;
        RECT 54.940 176.260 55.260 176.580 ;
        RECT 55.340 176.260 55.660 176.580 ;
        RECT 55.740 176.260 56.060 176.580 ;
        RECT 73.050 176.260 73.370 176.580 ;
        RECT 73.450 176.260 73.770 176.580 ;
        RECT 73.850 176.260 74.170 176.580 ;
        RECT 74.250 176.260 74.570 176.580 ;
        RECT 91.560 176.260 91.880 176.580 ;
        RECT 91.960 176.260 92.280 176.580 ;
        RECT 92.360 176.260 92.680 176.580 ;
        RECT 92.760 176.260 93.080 176.580 ;
        RECT 26.775 173.540 27.095 173.860 ;
        RECT 27.175 173.540 27.495 173.860 ;
        RECT 27.575 173.540 27.895 173.860 ;
        RECT 27.975 173.540 28.295 173.860 ;
        RECT 45.285 173.540 45.605 173.860 ;
        RECT 45.685 173.540 46.005 173.860 ;
        RECT 46.085 173.540 46.405 173.860 ;
        RECT 46.485 173.540 46.805 173.860 ;
        RECT 63.795 173.540 64.115 173.860 ;
        RECT 64.195 173.540 64.515 173.860 ;
        RECT 64.595 173.540 64.915 173.860 ;
        RECT 64.995 173.540 65.315 173.860 ;
        RECT 82.305 173.540 82.625 173.860 ;
        RECT 82.705 173.540 83.025 173.860 ;
        RECT 83.105 173.540 83.425 173.860 ;
        RECT 83.505 173.540 83.825 173.860 ;
        RECT 36.030 170.820 36.350 171.140 ;
        RECT 36.430 170.820 36.750 171.140 ;
        RECT 36.830 170.820 37.150 171.140 ;
        RECT 37.230 170.820 37.550 171.140 ;
        RECT 54.540 170.820 54.860 171.140 ;
        RECT 54.940 170.820 55.260 171.140 ;
        RECT 55.340 170.820 55.660 171.140 ;
        RECT 55.740 170.820 56.060 171.140 ;
        RECT 73.050 170.820 73.370 171.140 ;
        RECT 73.450 170.820 73.770 171.140 ;
        RECT 73.850 170.820 74.170 171.140 ;
        RECT 74.250 170.820 74.570 171.140 ;
        RECT 91.560 170.820 91.880 171.140 ;
        RECT 91.960 170.820 92.280 171.140 ;
        RECT 92.360 170.820 92.680 171.140 ;
        RECT 92.760 170.820 93.080 171.140 ;
        RECT 26.775 168.100 27.095 168.420 ;
        RECT 27.175 168.100 27.495 168.420 ;
        RECT 27.575 168.100 27.895 168.420 ;
        RECT 27.975 168.100 28.295 168.420 ;
        RECT 45.285 168.100 45.605 168.420 ;
        RECT 45.685 168.100 46.005 168.420 ;
        RECT 46.085 168.100 46.405 168.420 ;
        RECT 46.485 168.100 46.805 168.420 ;
        RECT 63.795 168.100 64.115 168.420 ;
        RECT 64.195 168.100 64.515 168.420 ;
        RECT 64.595 168.100 64.915 168.420 ;
        RECT 64.995 168.100 65.315 168.420 ;
        RECT 82.305 168.100 82.625 168.420 ;
        RECT 82.705 168.100 83.025 168.420 ;
        RECT 83.105 168.100 83.425 168.420 ;
        RECT 83.505 168.100 83.825 168.420 ;
        RECT 36.030 165.380 36.350 165.700 ;
        RECT 36.430 165.380 36.750 165.700 ;
        RECT 36.830 165.380 37.150 165.700 ;
        RECT 37.230 165.380 37.550 165.700 ;
        RECT 54.540 165.380 54.860 165.700 ;
        RECT 54.940 165.380 55.260 165.700 ;
        RECT 55.340 165.380 55.660 165.700 ;
        RECT 55.740 165.380 56.060 165.700 ;
        RECT 73.050 165.380 73.370 165.700 ;
        RECT 73.450 165.380 73.770 165.700 ;
        RECT 73.850 165.380 74.170 165.700 ;
        RECT 74.250 165.380 74.570 165.700 ;
        RECT 91.560 165.380 91.880 165.700 ;
        RECT 91.960 165.380 92.280 165.700 ;
        RECT 92.360 165.380 92.680 165.700 ;
        RECT 92.760 165.380 93.080 165.700 ;
        RECT 26.775 162.660 27.095 162.980 ;
        RECT 27.175 162.660 27.495 162.980 ;
        RECT 27.575 162.660 27.895 162.980 ;
        RECT 27.975 162.660 28.295 162.980 ;
        RECT 45.285 162.660 45.605 162.980 ;
        RECT 45.685 162.660 46.005 162.980 ;
        RECT 46.085 162.660 46.405 162.980 ;
        RECT 46.485 162.660 46.805 162.980 ;
        RECT 63.795 162.660 64.115 162.980 ;
        RECT 64.195 162.660 64.515 162.980 ;
        RECT 64.595 162.660 64.915 162.980 ;
        RECT 64.995 162.660 65.315 162.980 ;
        RECT 82.305 162.660 82.625 162.980 ;
        RECT 82.705 162.660 83.025 162.980 ;
        RECT 83.105 162.660 83.425 162.980 ;
        RECT 83.505 162.660 83.825 162.980 ;
        RECT 36.030 159.940 36.350 160.260 ;
        RECT 36.430 159.940 36.750 160.260 ;
        RECT 36.830 159.940 37.150 160.260 ;
        RECT 37.230 159.940 37.550 160.260 ;
        RECT 54.540 159.940 54.860 160.260 ;
        RECT 54.940 159.940 55.260 160.260 ;
        RECT 55.340 159.940 55.660 160.260 ;
        RECT 55.740 159.940 56.060 160.260 ;
        RECT 73.050 159.940 73.370 160.260 ;
        RECT 73.450 159.940 73.770 160.260 ;
        RECT 73.850 159.940 74.170 160.260 ;
        RECT 74.250 159.940 74.570 160.260 ;
        RECT 91.560 159.940 91.880 160.260 ;
        RECT 91.960 159.940 92.280 160.260 ;
        RECT 92.360 159.940 92.680 160.260 ;
        RECT 92.760 159.940 93.080 160.260 ;
        RECT 26.775 157.220 27.095 157.540 ;
        RECT 27.175 157.220 27.495 157.540 ;
        RECT 27.575 157.220 27.895 157.540 ;
        RECT 27.975 157.220 28.295 157.540 ;
        RECT 45.285 157.220 45.605 157.540 ;
        RECT 45.685 157.220 46.005 157.540 ;
        RECT 46.085 157.220 46.405 157.540 ;
        RECT 46.485 157.220 46.805 157.540 ;
        RECT 63.795 157.220 64.115 157.540 ;
        RECT 64.195 157.220 64.515 157.540 ;
        RECT 64.595 157.220 64.915 157.540 ;
        RECT 64.995 157.220 65.315 157.540 ;
        RECT 82.305 157.220 82.625 157.540 ;
        RECT 82.705 157.220 83.025 157.540 ;
        RECT 83.105 157.220 83.425 157.540 ;
        RECT 83.505 157.220 83.825 157.540 ;
        RECT 36.030 154.500 36.350 154.820 ;
        RECT 36.430 154.500 36.750 154.820 ;
        RECT 36.830 154.500 37.150 154.820 ;
        RECT 37.230 154.500 37.550 154.820 ;
        RECT 54.540 154.500 54.860 154.820 ;
        RECT 54.940 154.500 55.260 154.820 ;
        RECT 55.340 154.500 55.660 154.820 ;
        RECT 55.740 154.500 56.060 154.820 ;
        RECT 73.050 154.500 73.370 154.820 ;
        RECT 73.450 154.500 73.770 154.820 ;
        RECT 73.850 154.500 74.170 154.820 ;
        RECT 74.250 154.500 74.570 154.820 ;
        RECT 91.560 154.500 91.880 154.820 ;
        RECT 91.960 154.500 92.280 154.820 ;
        RECT 92.360 154.500 92.680 154.820 ;
        RECT 92.760 154.500 93.080 154.820 ;
        RECT 26.775 151.780 27.095 152.100 ;
        RECT 27.175 151.780 27.495 152.100 ;
        RECT 27.575 151.780 27.895 152.100 ;
        RECT 27.975 151.780 28.295 152.100 ;
        RECT 45.285 151.780 45.605 152.100 ;
        RECT 45.685 151.780 46.005 152.100 ;
        RECT 46.085 151.780 46.405 152.100 ;
        RECT 46.485 151.780 46.805 152.100 ;
        RECT 63.795 151.780 64.115 152.100 ;
        RECT 64.195 151.780 64.515 152.100 ;
        RECT 64.595 151.780 64.915 152.100 ;
        RECT 64.995 151.780 65.315 152.100 ;
        RECT 82.305 151.780 82.625 152.100 ;
        RECT 82.705 151.780 83.025 152.100 ;
        RECT 83.105 151.780 83.425 152.100 ;
        RECT 83.505 151.780 83.825 152.100 ;
        RECT 36.030 149.060 36.350 149.380 ;
        RECT 36.430 149.060 36.750 149.380 ;
        RECT 36.830 149.060 37.150 149.380 ;
        RECT 37.230 149.060 37.550 149.380 ;
        RECT 54.540 149.060 54.860 149.380 ;
        RECT 54.940 149.060 55.260 149.380 ;
        RECT 55.340 149.060 55.660 149.380 ;
        RECT 55.740 149.060 56.060 149.380 ;
        RECT 73.050 149.060 73.370 149.380 ;
        RECT 73.450 149.060 73.770 149.380 ;
        RECT 73.850 149.060 74.170 149.380 ;
        RECT 74.250 149.060 74.570 149.380 ;
        RECT 91.560 149.060 91.880 149.380 ;
        RECT 91.960 149.060 92.280 149.380 ;
        RECT 92.360 149.060 92.680 149.380 ;
        RECT 92.760 149.060 93.080 149.380 ;
        RECT 26.775 146.340 27.095 146.660 ;
        RECT 27.175 146.340 27.495 146.660 ;
        RECT 27.575 146.340 27.895 146.660 ;
        RECT 27.975 146.340 28.295 146.660 ;
        RECT 45.285 146.340 45.605 146.660 ;
        RECT 45.685 146.340 46.005 146.660 ;
        RECT 46.085 146.340 46.405 146.660 ;
        RECT 46.485 146.340 46.805 146.660 ;
        RECT 63.795 146.340 64.115 146.660 ;
        RECT 64.195 146.340 64.515 146.660 ;
        RECT 64.595 146.340 64.915 146.660 ;
        RECT 64.995 146.340 65.315 146.660 ;
        RECT 82.305 146.340 82.625 146.660 ;
        RECT 82.705 146.340 83.025 146.660 ;
        RECT 83.105 146.340 83.425 146.660 ;
        RECT 83.505 146.340 83.825 146.660 ;
        RECT 36.030 143.620 36.350 143.940 ;
        RECT 36.430 143.620 36.750 143.940 ;
        RECT 36.830 143.620 37.150 143.940 ;
        RECT 37.230 143.620 37.550 143.940 ;
        RECT 54.540 143.620 54.860 143.940 ;
        RECT 54.940 143.620 55.260 143.940 ;
        RECT 55.340 143.620 55.660 143.940 ;
        RECT 55.740 143.620 56.060 143.940 ;
        RECT 73.050 143.620 73.370 143.940 ;
        RECT 73.450 143.620 73.770 143.940 ;
        RECT 73.850 143.620 74.170 143.940 ;
        RECT 74.250 143.620 74.570 143.940 ;
        RECT 91.560 143.620 91.880 143.940 ;
        RECT 91.960 143.620 92.280 143.940 ;
        RECT 92.360 143.620 92.680 143.940 ;
        RECT 92.760 143.620 93.080 143.940 ;
        RECT 26.775 140.900 27.095 141.220 ;
        RECT 27.175 140.900 27.495 141.220 ;
        RECT 27.575 140.900 27.895 141.220 ;
        RECT 27.975 140.900 28.295 141.220 ;
        RECT 45.285 140.900 45.605 141.220 ;
        RECT 45.685 140.900 46.005 141.220 ;
        RECT 46.085 140.900 46.405 141.220 ;
        RECT 46.485 140.900 46.805 141.220 ;
        RECT 63.795 140.900 64.115 141.220 ;
        RECT 64.195 140.900 64.515 141.220 ;
        RECT 64.595 140.900 64.915 141.220 ;
        RECT 64.995 140.900 65.315 141.220 ;
        RECT 82.305 140.900 82.625 141.220 ;
        RECT 82.705 140.900 83.025 141.220 ;
        RECT 83.105 140.900 83.425 141.220 ;
        RECT 83.505 140.900 83.825 141.220 ;
        RECT 36.030 138.180 36.350 138.500 ;
        RECT 36.430 138.180 36.750 138.500 ;
        RECT 36.830 138.180 37.150 138.500 ;
        RECT 37.230 138.180 37.550 138.500 ;
        RECT 54.540 138.180 54.860 138.500 ;
        RECT 54.940 138.180 55.260 138.500 ;
        RECT 55.340 138.180 55.660 138.500 ;
        RECT 55.740 138.180 56.060 138.500 ;
        RECT 73.050 138.180 73.370 138.500 ;
        RECT 73.450 138.180 73.770 138.500 ;
        RECT 73.850 138.180 74.170 138.500 ;
        RECT 74.250 138.180 74.570 138.500 ;
        RECT 91.560 138.180 91.880 138.500 ;
        RECT 91.960 138.180 92.280 138.500 ;
        RECT 92.360 138.180 92.680 138.500 ;
        RECT 92.760 138.180 93.080 138.500 ;
        RECT 26.775 135.460 27.095 135.780 ;
        RECT 27.175 135.460 27.495 135.780 ;
        RECT 27.575 135.460 27.895 135.780 ;
        RECT 27.975 135.460 28.295 135.780 ;
        RECT 45.285 135.460 45.605 135.780 ;
        RECT 45.685 135.460 46.005 135.780 ;
        RECT 46.085 135.460 46.405 135.780 ;
        RECT 46.485 135.460 46.805 135.780 ;
        RECT 63.795 135.460 64.115 135.780 ;
        RECT 64.195 135.460 64.515 135.780 ;
        RECT 64.595 135.460 64.915 135.780 ;
        RECT 64.995 135.460 65.315 135.780 ;
        RECT 82.305 135.460 82.625 135.780 ;
        RECT 82.705 135.460 83.025 135.780 ;
        RECT 83.105 135.460 83.425 135.780 ;
        RECT 83.505 135.460 83.825 135.780 ;
        RECT 36.030 132.740 36.350 133.060 ;
        RECT 36.430 132.740 36.750 133.060 ;
        RECT 36.830 132.740 37.150 133.060 ;
        RECT 37.230 132.740 37.550 133.060 ;
        RECT 54.540 132.740 54.860 133.060 ;
        RECT 54.940 132.740 55.260 133.060 ;
        RECT 55.340 132.740 55.660 133.060 ;
        RECT 55.740 132.740 56.060 133.060 ;
        RECT 73.050 132.740 73.370 133.060 ;
        RECT 73.450 132.740 73.770 133.060 ;
        RECT 73.850 132.740 74.170 133.060 ;
        RECT 74.250 132.740 74.570 133.060 ;
        RECT 91.560 132.740 91.880 133.060 ;
        RECT 91.960 132.740 92.280 133.060 ;
        RECT 92.360 132.740 92.680 133.060 ;
        RECT 92.760 132.740 93.080 133.060 ;
        RECT 156.565 25.805 157.155 26.395 ;
      LAYER met4 ;
        RECT 26.735 136.300 28.335 206.580 ;
        RECT 26.700 132.660 28.335 136.300 ;
        RECT 35.990 135.350 37.590 206.580 ;
        RECT 45.245 136.300 46.845 206.580 ;
        RECT 35.950 132.660 37.590 135.350 ;
        RECT 45.200 132.660 46.845 136.300 ;
        RECT 54.500 135.550 56.100 206.580 ;
        RECT 63.755 137.800 65.355 206.580 ;
        RECT 54.500 132.660 56.150 135.550 ;
        RECT 63.755 132.660 65.400 137.800 ;
        RECT 73.010 135.850 74.610 206.580 ;
        RECT 0.950 124.900 1.000 126.500 ;
        RECT 2.500 124.900 2.550 126.500 ;
        RECT 26.700 124.900 28.300 132.660 ;
        RECT 35.950 121.450 37.450 132.660 ;
        RECT 45.200 124.900 46.800 132.660 ;
        RECT 54.650 121.450 56.150 132.660 ;
        RECT 63.800 124.900 65.400 132.660 ;
        RECT 72.950 132.660 74.610 135.850 ;
        RECT 82.265 138.500 83.865 206.580 ;
        RECT 82.265 132.660 83.900 138.500 ;
        RECT 91.520 132.660 93.120 206.580 ;
        RECT 72.950 121.450 74.450 132.660 ;
        RECT 82.300 124.900 83.900 132.660 ;
        RECT 9.940 119.950 93.950 121.450 ;
        RECT 156.560 1.000 157.160 26.400 ;
      LAYER via4 ;
        RECT 26.820 125.020 28.180 126.380 ;
        RECT 45.320 125.020 46.680 126.380 ;
        RECT 63.920 125.020 65.280 126.380 ;
        RECT 82.420 125.020 83.780 126.380 ;
      LAYER met5 ;
        RECT 0.830 126.500 2.670 126.620 ;
        RECT 0.830 124.900 92.700 126.500 ;
        RECT 0.830 124.780 2.670 124.900 ;
  END
END tt_um_mattvenn_r2r_dac
END LIBRARY

