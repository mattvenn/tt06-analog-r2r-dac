magic
tech sky130A
magscale 1 2
timestamp 1708001571
<< metal1 >>
rect 17138 20594 17148 20678
rect 17236 20594 17246 20678
rect 17166 20308 17210 20594
rect 17872 20578 17882 20690
rect 17996 20578 18006 20690
rect 17167 18815 17209 20308
rect 17905 19461 17947 20578
rect 18552 20576 18562 20688
rect 18676 20576 18686 20688
rect 19304 20651 19314 20694
rect 19086 20609 19314 20651
rect 17905 19419 18208 19461
rect 17167 18773 17787 18815
rect 16356 18130 16366 18360
rect 16602 18276 16612 18360
rect 17290 18276 17394 18448
rect 16602 18172 17394 18276
rect 16602 18130 16612 18172
rect 17290 18108 17394 18172
rect 17745 18155 17787 18773
rect 18166 18140 18208 19419
rect 18624 18128 18666 20576
rect 19086 18122 19128 20609
rect 19304 20582 19314 20609
rect 19428 20582 19438 20694
rect 17256 14970 17836 15140
rect 17455 12691 17621 14970
rect 18112 14204 18252 15106
rect 18584 14510 18724 15146
rect 19068 14688 19208 15158
rect 19068 14642 21200 14688
rect 19068 14562 21072 14642
rect 21162 14562 21200 14642
rect 19068 14548 21200 14562
rect 18584 14370 18944 14510
rect 18112 14064 18488 14204
rect 18584 14104 18724 14370
rect 17456 12324 17620 12691
rect 17456 12160 18272 12324
rect 18350 12290 18486 14064
rect 18806 12304 18942 14370
rect 19068 14116 19208 14548
rect 18350 12154 18740 12290
rect 18806 12168 19204 12304
<< via1 >>
rect 17148 20594 17236 20678
rect 17882 20578 17996 20690
rect 18562 20576 18676 20688
rect 16366 18130 16602 18360
rect 19314 20582 19428 20694
rect 21072 14562 21162 14642
<< metal2 >>
rect 17882 20690 17996 20700
rect 17148 20678 17236 20688
rect 17148 20584 17236 20594
rect 17882 20568 17996 20578
rect 18562 20688 18676 20698
rect 18562 20566 18676 20576
rect 19314 20694 19428 20704
rect 19314 20572 19428 20582
rect 16366 18360 16602 18370
rect 16366 18120 16602 18130
rect 21072 14642 21162 14652
rect 21072 14552 21162 14562
<< via2 >>
rect 17148 20594 17236 20678
rect 17882 20578 17996 20690
rect 18562 20576 18676 20688
rect 19314 20582 19428 20694
rect 16366 18130 16602 18360
rect 21072 14562 21162 14642
<< metal3 >>
rect 17872 20690 18006 20695
rect 19304 20694 19438 20699
rect 17138 20678 17246 20683
rect 17138 20594 17148 20678
rect 17236 20594 17246 20678
rect 17138 20589 17246 20594
rect 17872 20578 17882 20690
rect 17996 20578 18006 20690
rect 17872 20573 18006 20578
rect 18552 20688 18686 20693
rect 18552 20576 18562 20688
rect 18676 20576 18686 20688
rect 19304 20582 19314 20694
rect 19428 20582 19438 20694
rect 19304 20577 19438 20582
rect 18552 20571 18686 20576
rect 16356 18360 16612 18365
rect 16356 18130 16366 18360
rect 16602 18130 16612 18360
rect 16356 18125 16612 18130
rect 21062 14642 21172 14647
rect 21062 14562 21072 14642
rect 21162 14562 21172 14642
rect 21062 14557 21172 14562
<< via3 >>
rect 17148 20594 17236 20678
rect 17882 20578 17996 20690
rect 18562 20576 18676 20688
rect 19314 20582 19428 20694
rect 16366 18130 16602 18360
rect 21072 14562 21162 14642
<< metal4 >>
rect 200 200 500 45152
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 9800 18386 10100 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 25922 27354 45152
rect 17162 25862 27354 25922
rect 17162 20679 17222 25862
rect 28030 24710 28090 45152
rect 17912 24650 28090 24710
rect 17912 20691 17972 24650
rect 28766 23938 28826 45152
rect 18588 23878 28826 23938
rect 17881 20690 17997 20691
rect 17147 20678 17237 20679
rect 17147 20594 17148 20678
rect 17236 20594 17237 20678
rect 17147 20593 17237 20594
rect 17881 20578 17882 20690
rect 17996 20578 17997 20690
rect 18588 20689 18648 23878
rect 29502 23110 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 19334 23050 29562 23110
rect 19334 20695 19394 23050
rect 19313 20694 19429 20695
rect 17881 20577 17997 20578
rect 18561 20688 18677 20689
rect 18561 20576 18562 20688
rect 18676 20576 18677 20688
rect 19313 20582 19314 20694
rect 19428 20582 19429 20694
rect 19313 20581 19429 20582
rect 18561 20575 18677 20576
rect 9800 18360 16626 18386
rect 9800 18130 16366 18360
rect 16602 18130 16626 18360
rect 9800 18086 16626 18130
rect 200 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 9800 0 10100 18086
rect 21034 14642 31432 14660
rect 21034 14562 21072 14642
rect 21162 14562 31432 14642
rect 21034 14540 31432 14562
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31312 0 31432 14540
use sky130_fd_pr__res_generic_po_M7V662  2k
timestamp 1708000710
transform 1 0 17343 0 1 16639
box -33 -1799 33 1799
use sky130_fd_pr__res_generic_po_6GTJ3K  sky130_fd_pr__res_generic_po_6GTJ3K_0
timestamp 1708000710
transform 1 0 18185 0 1 13181
box -33 -1115 33 1115
use sky130_fd_pr__res_generic_po_6GTJ3K  sky130_fd_pr__res_generic_po_6GTJ3K_1
timestamp 1708000710
transform 1 0 18659 0 1 13211
box -33 -1115 33 1115
use sky130_fd_pr__res_generic_po_6GTJ3K  sky130_fd_pr__res_generic_po_6GTJ3K_2
timestamp 1708000710
transform 1 0 19133 0 1 13161
box -33 -1115 33 1115
use sky130_fd_pr__res_generic_po_M7V662  sky130_fd_pr__res_generic_po_M7V662_0
timestamp 1708000710
transform 1 0 17761 0 1 16631
box -33 -1799 33 1799
use sky130_fd_pr__res_generic_po_M7V662  sky130_fd_pr__res_generic_po_M7V662_1
timestamp 1708000710
transform 1 0 18185 0 1 16601
box -33 -1799 33 1799
use sky130_fd_pr__res_generic_po_M7V662  sky130_fd_pr__res_generic_po_M7V662_2
timestamp 1708000710
transform 1 0 18639 0 1 16601
box -33 -1799 33 1799
use sky130_fd_pr__res_generic_po_M7V662  sky130_fd_pr__res_generic_po_M7V662_3
timestamp 1708000710
transform 1 0 19113 0 1 16651
box -33 -1799 33 1799
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 200 0 500 45152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 0 10100 45152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
