.lib /home/matt/work/asic-workshop/shuttle-2404/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.include "../mag/tt_um_mattvenn_r2r_dac.sim.spice"

.param mc_mm_switch=1
.param mc_pr_switch=1

xtt clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6] ua[7] ui_in[4] ui_in[6] uio_in[0] uio_in[2] uio_in[3] uio_in[4] uio_in[5]
+ uio_in[6] uio_in[7] ui_in[3] ui_in[5] ui_in[7] ui_in[0] uio_in[1] ui_in[1] ui_in[2]
+ vcc 0 tt_um_mattvenn_r2r_dac_parax


* simulate tt output path
R1 "ua[0]" pin_out 500
C1 "ua[0]" 0 5p

* set ext data to be off, signal is generated inside
Vext_data uio_in[0] 0 0
Vload_div uio_in[1] 0 0

.param vcc=1.8
vcc vcc 0 {vcc}

* Digital clock signal
Vclk clk 0 PULSE {vcc} 0 0.5u 20p 20p 1u 2u

* reset signal with PULSE(V1 V2 Tdelay Trise Tfall Ton Tperiod)
* start at 0v, rise to 1.8v at 2u
Vreset rst_n 0 PULSE 0 {vcc} 2u 20p 20p 500u 1u

.control
tran 100n 40u 
write full_sim.raw
plot pin_out
.endc
.end
