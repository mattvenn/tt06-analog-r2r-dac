magic
tech sky130A
magscale 1 2
timestamp 1708461890
<< viali >>
rect 6101 15113 6135 15147
rect 8769 15113 8803 15147
rect 9965 15113 9999 15147
rect 11529 15113 11563 15147
rect 14841 15045 14875 15079
rect 8677 14977 8711 15011
rect 9873 14977 9907 15011
rect 11621 14977 11655 15011
rect 2421 14909 2455 14943
rect 3617 14909 3651 14943
rect 4905 14909 4939 14943
rect 5089 14909 5123 14943
rect 6101 14909 6135 14943
rect 6377 14909 6411 14943
rect 6469 14909 6503 14943
rect 7389 14909 7423 14943
rect 8401 14909 8435 14943
rect 9229 14909 9263 14943
rect 10149 14909 10183 14943
rect 10241 14909 10275 14943
rect 11897 14909 11931 14943
rect 11989 14909 12023 14943
rect 12541 14909 12575 14943
rect 13185 14909 13219 14943
rect 13369 14909 13403 14943
rect 13829 14909 13863 14943
rect 15025 14909 15059 14943
rect 3801 14841 3835 14875
rect 2145 14773 2179 14807
rect 2605 14773 2639 14807
rect 5825 14773 5859 14807
rect 6653 14773 6687 14807
rect 7573 14773 7607 14807
rect 8953 14773 8987 14807
rect 9045 14773 9079 14807
rect 9597 14773 9631 14807
rect 10425 14773 10459 14807
rect 11345 14773 11379 14807
rect 12173 14773 12207 14807
rect 12725 14773 12759 14807
rect 13277 14773 13311 14807
rect 14013 14773 14047 14807
rect 3525 14569 3559 14603
rect 5917 14569 5951 14603
rect 7021 14569 7055 14603
rect 8953 14569 8987 14603
rect 10977 14569 11011 14603
rect 13277 14569 13311 14603
rect 2053 14501 2087 14535
rect 3801 14501 3835 14535
rect 4528 14433 4562 14467
rect 6653 14433 6687 14467
rect 8145 14433 8179 14467
rect 8401 14433 8435 14467
rect 10077 14433 10111 14467
rect 10333 14433 10367 14467
rect 12090 14433 12124 14467
rect 12357 14433 12391 14467
rect 12791 14433 12825 14467
rect 12909 14433 12943 14467
rect 13001 14433 13035 14467
rect 13093 14433 13127 14467
rect 13369 14433 13403 14467
rect 15025 14433 15059 14467
rect 1777 14365 1811 14399
rect 4261 14365 4295 14399
rect 6285 14365 6319 14399
rect 6377 14365 6411 14399
rect 12633 14365 12667 14399
rect 13645 14365 13679 14399
rect 3985 14297 4019 14331
rect 5641 14229 5675 14263
rect 6561 14229 6595 14263
rect 6837 14229 6871 14263
rect 6745 14025 6779 14059
rect 8401 14025 8435 14059
rect 10241 14025 10275 14059
rect 11989 14025 12023 14059
rect 13185 14025 13219 14059
rect 13553 14025 13587 14059
rect 4905 13957 4939 13991
rect 9045 13889 9079 13923
rect 9597 13889 9631 13923
rect 10057 13889 10091 13923
rect 11345 13889 11379 13923
rect 11713 13889 11747 13923
rect 14749 13889 14783 13923
rect 2697 13821 2731 13855
rect 3525 13821 3559 13855
rect 3792 13821 3826 13855
rect 5549 13821 5583 13855
rect 5733 13821 5767 13855
rect 5825 13821 5859 13855
rect 6561 13821 6595 13855
rect 6837 13821 6871 13855
rect 8585 13821 8619 13855
rect 8677 13821 8711 13855
rect 9965 13821 9999 13855
rect 11805 13821 11839 13855
rect 13001 13821 13035 13855
rect 13185 13821 13219 13855
rect 13737 13821 13771 13855
rect 13829 13821 13863 13855
rect 2605 13753 2639 13787
rect 13553 13753 13587 13787
rect 6193 13685 6227 13719
rect 6285 13685 6319 13719
rect 14105 13685 14139 13719
rect 8217 13481 8251 13515
rect 8309 13481 8343 13515
rect 13185 13481 13219 13515
rect 6469 13345 6503 13379
rect 7849 13345 7883 13379
rect 8861 13345 8895 13379
rect 9873 13345 9907 13379
rect 9965 13345 9999 13379
rect 11621 13345 11655 13379
rect 12909 13345 12943 13379
rect 13277 13345 13311 13379
rect 13461 13345 13495 13379
rect 13553 13345 13587 13379
rect 13645 13345 13679 13379
rect 14013 13345 14047 13379
rect 14197 13345 14231 13379
rect 7757 13277 7791 13311
rect 8585 13277 8619 13311
rect 10333 13277 10367 13311
rect 11253 13277 11287 13311
rect 11713 13277 11747 13311
rect 13185 13277 13219 13311
rect 6561 13141 6595 13175
rect 7573 13141 7607 13175
rect 8769 13141 8803 13175
rect 9689 13141 9723 13175
rect 11897 13141 11931 13175
rect 13001 13141 13035 13175
rect 13921 13141 13955 13175
rect 14381 13141 14415 13175
rect 5549 12937 5583 12971
rect 13001 12937 13035 12971
rect 13553 12937 13587 12971
rect 6101 12869 6135 12903
rect 7941 12801 7975 12835
rect 10333 12801 10367 12835
rect 3433 12733 3467 12767
rect 5273 12733 5307 12767
rect 5825 12733 5859 12767
rect 7674 12733 7708 12767
rect 8861 12733 8895 12767
rect 12173 12733 12207 12767
rect 12725 12733 12759 12767
rect 13185 12733 13219 12767
rect 13369 12733 13403 12767
rect 13737 12733 13771 12767
rect 13921 12733 13955 12767
rect 14105 12733 14139 12767
rect 14197 12743 14231 12777
rect 14295 12733 14329 12767
rect 14473 12733 14507 12767
rect 3700 12665 3734 12699
rect 10066 12665 10100 12699
rect 11906 12665 11940 12699
rect 12541 12665 12575 12699
rect 13829 12665 13863 12699
rect 4813 12597 4847 12631
rect 5733 12597 5767 12631
rect 6285 12597 6319 12631
rect 6561 12597 6595 12631
rect 8769 12597 8803 12631
rect 8953 12597 8987 12631
rect 10793 12597 10827 12631
rect 12909 12597 12943 12631
rect 14381 12597 14415 12631
rect 9873 12393 9907 12427
rect 11161 12393 11195 12427
rect 2412 12325 2446 12359
rect 3801 12325 3835 12359
rect 6193 12325 6227 12359
rect 15025 12325 15059 12359
rect 3709 12257 3743 12291
rect 3893 12257 3927 12291
rect 4261 12257 4295 12291
rect 5917 12257 5951 12291
rect 6010 12257 6044 12291
rect 6285 12257 6319 12291
rect 6423 12257 6457 12291
rect 7205 12257 7239 12291
rect 7481 12257 7515 12291
rect 7573 12257 7607 12291
rect 9505 12257 9539 12291
rect 11713 12257 11747 12291
rect 13369 12257 13403 12291
rect 13645 12257 13679 12291
rect 2145 12189 2179 12223
rect 4905 12189 4939 12223
rect 9597 12189 9631 12223
rect 11437 12189 11471 12223
rect 3525 12121 3559 12155
rect 4353 12121 4387 12155
rect 5549 12053 5583 12087
rect 6561 12053 6595 12087
rect 7297 12053 7331 12087
rect 7757 12053 7791 12087
rect 9505 12053 9539 12087
rect 11437 12053 11471 12087
rect 2513 11849 2547 11883
rect 5641 11849 5675 11883
rect 5825 11849 5859 11883
rect 8217 11849 8251 11883
rect 8861 11849 8895 11883
rect 11897 11849 11931 11883
rect 4445 11781 4479 11815
rect 5457 11781 5491 11815
rect 8769 11781 8803 11815
rect 9229 11781 9263 11815
rect 10057 11781 10091 11815
rect 10977 11781 11011 11815
rect 3525 11713 3559 11747
rect 3801 11713 3835 11747
rect 9413 11713 9447 11747
rect 9781 11713 9815 11747
rect 2513 11645 2547 11679
rect 2697 11645 2731 11679
rect 3709 11645 3743 11679
rect 3893 11645 3927 11679
rect 3985 11645 4019 11679
rect 4169 11645 4203 11679
rect 4997 11645 5031 11679
rect 5733 11645 5767 11679
rect 6561 11645 6595 11679
rect 7573 11645 7607 11679
rect 7666 11645 7700 11679
rect 8079 11645 8113 11679
rect 8401 11645 8435 11679
rect 8677 11645 8711 11679
rect 9505 11645 9539 11679
rect 11437 11645 11471 11679
rect 12081 11645 12115 11679
rect 5181 11577 5215 11611
rect 7849 11577 7883 11611
rect 7941 11577 7975 11611
rect 9873 11577 9907 11611
rect 10425 11577 10459 11611
rect 10701 11577 10735 11611
rect 4629 11509 4663 11543
rect 4721 11509 4755 11543
rect 4813 11509 4847 11543
rect 6377 11509 6411 11543
rect 8493 11509 8527 11543
rect 9137 11509 9171 11543
rect 9965 11509 9999 11543
rect 11161 11509 11195 11543
rect 11345 11509 11379 11543
rect 11621 11509 11655 11543
rect 4169 11305 4203 11339
rect 5003 11305 5037 11339
rect 5089 11305 5123 11339
rect 10977 11305 11011 11339
rect 6276 11237 6310 11271
rect 12449 11237 12483 11271
rect 4905 11203 4939 11237
rect 2154 11169 2188 11203
rect 2421 11169 2455 11203
rect 3433 11169 3467 11203
rect 3525 11169 3559 11203
rect 3709 11169 3743 11203
rect 3801 11169 3835 11203
rect 3893 11169 3927 11203
rect 4077 11169 4111 11203
rect 4353 11169 4387 11203
rect 4804 11169 4838 11203
rect 5181 11169 5215 11203
rect 5457 11169 5491 11203
rect 8953 11169 8987 11203
rect 9229 11169 9263 11203
rect 9321 11169 9355 11203
rect 9781 11169 9815 11203
rect 9965 11169 9999 11203
rect 10057 11169 10091 11203
rect 10333 11169 10367 11203
rect 11161 11169 11195 11203
rect 11529 11169 11563 11203
rect 11989 11169 12023 11203
rect 12357 11169 12391 11203
rect 12541 11169 12575 11203
rect 12633 11169 12667 11203
rect 12726 11169 12760 11203
rect 12909 11169 12943 11203
rect 13001 11169 13035 11203
rect 13098 11169 13132 11203
rect 13369 11169 13403 11203
rect 3065 11101 3099 11135
rect 4537 11101 4571 11135
rect 4629 11101 4663 11135
rect 6009 11101 6043 11135
rect 9045 11101 9079 11135
rect 10793 11101 10827 11135
rect 11897 11101 11931 11135
rect 13645 11101 13679 11135
rect 4445 11033 4479 11067
rect 9505 11033 9539 11067
rect 9873 11033 9907 11067
rect 1041 10965 1075 10999
rect 2513 10965 2547 10999
rect 3249 10965 3283 10999
rect 3893 10965 3927 10999
rect 5365 10965 5399 10999
rect 7389 10965 7423 10999
rect 9597 10965 9631 10999
rect 10609 10965 10643 10999
rect 11161 10965 11195 10999
rect 11621 10965 11655 10999
rect 13277 10965 13311 10999
rect 14933 10965 14967 10999
rect 2329 10761 2363 10795
rect 3709 10761 3743 10795
rect 5089 10761 5123 10795
rect 6377 10761 6411 10795
rect 8125 10761 8159 10795
rect 9873 10761 9907 10795
rect 12909 10761 12943 10795
rect 13553 10761 13587 10795
rect 14289 10761 14323 10795
rect 14473 10761 14507 10795
rect 10517 10693 10551 10727
rect 11621 10693 11655 10727
rect 2605 10557 2639 10591
rect 2697 10557 2731 10591
rect 2881 10557 2915 10591
rect 4997 10557 5031 10591
rect 5273 10557 5307 10591
rect 5365 10557 5399 10591
rect 6101 10557 6135 10591
rect 6193 10557 6227 10591
rect 6469 10557 6503 10591
rect 6653 10557 6687 10591
rect 6955 10557 6989 10591
rect 7113 10557 7147 10591
rect 8217 10557 8251 10591
rect 8401 10557 8435 10591
rect 10793 10557 10827 10591
rect 10885 10557 10919 10591
rect 10977 10557 11011 10591
rect 11161 10557 11195 10591
rect 13093 10557 13127 10591
rect 13277 10557 13311 10591
rect 13369 10557 13403 10591
rect 13829 10557 13863 10591
rect 13921 10557 13955 10591
rect 14013 10557 14047 10591
rect 14197 10557 14231 10591
rect 2329 10489 2363 10523
rect 5549 10489 5583 10523
rect 5733 10489 5767 10523
rect 5917 10489 5951 10523
rect 6745 10489 6779 10523
rect 6837 10489 6871 10523
rect 11345 10489 11379 10523
rect 14657 10489 14691 10523
rect 2513 10421 2547 10455
rect 2789 10421 2823 10455
rect 14447 10421 14481 10455
rect 4353 10217 4387 10251
rect 5365 10217 5399 10251
rect 4521 10149 4555 10183
rect 4721 10149 4755 10183
rect 5273 10081 5307 10115
rect 5457 10081 5491 10115
rect 8769 10081 8803 10115
rect 8953 10081 8987 10115
rect 9045 10081 9079 10115
rect 9229 10081 9263 10115
rect 9413 10081 9447 10115
rect 11253 10081 11287 10115
rect 11345 10013 11379 10047
rect 11437 10013 11471 10047
rect 11529 10013 11563 10047
rect 8585 9945 8619 9979
rect 4537 9877 4571 9911
rect 9137 9877 9171 9911
rect 9689 9877 9723 9911
rect 11713 9877 11747 9911
rect 4905 9673 4939 9707
rect 5089 9673 5123 9707
rect 8585 9673 8619 9707
rect 9045 9673 9079 9707
rect 12541 9673 12575 9707
rect 3065 9605 3099 9639
rect 3525 9605 3559 9639
rect 5641 9605 5675 9639
rect 8769 9605 8803 9639
rect 12449 9605 12483 9639
rect 3709 9537 3743 9571
rect 8033 9537 8067 9571
rect 13093 9537 13127 9571
rect 14105 9537 14139 9571
rect 1685 9469 1719 9503
rect 3433 9469 3467 9503
rect 3617 9469 3651 9503
rect 3893 9469 3927 9503
rect 4077 9469 4111 9503
rect 5273 9469 5307 9503
rect 5457 9469 5491 9503
rect 5733 9469 5767 9503
rect 6469 9469 6503 9503
rect 6929 9469 6963 9503
rect 7113 9469 7147 9503
rect 7389 9469 7423 9503
rect 7849 9469 7883 9503
rect 7941 9469 7975 9503
rect 8125 9469 8159 9503
rect 9413 9469 9447 9503
rect 10977 9469 11011 9503
rect 11069 9469 11103 9503
rect 14381 9469 14415 9503
rect 14565 9469 14599 9503
rect 1952 9401 1986 9435
rect 4721 9401 4755 9435
rect 7021 9401 7055 9435
rect 7251 9401 7285 9435
rect 7665 9401 7699 9435
rect 8401 9401 8435 9435
rect 8861 9401 8895 9435
rect 9061 9401 9095 9435
rect 11336 9401 11370 9435
rect 13921 9401 13955 9435
rect 3249 9333 3283 9367
rect 4629 9333 4663 9367
rect 4921 9333 4955 9367
rect 5917 9333 5951 9367
rect 6285 9333 6319 9367
rect 6745 9333 6779 9367
rect 7481 9333 7515 9367
rect 8601 9333 8635 9367
rect 9229 9333 9263 9367
rect 9689 9333 9723 9367
rect 10885 9333 10919 9367
rect 13553 9333 13587 9367
rect 14013 9333 14047 9367
rect 14473 9333 14507 9367
rect 3341 9129 3375 9163
rect 3985 9129 4019 9163
rect 4905 9129 4939 9163
rect 7205 9129 7239 9163
rect 8585 9129 8619 9163
rect 10609 9129 10643 9163
rect 11713 9129 11747 9163
rect 6092 9061 6126 9095
rect 7297 9061 7331 9095
rect 9597 9061 9631 9095
rect 3249 8993 3283 9027
rect 3433 8993 3467 9027
rect 3893 8993 3927 9027
rect 4077 8993 4111 9027
rect 4813 8993 4847 9027
rect 9137 8993 9171 9027
rect 9229 8993 9263 9027
rect 9413 8993 9447 9027
rect 9689 8993 9723 9027
rect 9873 8993 9907 9027
rect 9965 8993 9999 9027
rect 10057 8993 10091 9027
rect 10425 8993 10459 9027
rect 10701 8993 10735 9027
rect 11897 8993 11931 9027
rect 12173 8993 12207 9027
rect 12357 8993 12391 9027
rect 12541 8993 12575 9027
rect 12725 8993 12759 9027
rect 13093 8993 13127 9027
rect 13277 8993 13311 9027
rect 13645 8993 13679 9027
rect 2605 8925 2639 8959
rect 5825 8925 5859 8959
rect 10977 8925 11011 8959
rect 11529 8925 11563 8959
rect 12817 8925 12851 8959
rect 12909 8925 12943 8959
rect 13369 8925 13403 8959
rect 11989 8857 12023 8891
rect 12081 8857 12115 8891
rect 1961 8789 1995 8823
rect 10333 8789 10367 8823
rect 10425 8789 10459 8823
rect 14933 8789 14967 8823
rect 2881 8585 2915 8619
rect 4445 8585 4479 8619
rect 5181 8585 5215 8619
rect 6285 8585 6319 8619
rect 11253 8585 11287 8619
rect 13185 8585 13219 8619
rect 3249 8517 3283 8551
rect 3985 8517 4019 8551
rect 4629 8517 4663 8551
rect 8677 8517 8711 8551
rect 9413 8517 9447 8551
rect 4261 8449 4295 8483
rect 6653 8449 6687 8483
rect 9873 8449 9907 8483
rect 13645 8449 13679 8483
rect 1501 8381 1535 8415
rect 3525 8381 3559 8415
rect 4537 8381 4571 8415
rect 4997 8381 5031 8415
rect 5457 8381 5491 8415
rect 6469 8381 6503 8415
rect 8585 8381 8619 8415
rect 8769 8381 8803 8415
rect 8861 8381 8895 8415
rect 9045 8381 9079 8415
rect 9137 8381 9171 8415
rect 9597 8381 9631 8415
rect 9689 8381 9723 8415
rect 10140 8381 10174 8415
rect 13185 8381 13219 8415
rect 13369 8381 13403 8415
rect 13553 8381 13587 8415
rect 13737 8381 13771 8415
rect 1768 8313 1802 8347
rect 3249 8313 3283 8347
rect 9413 8313 9447 8347
rect 3433 8245 3467 8279
rect 4813 8245 4847 8279
rect 4905 8245 4939 8279
rect 5641 8245 5675 8279
rect 8401 8245 8435 8279
rect 9229 8245 9263 8279
rect 2513 8041 2547 8075
rect 8769 8041 8803 8075
rect 4353 7973 4387 8007
rect 13185 7973 13219 8007
rect 2329 7905 2363 7939
rect 2513 7905 2547 7939
rect 4721 7905 4755 7939
rect 7389 7905 7423 7939
rect 7656 7905 7690 7939
rect 8861 7905 8895 7939
rect 9045 7905 9079 7939
rect 11989 7905 12023 7939
rect 12817 7905 12851 7939
rect 12909 7905 12943 7939
rect 13057 7905 13091 7939
rect 13277 7905 13311 7939
rect 13374 7905 13408 7939
rect 4537 7837 4571 7871
rect 4629 7837 4663 7871
rect 4813 7837 4847 7871
rect 11897 7837 11931 7871
rect 12081 7837 12115 7871
rect 12173 7837 12207 7871
rect 12725 7837 12759 7871
rect 3065 7769 3099 7803
rect 8953 7769 8987 7803
rect 12449 7769 12483 7803
rect 4997 7701 5031 7735
rect 12357 7701 12391 7735
rect 12633 7701 12667 7735
rect 13553 7701 13587 7735
rect 4353 7497 4387 7531
rect 4813 7497 4847 7531
rect 7849 7497 7883 7531
rect 11437 7497 11471 7531
rect 12173 7497 12207 7531
rect 13277 7497 13311 7531
rect 3801 7429 3835 7463
rect 6377 7429 6411 7463
rect 9689 7429 9723 7463
rect 9873 7429 9907 7463
rect 10149 7429 10183 7463
rect 4445 7361 4479 7395
rect 6837 7361 6871 7395
rect 7481 7361 7515 7395
rect 10057 7361 10091 7395
rect 12541 7361 12575 7395
rect 4629 7293 4663 7327
rect 4997 7293 5031 7327
rect 7665 7293 7699 7327
rect 7849 7293 7883 7327
rect 7941 7293 7975 7327
rect 9413 7293 9447 7327
rect 9689 7293 9723 7327
rect 9781 7293 9815 7327
rect 10425 7293 10459 7327
rect 10977 7293 11011 7327
rect 11161 7293 11195 7327
rect 11345 7293 11379 7327
rect 11437 7293 11471 7327
rect 11621 7293 11655 7327
rect 12265 7293 12299 7327
rect 12449 7293 12483 7327
rect 12633 7293 12667 7327
rect 13093 7293 13127 7327
rect 13829 7293 13863 7327
rect 13921 7293 13955 7327
rect 14013 7293 14047 7327
rect 14197 7293 14231 7327
rect 4077 7225 4111 7259
rect 5264 7225 5298 7259
rect 10057 7225 10091 7259
rect 10149 7225 10183 7259
rect 10333 7225 10367 7259
rect 11069 7225 11103 7259
rect 12909 7225 12943 7259
rect 3985 7157 4019 7191
rect 4169 7157 4203 7191
rect 8033 7157 8067 7191
rect 9505 7157 9539 7191
rect 10793 7157 10827 7191
rect 13553 7157 13587 7191
rect 2973 6953 3007 6987
rect 5365 6953 5399 6987
rect 12081 6953 12115 6987
rect 12541 6953 12575 6987
rect 12693 6885 12727 6919
rect 12909 6885 12943 6919
rect 2970 6817 3004 6851
rect 3900 6817 3934 6851
rect 4169 6817 4203 6851
rect 4353 6817 4387 6851
rect 5273 6817 5307 6851
rect 5457 6817 5491 6851
rect 6193 6817 6227 6851
rect 6377 6817 6411 6851
rect 6653 6817 6687 6851
rect 7113 6817 7147 6851
rect 11989 6817 12023 6851
rect 12265 6817 12299 6851
rect 13369 6817 13403 6851
rect 13645 6817 13679 6851
rect 15025 6817 15059 6851
rect 3433 6749 3467 6783
rect 3985 6749 4019 6783
rect 6285 6749 6319 6783
rect 6837 6749 6871 6783
rect 6929 6749 6963 6783
rect 6469 6681 6503 6715
rect 6745 6681 6779 6715
rect 12265 6681 12299 6715
rect 2789 6613 2823 6647
rect 3341 6613 3375 6647
rect 3525 6613 3559 6647
rect 4261 6613 4295 6647
rect 12725 6613 12759 6647
rect 4353 6409 4387 6443
rect 7021 6409 7055 6443
rect 9689 6409 9723 6443
rect 10977 6409 11011 6443
rect 14289 6409 14323 6443
rect 6469 6341 6503 6375
rect 8125 6341 8159 6375
rect 8493 6341 8527 6375
rect 9873 6341 9907 6375
rect 14841 6341 14875 6375
rect 1409 6273 1443 6307
rect 4169 6273 4203 6307
rect 4629 6273 4663 6307
rect 7849 6273 7883 6307
rect 11161 6273 11195 6307
rect 2881 6205 2915 6239
rect 3065 6205 3099 6239
rect 4445 6205 4479 6239
rect 4537 6205 4571 6239
rect 4721 6205 4755 6239
rect 5917 6205 5951 6239
rect 6009 6205 6043 6239
rect 6101 6205 6135 6239
rect 6193 6205 6227 6239
rect 6377 6205 6411 6239
rect 7297 6205 7331 6239
rect 7389 6205 7423 6239
rect 7757 6205 7791 6239
rect 8401 6205 8435 6239
rect 8920 6205 8954 6239
rect 9505 6205 9539 6239
rect 9781 6205 9815 6239
rect 10057 6205 10091 6239
rect 10149 6205 10183 6239
rect 10885 6205 10919 6239
rect 11253 6205 11287 6239
rect 11437 6205 11471 6239
rect 12725 6205 12759 6239
rect 13001 6205 13035 6239
rect 13185 6205 13219 6239
rect 13553 6205 13587 6239
rect 14197 6205 14231 6239
rect 14657 6205 14691 6239
rect 1676 6137 1710 6171
rect 2973 6137 3007 6171
rect 6745 6137 6779 6171
rect 9873 6137 9907 6171
rect 2789 6069 2823 6103
rect 3893 6069 3927 6103
rect 5733 6069 5767 6103
rect 6653 6069 6687 6103
rect 6837 6069 6871 6103
rect 8861 6069 8895 6103
rect 9045 6069 9079 6103
rect 9321 6069 9355 6103
rect 11161 6069 11195 6103
rect 11345 6069 11379 6103
rect 12541 6069 12575 6103
rect 14473 6069 14507 6103
rect 14565 6069 14599 6103
rect 6377 5865 6411 5899
rect 6540 5865 6574 5899
rect 7481 5865 7515 5899
rect 9137 5865 9171 5899
rect 10057 5865 10091 5899
rect 12173 5865 12207 5899
rect 3709 5797 3743 5831
rect 6745 5797 6779 5831
rect 7849 5797 7883 5831
rect 11529 5797 11563 5831
rect 3893 5729 3927 5763
rect 3985 5729 4019 5763
rect 4077 5729 4111 5763
rect 4261 5729 4295 5763
rect 4537 5729 4571 5763
rect 5089 5729 5123 5763
rect 5273 5729 5307 5763
rect 5457 5729 5491 5763
rect 6009 5729 6043 5763
rect 6193 5729 6227 5763
rect 6285 5729 6319 5763
rect 6837 5729 6871 5763
rect 7573 5729 7607 5763
rect 7757 5729 7791 5763
rect 11253 5729 11287 5763
rect 11345 5729 11379 5763
rect 12081 5729 12115 5763
rect 13093 5729 13127 5763
rect 4169 5661 4203 5695
rect 10609 5661 10643 5695
rect 12817 5661 12851 5695
rect 6009 5593 6043 5627
rect 3709 5525 3743 5559
rect 5457 5525 5491 5559
rect 6561 5525 6595 5559
rect 7757 5525 7791 5559
rect 11529 5525 11563 5559
rect 14381 5525 14415 5559
rect 4721 5321 4755 5355
rect 6377 5321 6411 5355
rect 6837 5321 6871 5355
rect 10333 5321 10367 5355
rect 12909 5321 12943 5355
rect 3341 5185 3375 5219
rect 11345 5185 11379 5219
rect 4997 5117 5031 5151
rect 5264 5117 5298 5151
rect 7950 5117 7984 5151
rect 8217 5117 8251 5151
rect 8953 5117 8987 5151
rect 11621 5117 11655 5151
rect 3608 5049 3642 5083
rect 9220 5049 9254 5083
rect 11253 4233 11287 4267
rect 9689 4097 9723 4131
rect 9965 4097 9999 4131
<< metal1 >>
rect 4982 15308 4988 15360
rect 5040 15348 5046 15360
rect 12158 15348 12164 15360
rect 5040 15320 12164 15348
rect 5040 15308 5046 15320
rect 12158 15308 12164 15320
rect 12216 15308 12222 15360
rect 552 15258 15364 15280
rect 552 15206 2249 15258
rect 2301 15206 2313 15258
rect 2365 15206 2377 15258
rect 2429 15206 2441 15258
rect 2493 15206 2505 15258
rect 2557 15206 5951 15258
rect 6003 15206 6015 15258
rect 6067 15206 6079 15258
rect 6131 15206 6143 15258
rect 6195 15206 6207 15258
rect 6259 15206 9653 15258
rect 9705 15206 9717 15258
rect 9769 15206 9781 15258
rect 9833 15206 9845 15258
rect 9897 15206 9909 15258
rect 9961 15206 13355 15258
rect 13407 15206 13419 15258
rect 13471 15206 13483 15258
rect 13535 15206 13547 15258
rect 13599 15206 13611 15258
rect 13663 15206 15364 15258
rect 552 15184 15364 15206
rect 6086 15104 6092 15156
rect 6144 15104 6150 15156
rect 6270 15104 6276 15156
rect 6328 15104 6334 15156
rect 6454 15104 6460 15156
rect 6512 15144 6518 15156
rect 8757 15147 8815 15153
rect 8757 15144 8769 15147
rect 6512 15116 8769 15144
rect 6512 15104 6518 15116
rect 8757 15113 8769 15116
rect 8803 15144 8815 15147
rect 9953 15147 10011 15153
rect 9953 15144 9965 15147
rect 8803 15116 9965 15144
rect 8803 15113 8815 15116
rect 8757 15107 8815 15113
rect 9953 15113 9965 15116
rect 9999 15144 10011 15147
rect 11422 15144 11428 15156
rect 9999 15116 11428 15144
rect 9999 15113 10011 15116
rect 9953 15107 10011 15113
rect 11422 15104 11428 15116
rect 11480 15144 11486 15156
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 11480 15116 11529 15144
rect 11480 15104 11486 15116
rect 11517 15113 11529 15116
rect 11563 15113 11575 15147
rect 11517 15107 11575 15113
rect 6288 15008 6316 15104
rect 10042 15036 10048 15088
rect 10100 15036 10106 15088
rect 11146 15036 11152 15088
rect 11204 15076 11210 15088
rect 11204 15048 12020 15076
rect 11204 15036 11210 15048
rect 8665 15011 8723 15017
rect 8665 15008 8677 15011
rect 6288 14980 6500 15008
rect 2130 14900 2136 14952
rect 2188 14940 2194 14952
rect 2409 14943 2467 14949
rect 2409 14940 2421 14943
rect 2188 14912 2421 14940
rect 2188 14900 2194 14912
rect 2409 14909 2421 14912
rect 2455 14909 2467 14943
rect 2409 14903 2467 14909
rect 3418 14900 3424 14952
rect 3476 14940 3482 14952
rect 3605 14943 3663 14949
rect 3605 14940 3617 14943
rect 3476 14912 3617 14940
rect 3476 14900 3482 14912
rect 3605 14909 3617 14912
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 4706 14900 4712 14952
rect 4764 14940 4770 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4764 14912 4905 14940
rect 4764 14900 4770 14912
rect 4893 14909 4905 14912
rect 4939 14909 4951 14943
rect 4893 14903 4951 14909
rect 5077 14943 5135 14949
rect 5077 14909 5089 14943
rect 5123 14940 5135 14943
rect 5994 14940 6000 14952
rect 5123 14912 6000 14940
rect 5123 14909 5135 14912
rect 5077 14903 5135 14909
rect 5994 14900 6000 14912
rect 6052 14900 6058 14952
rect 6089 14943 6147 14949
rect 6089 14909 6101 14943
rect 6135 14940 6147 14943
rect 6270 14940 6276 14952
rect 6135 14912 6276 14940
rect 6135 14909 6147 14912
rect 6089 14903 6147 14909
rect 6270 14900 6276 14912
rect 6328 14900 6334 14952
rect 6362 14900 6368 14952
rect 6420 14900 6426 14952
rect 6472 14949 6500 14980
rect 8496 14980 8677 15008
rect 6457 14943 6515 14949
rect 6457 14909 6469 14943
rect 6503 14909 6515 14943
rect 6457 14903 6515 14909
rect 7282 14900 7288 14952
rect 7340 14940 7346 14952
rect 7377 14943 7435 14949
rect 7377 14940 7389 14943
rect 7340 14912 7389 14940
rect 7340 14900 7346 14912
rect 7377 14909 7389 14912
rect 7423 14909 7435 14943
rect 7377 14903 7435 14909
rect 8386 14900 8392 14952
rect 8444 14900 8450 14952
rect 3789 14875 3847 14881
rect 3789 14841 3801 14875
rect 3835 14872 3847 14875
rect 4982 14872 4988 14884
rect 3835 14844 4988 14872
rect 3835 14841 3847 14844
rect 3789 14835 3847 14841
rect 4982 14832 4988 14844
rect 5040 14832 5046 14884
rect 6012 14872 6040 14900
rect 8496 14884 8524 14980
rect 8665 14977 8677 14980
rect 8711 15008 8723 15011
rect 9861 15011 9919 15017
rect 9861 15008 9873 15011
rect 8711 14980 9873 15008
rect 8711 14977 8723 14980
rect 8665 14971 8723 14977
rect 9861 14977 9873 14980
rect 9907 14977 9919 15011
rect 10060 15008 10088 15036
rect 11609 15011 11667 15017
rect 11609 15008 11621 15011
rect 10060 14980 10272 15008
rect 9861 14971 9919 14977
rect 8570 14900 8576 14952
rect 8628 14900 8634 14952
rect 9217 14943 9275 14949
rect 9217 14909 9229 14943
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 8478 14872 8484 14884
rect 5736 14844 5948 14872
rect 6012 14844 8484 14872
rect 5736 14816 5764 14844
rect 2130 14764 2136 14816
rect 2188 14764 2194 14816
rect 2590 14764 2596 14816
rect 2648 14764 2654 14816
rect 5718 14764 5724 14816
rect 5776 14764 5782 14816
rect 5810 14764 5816 14816
rect 5868 14764 5874 14816
rect 5920 14804 5948 14844
rect 8478 14832 8484 14844
rect 8536 14832 8542 14884
rect 8588 14872 8616 14900
rect 9232 14872 9260 14903
rect 8588 14844 9260 14872
rect 9876 14872 9904 14971
rect 10134 14900 10140 14952
rect 10192 14900 10198 14952
rect 10244 14949 10272 14980
rect 10336 14980 11621 15008
rect 10229 14943 10287 14949
rect 10229 14909 10241 14943
rect 10275 14909 10287 14943
rect 10229 14903 10287 14909
rect 10336 14872 10364 14980
rect 11609 14977 11621 14980
rect 11655 14977 11667 15011
rect 11609 14971 11667 14977
rect 11992 14949 12020 15048
rect 12802 15036 12808 15088
rect 12860 15076 12866 15088
rect 14829 15079 14887 15085
rect 14829 15076 14841 15079
rect 12860 15048 14841 15076
rect 12860 15036 12866 15048
rect 14829 15045 14841 15048
rect 14875 15045 14887 15079
rect 14829 15039 14887 15045
rect 11885 14943 11943 14949
rect 11885 14909 11897 14943
rect 11931 14909 11943 14943
rect 11885 14903 11943 14909
rect 11977 14943 12035 14949
rect 11977 14909 11989 14943
rect 12023 14909 12035 14943
rect 11977 14903 12035 14909
rect 9876 14844 10364 14872
rect 11900 14872 11928 14903
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 12529 14943 12587 14949
rect 12529 14940 12541 14943
rect 12492 14912 12541 14940
rect 12492 14900 12498 14912
rect 12529 14909 12541 14912
rect 12575 14909 12587 14943
rect 12529 14903 12587 14909
rect 13170 14900 13176 14952
rect 13228 14900 13234 14952
rect 13357 14943 13415 14949
rect 13357 14909 13369 14943
rect 13403 14909 13415 14943
rect 13357 14903 13415 14909
rect 13372 14872 13400 14903
rect 13722 14900 13728 14952
rect 13780 14940 13786 14952
rect 13817 14943 13875 14949
rect 13817 14940 13829 14943
rect 13780 14912 13829 14940
rect 13780 14900 13786 14912
rect 13817 14909 13829 14912
rect 13863 14909 13875 14943
rect 13817 14903 13875 14909
rect 15010 14900 15016 14952
rect 15068 14900 15074 14952
rect 11900 14844 12020 14872
rect 13372 14844 13860 14872
rect 11992 14816 12020 14844
rect 13832 14816 13860 14844
rect 6641 14807 6699 14813
rect 6641 14804 6653 14807
rect 5920 14776 6653 14804
rect 6641 14773 6653 14776
rect 6687 14773 6699 14807
rect 6641 14767 6699 14773
rect 7558 14764 7564 14816
rect 7616 14764 7622 14816
rect 8938 14764 8944 14816
rect 8996 14764 9002 14816
rect 9030 14764 9036 14816
rect 9088 14764 9094 14816
rect 9490 14764 9496 14816
rect 9548 14804 9554 14816
rect 9585 14807 9643 14813
rect 9585 14804 9597 14807
rect 9548 14776 9597 14804
rect 9548 14764 9554 14776
rect 9585 14773 9597 14776
rect 9631 14773 9643 14807
rect 9585 14767 9643 14773
rect 10410 14764 10416 14816
rect 10468 14764 10474 14816
rect 11330 14764 11336 14816
rect 11388 14764 11394 14816
rect 11974 14764 11980 14816
rect 12032 14764 12038 14816
rect 12161 14807 12219 14813
rect 12161 14773 12173 14807
rect 12207 14804 12219 14807
rect 12250 14804 12256 14816
rect 12207 14776 12256 14804
rect 12207 14773 12219 14776
rect 12161 14767 12219 14773
rect 12250 14764 12256 14776
rect 12308 14764 12314 14816
rect 12710 14764 12716 14816
rect 12768 14764 12774 14816
rect 13262 14764 13268 14816
rect 13320 14764 13326 14816
rect 13814 14764 13820 14816
rect 13872 14764 13878 14816
rect 14001 14807 14059 14813
rect 14001 14773 14013 14807
rect 14047 14804 14059 14807
rect 14182 14804 14188 14816
rect 14047 14776 14188 14804
rect 14047 14773 14059 14776
rect 14001 14767 14059 14773
rect 14182 14764 14188 14776
rect 14240 14764 14246 14816
rect 552 14714 15520 14736
rect 552 14662 4100 14714
rect 4152 14662 4164 14714
rect 4216 14662 4228 14714
rect 4280 14662 4292 14714
rect 4344 14662 4356 14714
rect 4408 14662 7802 14714
rect 7854 14662 7866 14714
rect 7918 14662 7930 14714
rect 7982 14662 7994 14714
rect 8046 14662 8058 14714
rect 8110 14662 11504 14714
rect 11556 14662 11568 14714
rect 11620 14662 11632 14714
rect 11684 14662 11696 14714
rect 11748 14662 11760 14714
rect 11812 14662 15206 14714
rect 15258 14662 15270 14714
rect 15322 14662 15334 14714
rect 15386 14662 15398 14714
rect 15450 14662 15462 14714
rect 15514 14662 15520 14714
rect 552 14640 15520 14662
rect 2130 14560 2136 14612
rect 2188 14560 2194 14612
rect 3513 14603 3571 14609
rect 3513 14569 3525 14603
rect 3559 14569 3571 14603
rect 3513 14563 3571 14569
rect 2041 14535 2099 14541
rect 2041 14501 2053 14535
rect 2087 14532 2099 14535
rect 2148 14532 2176 14560
rect 2087 14504 2176 14532
rect 2087 14501 2099 14504
rect 2041 14495 2099 14501
rect 2682 14492 2688 14544
rect 2740 14492 2746 14544
rect 3528 14532 3556 14563
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 5905 14603 5963 14609
rect 5905 14600 5917 14603
rect 5868 14572 5917 14600
rect 5868 14560 5874 14572
rect 5905 14569 5917 14572
rect 5951 14569 5963 14603
rect 5905 14563 5963 14569
rect 7009 14603 7067 14609
rect 7009 14569 7021 14603
rect 7055 14600 7067 14603
rect 7374 14600 7380 14612
rect 7055 14572 7380 14600
rect 7055 14569 7067 14572
rect 7009 14563 7067 14569
rect 7374 14560 7380 14572
rect 7432 14600 7438 14612
rect 8386 14600 8392 14612
rect 7432 14572 8392 14600
rect 7432 14560 7438 14572
rect 8386 14560 8392 14572
rect 8444 14560 8450 14612
rect 8941 14603 8999 14609
rect 8941 14569 8953 14603
rect 8987 14600 8999 14603
rect 9398 14600 9404 14612
rect 8987 14572 9404 14600
rect 8987 14569 8999 14572
rect 8941 14563 8999 14569
rect 9398 14560 9404 14572
rect 9456 14600 9462 14612
rect 10134 14600 10140 14612
rect 9456 14572 10140 14600
rect 9456 14560 9462 14572
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 10965 14603 11023 14609
rect 10965 14569 10977 14603
rect 11011 14600 11023 14603
rect 11974 14600 11980 14612
rect 11011 14572 11980 14600
rect 11011 14569 11023 14572
rect 10965 14563 11023 14569
rect 11974 14560 11980 14572
rect 12032 14560 12038 14612
rect 13170 14560 13176 14612
rect 13228 14600 13234 14612
rect 13265 14603 13323 14609
rect 13265 14600 13277 14603
rect 13228 14572 13277 14600
rect 13228 14560 13234 14572
rect 13265 14569 13277 14572
rect 13311 14569 13323 14603
rect 13265 14563 13323 14569
rect 3789 14535 3847 14541
rect 3789 14532 3801 14535
rect 3528 14504 3801 14532
rect 3789 14501 3801 14504
rect 3835 14532 3847 14535
rect 6454 14532 6460 14544
rect 3835 14504 6460 14532
rect 3835 14501 3847 14504
rect 3789 14495 3847 14501
rect 6454 14492 6460 14504
rect 6512 14492 6518 14544
rect 8404 14504 13400 14532
rect 4516 14467 4574 14473
rect 4516 14433 4528 14467
rect 4562 14464 4574 14467
rect 5534 14464 5540 14476
rect 4562 14436 5540 14464
rect 4562 14433 4574 14436
rect 4516 14427 4574 14433
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 5994 14424 6000 14476
rect 6052 14464 6058 14476
rect 6641 14467 6699 14473
rect 6641 14464 6653 14467
rect 6052 14436 6653 14464
rect 6052 14424 6058 14436
rect 6641 14433 6653 14436
rect 6687 14433 6699 14467
rect 7558 14464 7564 14476
rect 6641 14427 6699 14433
rect 7392 14436 7564 14464
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 3326 14396 3332 14408
rect 1811 14368 3332 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 3326 14356 3332 14368
rect 3384 14396 3390 14408
rect 4249 14399 4307 14405
rect 4249 14396 4261 14399
rect 3384 14368 4261 14396
rect 3384 14356 3390 14368
rect 4249 14365 4261 14368
rect 4295 14365 4307 14399
rect 4249 14359 4307 14365
rect 6270 14356 6276 14408
rect 6328 14356 6334 14408
rect 6365 14399 6423 14405
rect 6365 14365 6377 14399
rect 6411 14396 6423 14399
rect 7392 14396 7420 14436
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 8133 14467 8191 14473
rect 8133 14433 8145 14467
rect 8179 14464 8191 14467
rect 8294 14464 8300 14476
rect 8179 14436 8300 14464
rect 8179 14433 8191 14436
rect 8133 14427 8191 14433
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 8404 14473 8432 14504
rect 10336 14476 10364 14504
rect 8389 14467 8447 14473
rect 8389 14433 8401 14467
rect 8435 14433 8447 14467
rect 8389 14427 8447 14433
rect 10065 14467 10123 14473
rect 10065 14433 10077 14467
rect 10111 14464 10123 14467
rect 10226 14464 10232 14476
rect 10111 14436 10232 14464
rect 10111 14433 10123 14436
rect 10065 14427 10123 14433
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 10318 14424 10324 14476
rect 10376 14424 10382 14476
rect 12066 14424 12072 14476
rect 12124 14473 12130 14476
rect 12360 14473 12388 14504
rect 12802 14473 12808 14476
rect 12124 14427 12136 14473
rect 12345 14467 12403 14473
rect 12345 14433 12357 14467
rect 12391 14433 12403 14467
rect 12345 14427 12403 14433
rect 12779 14467 12808 14473
rect 12779 14433 12791 14467
rect 12779 14427 12808 14433
rect 12124 14424 12130 14427
rect 12802 14424 12808 14427
rect 12860 14424 12866 14476
rect 12894 14424 12900 14476
rect 12952 14424 12958 14476
rect 12986 14424 12992 14476
rect 13044 14424 13050 14476
rect 13078 14424 13084 14476
rect 13136 14424 13142 14476
rect 13372 14473 13400 14504
rect 13357 14467 13415 14473
rect 13357 14433 13369 14467
rect 13403 14433 13415 14467
rect 13357 14427 13415 14433
rect 15010 14424 15016 14476
rect 15068 14424 15074 14476
rect 6411 14368 7420 14396
rect 12621 14399 12679 14405
rect 6411 14365 6423 14368
rect 6365 14359 6423 14365
rect 12621 14365 12633 14399
rect 12667 14365 12679 14399
rect 12621 14359 12679 14365
rect 13633 14399 13691 14405
rect 13633 14365 13645 14399
rect 13679 14396 13691 14399
rect 13722 14396 13728 14408
rect 13679 14368 13728 14396
rect 13679 14365 13691 14368
rect 13633 14359 13691 14365
rect 3878 14328 3884 14340
rect 3160 14300 3884 14328
rect 3160 14272 3188 14300
rect 3878 14288 3884 14300
rect 3936 14328 3942 14340
rect 3973 14331 4031 14337
rect 3973 14328 3985 14331
rect 3936 14300 3985 14328
rect 3936 14288 3942 14300
rect 3973 14297 3985 14300
rect 4019 14297 4031 14331
rect 6288 14328 6316 14356
rect 6288 14300 6868 14328
rect 3973 14291 4031 14297
rect 3142 14220 3148 14272
rect 3200 14220 3206 14272
rect 5629 14263 5687 14269
rect 5629 14229 5641 14263
rect 5675 14260 5687 14263
rect 5810 14260 5816 14272
rect 5675 14232 5816 14260
rect 5675 14229 5687 14232
rect 5629 14223 5687 14229
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 6086 14220 6092 14272
rect 6144 14260 6150 14272
rect 6270 14260 6276 14272
rect 6144 14232 6276 14260
rect 6144 14220 6150 14232
rect 6270 14220 6276 14232
rect 6328 14220 6334 14272
rect 6546 14220 6552 14272
rect 6604 14220 6610 14272
rect 6840 14269 6868 14300
rect 6825 14263 6883 14269
rect 6825 14229 6837 14263
rect 6871 14260 6883 14263
rect 6914 14260 6920 14272
rect 6871 14232 6920 14260
rect 6871 14229 6883 14232
rect 6825 14223 6883 14229
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 12434 14220 12440 14272
rect 12492 14260 12498 14272
rect 12636 14260 12664 14359
rect 13722 14356 13728 14368
rect 13780 14356 13786 14408
rect 13998 14260 14004 14272
rect 12492 14232 14004 14260
rect 12492 14220 12498 14232
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 552 14170 15364 14192
rect 552 14118 2249 14170
rect 2301 14118 2313 14170
rect 2365 14118 2377 14170
rect 2429 14118 2441 14170
rect 2493 14118 2505 14170
rect 2557 14118 5951 14170
rect 6003 14118 6015 14170
rect 6067 14118 6079 14170
rect 6131 14118 6143 14170
rect 6195 14118 6207 14170
rect 6259 14118 9653 14170
rect 9705 14118 9717 14170
rect 9769 14118 9781 14170
rect 9833 14118 9845 14170
rect 9897 14118 9909 14170
rect 9961 14118 13355 14170
rect 13407 14118 13419 14170
rect 13471 14118 13483 14170
rect 13535 14118 13547 14170
rect 13599 14118 13611 14170
rect 13663 14118 15364 14170
rect 552 14096 15364 14118
rect 2590 14016 2596 14068
rect 2648 14016 2654 14068
rect 2682 14016 2688 14068
rect 2740 14016 2746 14068
rect 3878 14016 3884 14068
rect 3936 14056 3942 14068
rect 6270 14056 6276 14068
rect 3936 14028 6276 14056
rect 3936 14016 3942 14028
rect 6270 14016 6276 14028
rect 6328 14056 6334 14068
rect 6733 14059 6791 14065
rect 6733 14056 6745 14059
rect 6328 14028 6745 14056
rect 6328 14016 6334 14028
rect 6733 14025 6745 14028
rect 6779 14025 6791 14059
rect 6733 14019 6791 14025
rect 2608 13852 2636 14016
rect 2700 13920 2728 14016
rect 4893 13991 4951 13997
rect 4893 13957 4905 13991
rect 4939 13988 4951 13991
rect 5626 13988 5632 14000
rect 4939 13960 5632 13988
rect 4939 13957 4951 13960
rect 4893 13951 4951 13957
rect 5626 13948 5632 13960
rect 5684 13988 5690 14000
rect 6362 13988 6368 14000
rect 5684 13960 6368 13988
rect 5684 13948 5690 13960
rect 6362 13948 6368 13960
rect 6420 13948 6426 14000
rect 6546 13948 6552 14000
rect 6604 13948 6610 14000
rect 6748 13988 6776 14019
rect 8294 14016 8300 14068
rect 8352 14056 8358 14068
rect 8389 14059 8447 14065
rect 8389 14056 8401 14059
rect 8352 14028 8401 14056
rect 8352 14016 8358 14028
rect 8389 14025 8401 14028
rect 8435 14025 8447 14059
rect 8389 14019 8447 14025
rect 8570 14016 8576 14068
rect 8628 14016 8634 14068
rect 10226 14016 10232 14068
rect 10284 14016 10290 14068
rect 11977 14059 12035 14065
rect 11977 14025 11989 14059
rect 12023 14056 12035 14059
rect 12066 14056 12072 14068
rect 12023 14028 12072 14056
rect 12023 14025 12035 14028
rect 11977 14019 12035 14025
rect 12066 14016 12072 14028
rect 12124 14016 12130 14068
rect 13078 14016 13084 14068
rect 13136 14056 13142 14068
rect 13173 14059 13231 14065
rect 13173 14056 13185 14059
rect 13136 14028 13185 14056
rect 13136 14016 13142 14028
rect 13173 14025 13185 14028
rect 13219 14025 13231 14059
rect 13173 14019 13231 14025
rect 13541 14059 13599 14065
rect 13541 14025 13553 14059
rect 13587 14056 13599 14059
rect 13722 14056 13728 14068
rect 13587 14028 13728 14056
rect 13587 14025 13599 14028
rect 13541 14019 13599 14025
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 8588 13988 8616 14016
rect 12250 13988 12256 14000
rect 6748 13960 8616 13988
rect 10060 13960 12256 13988
rect 6564 13920 6592 13948
rect 6914 13920 6920 13932
rect 2700 13892 2820 13920
rect 2685 13855 2743 13861
rect 2685 13852 2697 13855
rect 2608 13824 2697 13852
rect 2685 13821 2697 13824
rect 2731 13821 2743 13855
rect 2685 13815 2743 13821
rect 2593 13787 2651 13793
rect 2593 13753 2605 13787
rect 2639 13784 2651 13787
rect 2792 13784 2820 13892
rect 5184 13892 6592 13920
rect 6748 13892 6920 13920
rect 3326 13812 3332 13864
rect 3384 13852 3390 13864
rect 3513 13855 3571 13861
rect 3513 13852 3525 13855
rect 3384 13824 3525 13852
rect 3384 13812 3390 13824
rect 3513 13821 3525 13824
rect 3559 13821 3571 13855
rect 3513 13815 3571 13821
rect 3780 13855 3838 13861
rect 3780 13821 3792 13855
rect 3826 13852 3838 13855
rect 5184 13852 5212 13892
rect 3826 13824 5212 13852
rect 3826 13821 3838 13824
rect 3780 13815 3838 13821
rect 5534 13812 5540 13864
rect 5592 13812 5598 13864
rect 5718 13812 5724 13864
rect 5776 13812 5782 13864
rect 5813 13855 5871 13861
rect 5813 13821 5825 13855
rect 5859 13852 5871 13855
rect 6549 13855 6607 13861
rect 6549 13852 6561 13855
rect 5859 13824 6561 13852
rect 5859 13821 5871 13824
rect 5813 13815 5871 13821
rect 6549 13821 6561 13824
rect 6595 13852 6607 13855
rect 6748 13852 6776 13892
rect 6914 13880 6920 13892
rect 6972 13920 6978 13932
rect 6972 13892 8708 13920
rect 6972 13880 6978 13892
rect 8680 13864 8708 13892
rect 8938 13880 8944 13932
rect 8996 13920 9002 13932
rect 9033 13923 9091 13929
rect 9033 13920 9045 13923
rect 8996 13892 9045 13920
rect 8996 13880 9002 13892
rect 9033 13889 9045 13892
rect 9079 13889 9091 13923
rect 9033 13883 9091 13889
rect 9490 13880 9496 13932
rect 9548 13920 9554 13932
rect 10060 13929 10088 13960
rect 12250 13948 12256 13960
rect 12308 13948 12314 14000
rect 9585 13923 9643 13929
rect 9585 13920 9597 13923
rect 9548 13892 9597 13920
rect 9548 13880 9554 13892
rect 9585 13889 9597 13892
rect 9631 13889 9643 13923
rect 9585 13883 9643 13889
rect 10045 13923 10103 13929
rect 10045 13889 10057 13923
rect 10091 13889 10103 13923
rect 10045 13883 10103 13889
rect 11330 13880 11336 13932
rect 11388 13880 11394 13932
rect 11701 13923 11759 13929
rect 11701 13889 11713 13923
rect 11747 13920 11759 13923
rect 12802 13920 12808 13932
rect 11747 13892 12808 13920
rect 11747 13889 11759 13892
rect 11701 13883 11759 13889
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 14737 13923 14795 13929
rect 14737 13920 14749 13923
rect 13188 13892 14749 13920
rect 6595 13824 6776 13852
rect 6825 13855 6883 13861
rect 6595 13821 6607 13824
rect 6549 13815 6607 13821
rect 6825 13821 6837 13855
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 8573 13855 8631 13861
rect 8573 13821 8585 13855
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 6840 13784 6868 13815
rect 2639 13756 2820 13784
rect 5828 13756 6868 13784
rect 8588 13784 8616 13815
rect 8662 13812 8668 13864
rect 8720 13852 8726 13864
rect 9950 13852 9956 13864
rect 8720 13824 9956 13852
rect 8720 13812 8726 13824
rect 9950 13812 9956 13824
rect 10008 13812 10014 13864
rect 10410 13812 10416 13864
rect 10468 13812 10474 13864
rect 11793 13855 11851 13861
rect 11793 13821 11805 13855
rect 11839 13852 11851 13855
rect 11882 13852 11888 13864
rect 11839 13824 11888 13852
rect 11839 13821 11851 13824
rect 11793 13815 11851 13821
rect 11882 13812 11888 13824
rect 11940 13812 11946 13864
rect 12158 13812 12164 13864
rect 12216 13852 12222 13864
rect 13188 13861 13216 13892
rect 14737 13889 14749 13892
rect 14783 13920 14795 13923
rect 15010 13920 15016 13932
rect 14783 13892 15016 13920
rect 14783 13889 14795 13892
rect 14737 13883 14795 13889
rect 15010 13880 15016 13892
rect 15068 13880 15074 13932
rect 12989 13855 13047 13861
rect 12989 13852 13001 13855
rect 12216 13824 13001 13852
rect 12216 13812 12222 13824
rect 12989 13821 13001 13824
rect 13035 13821 13047 13855
rect 12989 13815 13047 13821
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13821 13231 13855
rect 13173 13815 13231 13821
rect 13262 13812 13268 13864
rect 13320 13852 13326 13864
rect 13725 13855 13783 13861
rect 13725 13852 13737 13855
rect 13320 13824 13737 13852
rect 13320 13812 13326 13824
rect 13725 13821 13737 13824
rect 13771 13821 13783 13855
rect 13725 13815 13783 13821
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 10428 13784 10456 13812
rect 13541 13787 13599 13793
rect 13541 13784 13553 13787
rect 8588 13756 10456 13784
rect 13280 13756 13553 13784
rect 2639 13753 2651 13756
rect 2593 13747 2651 13753
rect 5828 13728 5856 13756
rect 13280 13728 13308 13756
rect 13541 13753 13553 13756
rect 13587 13753 13599 13787
rect 13541 13747 13599 13753
rect 5810 13676 5816 13728
rect 5868 13676 5874 13728
rect 6181 13719 6239 13725
rect 6181 13685 6193 13719
rect 6227 13716 6239 13719
rect 6273 13719 6331 13725
rect 6273 13716 6285 13719
rect 6227 13688 6285 13716
rect 6227 13685 6239 13688
rect 6181 13679 6239 13685
rect 6273 13685 6285 13688
rect 6319 13685 6331 13719
rect 6273 13679 6331 13685
rect 7558 13676 7564 13728
rect 7616 13716 7622 13728
rect 10502 13716 10508 13728
rect 7616 13688 10508 13716
rect 7616 13676 7622 13688
rect 10502 13676 10508 13688
rect 10560 13676 10566 13728
rect 13262 13676 13268 13728
rect 13320 13676 13326 13728
rect 13354 13676 13360 13728
rect 13412 13716 13418 13728
rect 14093 13719 14151 13725
rect 14093 13716 14105 13719
rect 13412 13688 14105 13716
rect 13412 13676 13418 13688
rect 14093 13685 14105 13688
rect 14139 13685 14151 13719
rect 14093 13679 14151 13685
rect 552 13626 15520 13648
rect 552 13574 4100 13626
rect 4152 13574 4164 13626
rect 4216 13574 4228 13626
rect 4280 13574 4292 13626
rect 4344 13574 4356 13626
rect 4408 13574 7802 13626
rect 7854 13574 7866 13626
rect 7918 13574 7930 13626
rect 7982 13574 7994 13626
rect 8046 13574 8058 13626
rect 8110 13574 11504 13626
rect 11556 13574 11568 13626
rect 11620 13574 11632 13626
rect 11684 13574 11696 13626
rect 11748 13574 11760 13626
rect 11812 13574 15206 13626
rect 15258 13574 15270 13626
rect 15322 13574 15334 13626
rect 15386 13574 15398 13626
rect 15450 13574 15462 13626
rect 15514 13574 15520 13626
rect 552 13552 15520 13574
rect 8205 13515 8263 13521
rect 8205 13481 8217 13515
rect 8251 13512 8263 13515
rect 8297 13515 8355 13521
rect 8297 13512 8309 13515
rect 8251 13484 8309 13512
rect 8251 13481 8263 13484
rect 8205 13475 8263 13481
rect 8297 13481 8309 13484
rect 8343 13481 8355 13515
rect 12710 13512 12716 13524
rect 8297 13475 8355 13481
rect 9876 13484 12716 13512
rect 6454 13336 6460 13388
rect 6512 13336 6518 13388
rect 7837 13379 7895 13385
rect 7837 13345 7849 13379
rect 7883 13376 7895 13379
rect 8662 13376 8668 13388
rect 7883 13348 8668 13376
rect 7883 13345 7895 13348
rect 7837 13339 7895 13345
rect 8662 13336 8668 13348
rect 8720 13336 8726 13388
rect 8846 13336 8852 13388
rect 8904 13336 8910 13388
rect 9876 13385 9904 13484
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 13173 13515 13231 13521
rect 13173 13481 13185 13515
rect 13219 13512 13231 13515
rect 13814 13512 13820 13524
rect 13219 13484 13820 13512
rect 13219 13481 13231 13484
rect 13173 13475 13231 13481
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 13722 13444 13728 13456
rect 13556 13416 13728 13444
rect 9861 13379 9919 13385
rect 9861 13345 9873 13379
rect 9907 13345 9919 13379
rect 9861 13339 9919 13345
rect 9950 13336 9956 13388
rect 10008 13376 10014 13388
rect 11609 13379 11667 13385
rect 11609 13376 11621 13379
rect 10008 13348 11621 13376
rect 10008 13336 10014 13348
rect 11609 13345 11621 13348
rect 11655 13376 11667 13379
rect 11882 13376 11888 13388
rect 11655 13348 11888 13376
rect 11655 13345 11667 13348
rect 11609 13339 11667 13345
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 12618 13336 12624 13388
rect 12676 13376 12682 13388
rect 13556 13385 13584 13416
rect 13722 13404 13728 13416
rect 13780 13404 13786 13456
rect 13924 13416 14504 13444
rect 12897 13379 12955 13385
rect 12897 13376 12909 13379
rect 12676 13348 12909 13376
rect 12676 13336 12682 13348
rect 12897 13345 12909 13348
rect 12943 13345 12955 13379
rect 13265 13379 13323 13385
rect 13265 13376 13277 13379
rect 12897 13339 12955 13345
rect 13004 13348 13277 13376
rect 7745 13311 7803 13317
rect 7745 13277 7757 13311
rect 7791 13277 7803 13311
rect 7745 13271 7803 13277
rect 7760 13240 7788 13271
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 8573 13311 8631 13317
rect 8573 13308 8585 13311
rect 8536 13280 8585 13308
rect 8536 13268 8542 13280
rect 8573 13277 8585 13280
rect 8619 13277 8631 13311
rect 8573 13271 8631 13277
rect 10134 13268 10140 13320
rect 10192 13308 10198 13320
rect 10321 13311 10379 13317
rect 10321 13308 10333 13311
rect 10192 13280 10333 13308
rect 10192 13268 10198 13280
rect 10321 13277 10333 13280
rect 10367 13277 10379 13311
rect 10321 13271 10379 13277
rect 11238 13268 11244 13320
rect 11296 13268 11302 13320
rect 11701 13311 11759 13317
rect 11701 13277 11713 13311
rect 11747 13277 11759 13311
rect 11701 13271 11759 13277
rect 9030 13240 9036 13252
rect 7760 13212 9036 13240
rect 8588 13184 8616 13212
rect 9030 13200 9036 13212
rect 9088 13200 9094 13252
rect 11716 13240 11744 13271
rect 12342 13268 12348 13320
rect 12400 13308 12406 13320
rect 13004 13308 13032 13348
rect 13265 13345 13277 13348
rect 13311 13345 13323 13379
rect 13265 13339 13323 13345
rect 13449 13379 13507 13385
rect 13449 13345 13461 13379
rect 13495 13345 13507 13379
rect 13449 13339 13507 13345
rect 13541 13379 13599 13385
rect 13541 13345 13553 13379
rect 13587 13345 13599 13379
rect 13541 13339 13599 13345
rect 13633 13379 13691 13385
rect 13633 13345 13645 13379
rect 13679 13376 13691 13379
rect 13924 13376 13952 13416
rect 14476 13388 14504 13416
rect 13679 13348 13952 13376
rect 13679 13345 13691 13348
rect 13633 13339 13691 13345
rect 12400 13280 13032 13308
rect 13173 13311 13231 13317
rect 12400 13268 12406 13280
rect 13173 13277 13185 13311
rect 13219 13308 13231 13311
rect 13354 13308 13360 13320
rect 13219 13280 13360 13308
rect 13219 13277 13231 13280
rect 13173 13271 13231 13277
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 13464 13308 13492 13339
rect 13998 13336 14004 13388
rect 14056 13336 14062 13388
rect 14182 13336 14188 13388
rect 14240 13336 14246 13388
rect 14458 13336 14464 13388
rect 14516 13336 14522 13388
rect 13722 13308 13728 13320
rect 13464 13280 13728 13308
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 14200 13240 14228 13336
rect 11716 13212 14228 13240
rect 6454 13132 6460 13184
rect 6512 13172 6518 13184
rect 6549 13175 6607 13181
rect 6549 13172 6561 13175
rect 6512 13144 6561 13172
rect 6512 13132 6518 13144
rect 6549 13141 6561 13144
rect 6595 13141 6607 13175
rect 6549 13135 6607 13141
rect 7561 13175 7619 13181
rect 7561 13141 7573 13175
rect 7607 13172 7619 13175
rect 7650 13172 7656 13184
rect 7607 13144 7656 13172
rect 7607 13141 7619 13144
rect 7561 13135 7619 13141
rect 7650 13132 7656 13144
rect 7708 13132 7714 13184
rect 8570 13132 8576 13184
rect 8628 13132 8634 13184
rect 8662 13132 8668 13184
rect 8720 13172 8726 13184
rect 8757 13175 8815 13181
rect 8757 13172 8769 13175
rect 8720 13144 8769 13172
rect 8720 13132 8726 13144
rect 8757 13141 8769 13144
rect 8803 13172 8815 13175
rect 9490 13172 9496 13184
rect 8803 13144 9496 13172
rect 8803 13141 8815 13144
rect 8757 13135 8815 13141
rect 9490 13132 9496 13144
rect 9548 13132 9554 13184
rect 9677 13175 9735 13181
rect 9677 13141 9689 13175
rect 9723 13172 9735 13175
rect 10042 13172 10048 13184
rect 9723 13144 10048 13172
rect 9723 13141 9735 13144
rect 9677 13135 9735 13141
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 11882 13132 11888 13184
rect 11940 13132 11946 13184
rect 12986 13132 12992 13184
rect 13044 13132 13050 13184
rect 13906 13132 13912 13184
rect 13964 13132 13970 13184
rect 14182 13132 14188 13184
rect 14240 13172 14246 13184
rect 14369 13175 14427 13181
rect 14369 13172 14381 13175
rect 14240 13144 14381 13172
rect 14240 13132 14246 13144
rect 14369 13141 14381 13144
rect 14415 13141 14427 13175
rect 14369 13135 14427 13141
rect 552 13082 15364 13104
rect 552 13030 2249 13082
rect 2301 13030 2313 13082
rect 2365 13030 2377 13082
rect 2429 13030 2441 13082
rect 2493 13030 2505 13082
rect 2557 13030 5951 13082
rect 6003 13030 6015 13082
rect 6067 13030 6079 13082
rect 6131 13030 6143 13082
rect 6195 13030 6207 13082
rect 6259 13030 9653 13082
rect 9705 13030 9717 13082
rect 9769 13030 9781 13082
rect 9833 13030 9845 13082
rect 9897 13030 9909 13082
rect 9961 13030 13355 13082
rect 13407 13030 13419 13082
rect 13471 13030 13483 13082
rect 13535 13030 13547 13082
rect 13599 13030 13611 13082
rect 13663 13030 15364 13082
rect 552 13008 15364 13030
rect 5537 12971 5595 12977
rect 5537 12937 5549 12971
rect 5583 12968 5595 12971
rect 5626 12968 5632 12980
rect 5583 12940 5632 12968
rect 5583 12937 5595 12940
rect 5537 12931 5595 12937
rect 5626 12928 5632 12940
rect 5684 12928 5690 12980
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 5776 12940 9352 12968
rect 5776 12928 5782 12940
rect 5644 12900 5672 12928
rect 9324 12912 9352 12940
rect 12986 12928 12992 12980
rect 13044 12928 13050 12980
rect 13541 12971 13599 12977
rect 13541 12937 13553 12971
rect 13587 12968 13599 12971
rect 13722 12968 13728 12980
rect 13587 12940 13728 12968
rect 13587 12937 13599 12940
rect 13541 12931 13599 12937
rect 13722 12928 13728 12940
rect 13780 12928 13786 12980
rect 6089 12903 6147 12909
rect 6089 12900 6101 12903
rect 5644 12872 6101 12900
rect 6089 12869 6101 12872
rect 6135 12869 6147 12903
rect 6089 12863 6147 12869
rect 9306 12860 9312 12912
rect 9364 12860 9370 12912
rect 12618 12860 12624 12912
rect 12676 12900 12682 12912
rect 12676 12872 14044 12900
rect 12676 12860 12682 12872
rect 7929 12835 7987 12841
rect 7929 12801 7941 12835
rect 7975 12832 7987 12835
rect 7975 12804 9352 12832
rect 7975 12801 7987 12804
rect 7929 12795 7987 12801
rect 3326 12724 3332 12776
rect 3384 12764 3390 12776
rect 3421 12767 3479 12773
rect 3421 12764 3433 12767
rect 3384 12736 3433 12764
rect 3384 12724 3390 12736
rect 3421 12733 3433 12736
rect 3467 12733 3479 12767
rect 5261 12767 5319 12773
rect 5261 12764 5273 12767
rect 3421 12727 3479 12733
rect 4816 12736 5273 12764
rect 3688 12699 3746 12705
rect 3688 12665 3700 12699
rect 3734 12696 3746 12699
rect 3786 12696 3792 12708
rect 3734 12668 3792 12696
rect 3734 12665 3746 12668
rect 3688 12659 3746 12665
rect 3786 12656 3792 12668
rect 3844 12656 3850 12708
rect 4706 12588 4712 12640
rect 4764 12628 4770 12640
rect 4816 12637 4844 12736
rect 5261 12733 5273 12736
rect 5307 12764 5319 12767
rect 5813 12767 5871 12773
rect 5813 12764 5825 12767
rect 5307 12736 5825 12764
rect 5307 12733 5319 12736
rect 5261 12727 5319 12733
rect 5813 12733 5825 12736
rect 5859 12733 5871 12767
rect 5813 12727 5871 12733
rect 7650 12724 7656 12776
rect 7708 12773 7714 12776
rect 7708 12764 7720 12773
rect 8849 12767 8907 12773
rect 7708 12736 7753 12764
rect 7708 12727 7720 12736
rect 8849 12733 8861 12767
rect 8895 12764 8907 12767
rect 9324 12764 9352 12804
rect 10318 12792 10324 12844
rect 10376 12792 10382 12844
rect 13372 12804 13952 12832
rect 10336 12764 10364 12792
rect 12158 12764 12164 12776
rect 8895 12736 8984 12764
rect 9324 12736 12164 12764
rect 8895 12733 8907 12736
rect 8849 12727 8907 12733
rect 7708 12724 7714 12727
rect 4801 12631 4859 12637
rect 4801 12628 4813 12631
rect 4764 12600 4813 12628
rect 4764 12588 4770 12600
rect 4801 12597 4813 12600
rect 4847 12597 4859 12631
rect 4801 12591 4859 12597
rect 5718 12588 5724 12640
rect 5776 12588 5782 12640
rect 5902 12588 5908 12640
rect 5960 12628 5966 12640
rect 6273 12631 6331 12637
rect 6273 12628 6285 12631
rect 5960 12600 6285 12628
rect 5960 12588 5966 12600
rect 6273 12597 6285 12600
rect 6319 12597 6331 12631
rect 6273 12591 6331 12597
rect 6549 12631 6607 12637
rect 6549 12597 6561 12631
rect 6595 12628 6607 12631
rect 7558 12628 7564 12640
rect 6595 12600 7564 12628
rect 6595 12597 6607 12600
rect 6549 12591 6607 12597
rect 7558 12588 7564 12600
rect 7616 12588 7622 12640
rect 8754 12588 8760 12640
rect 8812 12588 8818 12640
rect 8956 12637 8984 12736
rect 12158 12724 12164 12736
rect 12216 12724 12222 12776
rect 12713 12767 12771 12773
rect 12713 12733 12725 12767
rect 12759 12764 12771 12767
rect 12986 12764 12992 12776
rect 12759 12736 12992 12764
rect 12759 12733 12771 12736
rect 12713 12727 12771 12733
rect 12986 12724 12992 12736
rect 13044 12724 13050 12776
rect 13372 12773 13400 12804
rect 13173 12767 13231 12773
rect 13173 12733 13185 12767
rect 13219 12733 13231 12767
rect 13173 12727 13231 12733
rect 13357 12767 13415 12773
rect 13357 12733 13369 12767
rect 13403 12733 13415 12767
rect 13357 12727 13415 12733
rect 10042 12656 10048 12708
rect 10100 12705 10106 12708
rect 10100 12696 10112 12705
rect 10100 12668 10145 12696
rect 10100 12659 10112 12668
rect 10100 12656 10106 12659
rect 11882 12656 11888 12708
rect 11940 12705 11946 12708
rect 11940 12696 11952 12705
rect 12529 12699 12587 12705
rect 11940 12668 11985 12696
rect 11940 12659 11952 12668
rect 12529 12665 12541 12699
rect 12575 12696 12587 12699
rect 13078 12696 13084 12708
rect 12575 12668 13084 12696
rect 12575 12665 12587 12668
rect 12529 12659 12587 12665
rect 11940 12656 11946 12659
rect 13078 12656 13084 12668
rect 13136 12656 13142 12708
rect 13188 12696 13216 12727
rect 13722 12724 13728 12776
rect 13780 12724 13786 12776
rect 13924 12773 13952 12804
rect 13909 12767 13967 12773
rect 13909 12733 13921 12767
rect 13955 12733 13967 12767
rect 14016 12764 14044 12872
rect 14093 12767 14151 12773
rect 14093 12764 14105 12767
rect 14016 12736 14105 12764
rect 13909 12727 13967 12733
rect 14093 12733 14105 12736
rect 14139 12733 14151 12767
rect 14182 12734 14188 12786
rect 14240 12734 14246 12786
rect 14093 12727 14151 12733
rect 13446 12696 13452 12708
rect 13188 12668 13452 12696
rect 13446 12656 13452 12668
rect 13504 12656 13510 12708
rect 13817 12699 13875 12705
rect 13817 12665 13829 12699
rect 13863 12665 13875 12699
rect 13924 12696 13952 12727
rect 14274 12724 14280 12776
rect 14332 12773 14338 12776
rect 14332 12764 14341 12773
rect 14332 12736 14377 12764
rect 14332 12727 14341 12736
rect 14332 12724 14338 12727
rect 14458 12724 14464 12776
rect 14516 12764 14522 12776
rect 14516 12736 15056 12764
rect 14516 12724 14522 12736
rect 15028 12708 15056 12736
rect 13924 12668 14504 12696
rect 13817 12659 13875 12665
rect 8941 12631 8999 12637
rect 8941 12597 8953 12631
rect 8987 12628 8999 12631
rect 9030 12628 9036 12640
rect 8987 12600 9036 12628
rect 8987 12597 8999 12600
rect 8941 12591 8999 12597
rect 9030 12588 9036 12600
rect 9088 12588 9094 12640
rect 10594 12588 10600 12640
rect 10652 12628 10658 12640
rect 10781 12631 10839 12637
rect 10781 12628 10793 12631
rect 10652 12600 10793 12628
rect 10652 12588 10658 12600
rect 10781 12597 10793 12600
rect 10827 12597 10839 12631
rect 10781 12591 10839 12597
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13538 12628 13544 12640
rect 12943 12600 13544 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13538 12588 13544 12600
rect 13596 12588 13602 12640
rect 13832 12628 13860 12659
rect 14476 12640 14504 12668
rect 15010 12656 15016 12708
rect 15068 12656 15074 12708
rect 13998 12628 14004 12640
rect 13832 12600 14004 12628
rect 13998 12588 14004 12600
rect 14056 12628 14062 12640
rect 14369 12631 14427 12637
rect 14369 12628 14381 12631
rect 14056 12600 14381 12628
rect 14056 12588 14062 12600
rect 14369 12597 14381 12600
rect 14415 12597 14427 12631
rect 14369 12591 14427 12597
rect 14458 12588 14464 12640
rect 14516 12588 14522 12640
rect 552 12538 15520 12560
rect 552 12486 4100 12538
rect 4152 12486 4164 12538
rect 4216 12486 4228 12538
rect 4280 12486 4292 12538
rect 4344 12486 4356 12538
rect 4408 12486 7802 12538
rect 7854 12486 7866 12538
rect 7918 12486 7930 12538
rect 7982 12486 7994 12538
rect 8046 12486 8058 12538
rect 8110 12486 11504 12538
rect 11556 12486 11568 12538
rect 11620 12486 11632 12538
rect 11684 12486 11696 12538
rect 11748 12486 11760 12538
rect 11812 12486 15206 12538
rect 15258 12486 15270 12538
rect 15322 12486 15334 12538
rect 15386 12486 15398 12538
rect 15450 12486 15462 12538
rect 15514 12486 15520 12538
rect 552 12464 15520 12486
rect 842 12384 848 12436
rect 900 12424 906 12436
rect 7282 12424 7288 12436
rect 900 12396 7288 12424
rect 900 12384 906 12396
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 9861 12427 9919 12433
rect 9861 12393 9873 12427
rect 9907 12424 9919 12427
rect 10134 12424 10140 12436
rect 9907 12396 10140 12424
rect 9907 12393 9919 12396
rect 9861 12387 9919 12393
rect 10134 12384 10140 12396
rect 10192 12384 10198 12436
rect 11149 12427 11207 12433
rect 11149 12393 11161 12427
rect 11195 12424 11207 12427
rect 11238 12424 11244 12436
rect 11195 12396 11244 12424
rect 11195 12393 11207 12396
rect 11149 12387 11207 12393
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 13078 12384 13084 12436
rect 13136 12424 13142 12436
rect 14274 12424 14280 12436
rect 13136 12396 14280 12424
rect 13136 12384 13142 12396
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 2400 12359 2458 12365
rect 2400 12325 2412 12359
rect 2446 12356 2458 12359
rect 2590 12356 2596 12368
rect 2446 12328 2596 12356
rect 2446 12325 2458 12328
rect 2400 12319 2458 12325
rect 2590 12316 2596 12328
rect 2648 12316 2654 12368
rect 3786 12316 3792 12368
rect 3844 12316 3850 12368
rect 5718 12316 5724 12368
rect 5776 12356 5782 12368
rect 6181 12359 6239 12365
rect 6181 12356 6193 12359
rect 5776 12328 6193 12356
rect 5776 12316 5782 12328
rect 6181 12325 6193 12328
rect 6227 12325 6239 12359
rect 6181 12319 6239 12325
rect 7116 12328 7604 12356
rect 3602 12248 3608 12300
rect 3660 12288 3666 12300
rect 3697 12291 3755 12297
rect 3697 12288 3709 12291
rect 3660 12260 3709 12288
rect 3660 12248 3666 12260
rect 3697 12257 3709 12260
rect 3743 12257 3755 12291
rect 3697 12251 3755 12257
rect 3878 12248 3884 12300
rect 3936 12248 3942 12300
rect 4249 12291 4307 12297
rect 4249 12257 4261 12291
rect 4295 12257 4307 12291
rect 4249 12251 4307 12257
rect 2130 12180 2136 12232
rect 2188 12180 2194 12232
rect 4264 12220 4292 12251
rect 5902 12248 5908 12300
rect 5960 12248 5966 12300
rect 5998 12291 6056 12297
rect 5998 12257 6010 12291
rect 6044 12257 6056 12291
rect 5998 12251 6056 12257
rect 3528 12192 4292 12220
rect 3528 12164 3556 12192
rect 4706 12180 4712 12232
rect 4764 12220 4770 12232
rect 4893 12223 4951 12229
rect 4893 12220 4905 12223
rect 4764 12192 4905 12220
rect 4764 12180 4770 12192
rect 4893 12189 4905 12192
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 6012 12220 6040 12251
rect 6270 12248 6276 12300
rect 6328 12248 6334 12300
rect 6411 12291 6469 12297
rect 6411 12257 6423 12291
rect 6457 12288 6469 12291
rect 7116 12288 7144 12328
rect 7576 12300 7604 12328
rect 15010 12316 15016 12368
rect 15068 12316 15074 12368
rect 6457 12260 7144 12288
rect 7193 12291 7251 12297
rect 6457 12257 6469 12260
rect 6411 12251 6469 12257
rect 7193 12257 7205 12291
rect 7239 12257 7251 12291
rect 7193 12251 7251 12257
rect 5684 12192 6040 12220
rect 5684 12180 5690 12192
rect 3510 12112 3516 12164
rect 3568 12112 3574 12164
rect 4338 12112 4344 12164
rect 4396 12152 4402 12164
rect 7208 12152 7236 12251
rect 7466 12248 7472 12300
rect 7524 12248 7530 12300
rect 7558 12248 7564 12300
rect 7616 12288 7622 12300
rect 8846 12288 8852 12300
rect 7616 12260 8852 12288
rect 7616 12248 7622 12260
rect 8846 12248 8852 12260
rect 8904 12248 8910 12300
rect 9490 12248 9496 12300
rect 9548 12288 9554 12300
rect 10226 12288 10232 12300
rect 9548 12260 10232 12288
rect 9548 12248 9554 12260
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 10594 12248 10600 12300
rect 10652 12288 10658 12300
rect 11701 12291 11759 12297
rect 11701 12288 11713 12291
rect 10652 12260 11713 12288
rect 10652 12248 10658 12260
rect 11701 12257 11713 12260
rect 11747 12257 11759 12291
rect 11701 12251 11759 12257
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 13262 12288 13268 12300
rect 12216 12260 13268 12288
rect 12216 12248 12222 12260
rect 13262 12248 13268 12260
rect 13320 12288 13326 12300
rect 13357 12291 13415 12297
rect 13357 12288 13369 12291
rect 13320 12260 13369 12288
rect 13320 12248 13326 12260
rect 13357 12257 13369 12260
rect 13403 12257 13415 12291
rect 13357 12251 13415 12257
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 13906 12288 13912 12300
rect 13679 12260 13912 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 13906 12248 13912 12260
rect 13964 12248 13970 12300
rect 8478 12180 8484 12232
rect 8536 12220 8542 12232
rect 9585 12223 9643 12229
rect 9585 12220 9597 12223
rect 8536 12192 9597 12220
rect 8536 12180 8542 12192
rect 9585 12189 9597 12192
rect 9631 12220 9643 12223
rect 11425 12223 11483 12229
rect 11425 12220 11437 12223
rect 9631 12192 11437 12220
rect 9631 12189 9643 12192
rect 9585 12183 9643 12189
rect 11425 12189 11437 12192
rect 11471 12189 11483 12223
rect 11425 12183 11483 12189
rect 14090 12180 14096 12232
rect 14148 12220 14154 12232
rect 14458 12220 14464 12232
rect 14148 12192 14464 12220
rect 14148 12180 14154 12192
rect 14458 12180 14464 12192
rect 14516 12180 14522 12232
rect 7650 12152 7656 12164
rect 4396 12124 7656 12152
rect 4396 12112 4402 12124
rect 7650 12112 7656 12124
rect 7708 12112 7714 12164
rect 8110 12112 8116 12164
rect 8168 12152 8174 12164
rect 9398 12152 9404 12164
rect 8168 12124 9404 12152
rect 8168 12112 8174 12124
rect 9398 12112 9404 12124
rect 9456 12112 9462 12164
rect 5534 12044 5540 12096
rect 5592 12044 5598 12096
rect 6549 12087 6607 12093
rect 6549 12053 6561 12087
rect 6595 12084 6607 12087
rect 7190 12084 7196 12096
rect 6595 12056 7196 12084
rect 6595 12053 6607 12056
rect 6549 12047 6607 12053
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 7285 12087 7343 12093
rect 7285 12053 7297 12087
rect 7331 12084 7343 12087
rect 7374 12084 7380 12096
rect 7331 12056 7380 12084
rect 7331 12053 7343 12056
rect 7285 12047 7343 12053
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 7745 12087 7803 12093
rect 7745 12053 7757 12087
rect 7791 12084 7803 12087
rect 8202 12084 8208 12096
rect 7791 12056 8208 12084
rect 7791 12053 7803 12056
rect 7745 12047 7803 12053
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 8754 12044 8760 12096
rect 8812 12084 8818 12096
rect 9490 12084 9496 12096
rect 8812 12056 9496 12084
rect 8812 12044 8818 12056
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 11422 12044 11428 12096
rect 11480 12044 11486 12096
rect 552 11994 15364 12016
rect 552 11942 2249 11994
rect 2301 11942 2313 11994
rect 2365 11942 2377 11994
rect 2429 11942 2441 11994
rect 2493 11942 2505 11994
rect 2557 11942 5951 11994
rect 6003 11942 6015 11994
rect 6067 11942 6079 11994
rect 6131 11942 6143 11994
rect 6195 11942 6207 11994
rect 6259 11942 9653 11994
rect 9705 11942 9717 11994
rect 9769 11942 9781 11994
rect 9833 11942 9845 11994
rect 9897 11942 9909 11994
rect 9961 11942 13355 11994
rect 13407 11942 13419 11994
rect 13471 11942 13483 11994
rect 13535 11942 13547 11994
rect 13599 11942 13611 11994
rect 13663 11942 15364 11994
rect 552 11920 15364 11942
rect 2501 11883 2559 11889
rect 2501 11849 2513 11883
rect 2547 11880 2559 11883
rect 2590 11880 2596 11892
rect 2547 11852 2596 11880
rect 2547 11849 2559 11852
rect 2501 11843 2559 11849
rect 2590 11840 2596 11852
rect 2648 11840 2654 11892
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 3568 11852 4476 11880
rect 3568 11840 3574 11852
rect 3694 11772 3700 11824
rect 3752 11812 3758 11824
rect 3970 11812 3976 11824
rect 3752 11784 3976 11812
rect 3752 11772 3758 11784
rect 3970 11772 3976 11784
rect 4028 11772 4034 11824
rect 4448 11821 4476 11852
rect 5626 11840 5632 11892
rect 5684 11840 5690 11892
rect 5813 11883 5871 11889
rect 5813 11849 5825 11883
rect 5859 11880 5871 11883
rect 6270 11880 6276 11892
rect 5859 11852 6276 11880
rect 5859 11849 5871 11852
rect 5813 11843 5871 11849
rect 6270 11840 6276 11852
rect 6328 11880 6334 11892
rect 7466 11880 7472 11892
rect 6328 11852 7472 11880
rect 6328 11840 6334 11852
rect 7466 11840 7472 11852
rect 7524 11840 7530 11892
rect 8205 11883 8263 11889
rect 8205 11849 8217 11883
rect 8251 11880 8263 11883
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 8251 11852 8861 11880
rect 8251 11849 8263 11852
rect 8205 11843 8263 11849
rect 8849 11849 8861 11852
rect 8895 11849 8907 11883
rect 8849 11843 8907 11849
rect 9030 11840 9036 11892
rect 9088 11880 9094 11892
rect 9088 11852 9352 11880
rect 9088 11840 9094 11852
rect 4433 11815 4491 11821
rect 4433 11781 4445 11815
rect 4479 11812 4491 11815
rect 4890 11812 4896 11824
rect 4479 11784 4896 11812
rect 4479 11781 4491 11784
rect 4433 11775 4491 11781
rect 4890 11772 4896 11784
rect 4948 11772 4954 11824
rect 5445 11815 5503 11821
rect 5445 11781 5457 11815
rect 5491 11812 5503 11815
rect 5718 11812 5724 11824
rect 5491 11784 5724 11812
rect 5491 11781 5503 11784
rect 5445 11775 5503 11781
rect 5718 11772 5724 11784
rect 5776 11772 5782 11824
rect 8757 11815 8815 11821
rect 8757 11781 8769 11815
rect 8803 11812 8815 11815
rect 9217 11815 9275 11821
rect 9217 11812 9229 11815
rect 8803 11784 9229 11812
rect 8803 11781 8815 11784
rect 8757 11775 8815 11781
rect 9217 11781 9229 11784
rect 9263 11781 9275 11815
rect 9324 11812 9352 11852
rect 11882 11840 11888 11892
rect 11940 11840 11946 11892
rect 12066 11840 12072 11892
rect 12124 11840 12130 11892
rect 10045 11815 10103 11821
rect 10045 11812 10057 11815
rect 9324 11784 10057 11812
rect 9217 11775 9275 11781
rect 10045 11781 10057 11784
rect 10091 11781 10103 11815
rect 10045 11775 10103 11781
rect 10594 11772 10600 11824
rect 10652 11812 10658 11824
rect 10965 11815 11023 11821
rect 10965 11812 10977 11815
rect 10652 11784 10977 11812
rect 10652 11772 10658 11784
rect 10965 11781 10977 11784
rect 11011 11781 11023 11815
rect 10965 11775 11023 11781
rect 3513 11747 3571 11753
rect 3513 11744 3525 11747
rect 2516 11716 3525 11744
rect 2516 11685 2544 11716
rect 3513 11713 3525 11716
rect 3559 11713 3571 11747
rect 3513 11707 3571 11713
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11744 3847 11747
rect 4062 11744 4068 11756
rect 3835 11716 4068 11744
rect 3835 11713 3847 11716
rect 3789 11707 3847 11713
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 7576 11716 9168 11744
rect 2501 11679 2559 11685
rect 2501 11645 2513 11679
rect 2547 11645 2559 11679
rect 2501 11639 2559 11645
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11676 2743 11679
rect 3602 11676 3608 11688
rect 2731 11648 3608 11676
rect 2731 11645 2743 11648
rect 2685 11639 2743 11645
rect 3602 11636 3608 11648
rect 3660 11636 3666 11688
rect 3697 11679 3755 11685
rect 3697 11645 3709 11679
rect 3743 11645 3755 11679
rect 3697 11639 3755 11645
rect 3881 11679 3939 11685
rect 3881 11645 3893 11679
rect 3927 11645 3939 11679
rect 3881 11639 3939 11645
rect 3712 11608 3740 11639
rect 3786 11608 3792 11620
rect 3712 11580 3792 11608
rect 3786 11568 3792 11580
rect 3844 11568 3850 11620
rect 3896 11608 3924 11639
rect 3970 11636 3976 11688
rect 4028 11636 4034 11688
rect 4157 11679 4215 11685
rect 4157 11645 4169 11679
rect 4203 11676 4215 11679
rect 4338 11676 4344 11688
rect 4203 11648 4344 11676
rect 4203 11645 4215 11648
rect 4157 11639 4215 11645
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 4798 11636 4804 11688
rect 4856 11676 4862 11688
rect 4985 11679 5043 11685
rect 4985 11676 4997 11679
rect 4856 11648 4997 11676
rect 4856 11636 4862 11648
rect 4985 11645 4997 11648
rect 5031 11645 5043 11679
rect 5721 11679 5779 11685
rect 5721 11676 5733 11679
rect 4985 11639 5043 11645
rect 5092 11648 5733 11676
rect 5092 11608 5120 11648
rect 5721 11645 5733 11648
rect 5767 11645 5779 11679
rect 5721 11639 5779 11645
rect 6546 11636 6552 11688
rect 6604 11636 6610 11688
rect 7190 11636 7196 11688
rect 7248 11636 7254 11688
rect 7374 11636 7380 11688
rect 7432 11636 7438 11688
rect 7576 11685 7604 11716
rect 7561 11679 7619 11685
rect 7561 11645 7573 11679
rect 7607 11645 7619 11679
rect 7561 11639 7619 11645
rect 7650 11636 7656 11688
rect 7708 11676 7714 11688
rect 8110 11685 8116 11688
rect 8067 11679 8116 11685
rect 7708 11648 7753 11676
rect 7708 11636 7714 11648
rect 8067 11645 8079 11679
rect 8113 11645 8116 11679
rect 8067 11639 8116 11645
rect 8110 11636 8116 11639
rect 8168 11636 8174 11688
rect 8202 11636 8208 11688
rect 8260 11676 8266 11688
rect 8389 11679 8447 11685
rect 8389 11676 8401 11679
rect 8260 11648 8401 11676
rect 8260 11636 8266 11648
rect 8389 11645 8401 11648
rect 8435 11645 8447 11679
rect 8389 11639 8447 11645
rect 8662 11636 8668 11688
rect 8720 11636 8726 11688
rect 9140 11676 9168 11716
rect 9398 11704 9404 11756
rect 9456 11704 9462 11756
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9640 11716 9781 11744
rect 9640 11704 9646 11716
rect 9769 11713 9781 11716
rect 9815 11713 9827 11747
rect 12084 11744 12112 11840
rect 9769 11707 9827 11713
rect 11440 11716 12112 11744
rect 9493 11679 9551 11685
rect 9140 11648 9260 11676
rect 3896 11580 4016 11608
rect 3988 11540 4016 11580
rect 4632 11580 5120 11608
rect 5169 11611 5227 11617
rect 4632 11552 4660 11580
rect 5169 11577 5181 11611
rect 5215 11608 5227 11611
rect 5442 11608 5448 11620
rect 5215 11580 5448 11608
rect 5215 11577 5227 11580
rect 5169 11571 5227 11577
rect 4522 11540 4528 11552
rect 3988 11512 4528 11540
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 4614 11500 4620 11552
rect 4672 11500 4678 11552
rect 4706 11500 4712 11552
rect 4764 11500 4770 11552
rect 4801 11543 4859 11549
rect 4801 11509 4813 11543
rect 4847 11540 4859 11543
rect 5184 11540 5212 11571
rect 5442 11568 5448 11580
rect 5500 11568 5506 11620
rect 4847 11512 5212 11540
rect 4847 11509 4859 11512
rect 4801 11503 4859 11509
rect 6362 11500 6368 11552
rect 6420 11500 6426 11552
rect 7208 11540 7236 11636
rect 7392 11608 7420 11636
rect 7837 11611 7895 11617
rect 7837 11608 7849 11611
rect 7392 11580 7849 11608
rect 7837 11577 7849 11580
rect 7883 11577 7895 11611
rect 7837 11571 7895 11577
rect 7929 11611 7987 11617
rect 7929 11577 7941 11611
rect 7975 11608 7987 11611
rect 8294 11608 8300 11620
rect 7975 11580 8300 11608
rect 7975 11577 7987 11580
rect 7929 11571 7987 11577
rect 8294 11568 8300 11580
rect 8352 11568 8358 11620
rect 8481 11543 8539 11549
rect 8481 11540 8493 11543
rect 7208 11512 8493 11540
rect 8481 11509 8493 11512
rect 8527 11509 8539 11543
rect 8481 11503 8539 11509
rect 9122 11500 9128 11552
rect 9180 11500 9186 11552
rect 9232 11540 9260 11648
rect 9493 11645 9505 11679
rect 9539 11676 9551 11679
rect 9674 11676 9680 11688
rect 9539 11648 9680 11676
rect 9539 11645 9551 11648
rect 9493 11639 9551 11645
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 11440 11685 11468 11716
rect 11425 11679 11483 11685
rect 11425 11645 11437 11679
rect 11471 11645 11483 11679
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 11425 11639 11483 11645
rect 11992 11648 12081 11676
rect 9582 11568 9588 11620
rect 9640 11608 9646 11620
rect 9861 11611 9919 11617
rect 9861 11608 9873 11611
rect 9640 11580 9873 11608
rect 9640 11568 9646 11580
rect 9861 11577 9873 11580
rect 9907 11608 9919 11611
rect 10413 11611 10471 11617
rect 10413 11608 10425 11611
rect 9907 11580 10425 11608
rect 9907 11577 9919 11580
rect 9861 11571 9919 11577
rect 10413 11577 10425 11580
rect 10459 11577 10471 11611
rect 10413 11571 10471 11577
rect 10686 11568 10692 11620
rect 10744 11568 10750 11620
rect 11992 11552 12020 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 9950 11540 9956 11552
rect 9232 11512 9956 11540
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 11146 11500 11152 11552
rect 11204 11500 11210 11552
rect 11330 11500 11336 11552
rect 11388 11500 11394 11552
rect 11422 11500 11428 11552
rect 11480 11540 11486 11552
rect 11609 11543 11667 11549
rect 11609 11540 11621 11543
rect 11480 11512 11621 11540
rect 11480 11500 11486 11512
rect 11609 11509 11621 11512
rect 11655 11509 11667 11543
rect 11609 11503 11667 11509
rect 11974 11500 11980 11552
rect 12032 11500 12038 11552
rect 552 11450 15520 11472
rect 552 11398 4100 11450
rect 4152 11398 4164 11450
rect 4216 11398 4228 11450
rect 4280 11398 4292 11450
rect 4344 11398 4356 11450
rect 4408 11398 7802 11450
rect 7854 11398 7866 11450
rect 7918 11398 7930 11450
rect 7982 11398 7994 11450
rect 8046 11398 8058 11450
rect 8110 11398 11504 11450
rect 11556 11398 11568 11450
rect 11620 11398 11632 11450
rect 11684 11398 11696 11450
rect 11748 11398 11760 11450
rect 11812 11398 15206 11450
rect 15258 11398 15270 11450
rect 15322 11398 15334 11450
rect 15386 11398 15398 11450
rect 15450 11398 15462 11450
rect 15514 11398 15520 11450
rect 552 11376 15520 11398
rect 2130 11296 2136 11348
rect 2188 11336 2194 11348
rect 2188 11308 2452 11336
rect 2188 11296 2194 11308
rect 2130 11160 2136 11212
rect 2188 11209 2194 11212
rect 2424 11209 2452 11308
rect 3878 11296 3884 11348
rect 3936 11336 3942 11348
rect 4157 11339 4215 11345
rect 4157 11336 4169 11339
rect 3936 11308 4169 11336
rect 3936 11296 3942 11308
rect 4157 11305 4169 11308
rect 4203 11305 4215 11339
rect 4991 11339 5049 11345
rect 4991 11336 5003 11339
rect 4157 11299 4215 11305
rect 4356 11308 5003 11336
rect 3436 11240 3924 11268
rect 2188 11200 2200 11209
rect 2409 11203 2467 11209
rect 2188 11172 2233 11200
rect 2188 11163 2200 11172
rect 2409 11169 2421 11203
rect 2455 11200 2467 11203
rect 3326 11200 3332 11212
rect 2455 11172 3332 11200
rect 2455 11169 2467 11172
rect 2409 11163 2467 11169
rect 2188 11160 2194 11163
rect 3326 11160 3332 11172
rect 3384 11160 3390 11212
rect 3436 11209 3464 11240
rect 3421 11203 3479 11209
rect 3421 11169 3433 11203
rect 3467 11169 3479 11203
rect 3421 11163 3479 11169
rect 3510 11160 3516 11212
rect 3568 11160 3574 11212
rect 3697 11203 3755 11209
rect 3697 11169 3709 11203
rect 3743 11169 3755 11203
rect 3697 11163 3755 11169
rect 3053 11135 3111 11141
rect 3053 11132 3065 11135
rect 2424 11104 3065 11132
rect 1029 10999 1087 11005
rect 1029 10965 1041 10999
rect 1075 10996 1087 10999
rect 2424 10996 2452 11104
rect 3053 11101 3065 11104
rect 3099 11101 3111 11135
rect 3053 11095 3111 11101
rect 3068 11064 3096 11095
rect 3528 11064 3556 11160
rect 3068 11036 3556 11064
rect 1075 10968 2452 10996
rect 2501 10999 2559 11005
rect 1075 10965 1087 10968
rect 1029 10959 1087 10965
rect 2501 10965 2513 10999
rect 2547 10996 2559 10999
rect 2682 10996 2688 11008
rect 2547 10968 2688 10996
rect 2547 10965 2559 10968
rect 2501 10959 2559 10965
rect 2682 10956 2688 10968
rect 2740 10956 2746 11008
rect 3234 10956 3240 11008
rect 3292 10956 3298 11008
rect 3712 10996 3740 11163
rect 3786 11160 3792 11212
rect 3844 11160 3850 11212
rect 3896 11209 3924 11240
rect 3970 11228 3976 11280
rect 4028 11268 4034 11280
rect 4356 11268 4384 11308
rect 4991 11305 5003 11308
rect 5037 11305 5049 11339
rect 4991 11299 5049 11305
rect 5077 11339 5135 11345
rect 5077 11305 5089 11339
rect 5123 11336 5135 11339
rect 5258 11336 5264 11348
rect 5123 11308 5264 11336
rect 5123 11305 5135 11308
rect 5077 11299 5135 11305
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 10965 11339 11023 11345
rect 10965 11336 10977 11339
rect 8720 11308 10977 11336
rect 8720 11296 8726 11308
rect 4028 11240 4384 11268
rect 6264 11271 6322 11277
rect 4028 11228 4034 11240
rect 3881 11203 3939 11209
rect 3881 11169 3893 11203
rect 3927 11200 3939 11203
rect 3927 11172 4016 11200
rect 3927 11169 3939 11172
rect 3881 11163 3939 11169
rect 3988 11132 4016 11172
rect 4062 11160 4068 11212
rect 4120 11160 4126 11212
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11169 4399 11203
rect 4792 11203 4850 11209
rect 4792 11200 4804 11203
rect 4341 11163 4399 11169
rect 4724 11172 4804 11200
rect 4356 11132 4384 11163
rect 3988 11104 4108 11132
rect 3881 10999 3939 11005
rect 3881 10996 3893 10999
rect 3712 10968 3893 10996
rect 3881 10965 3893 10968
rect 3927 10965 3939 10999
rect 3881 10959 3939 10965
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 4080 10996 4108 11104
rect 4264 11104 4384 11132
rect 4264 11076 4292 11104
rect 4522 11092 4528 11144
rect 4580 11092 4586 11144
rect 4614 11092 4620 11144
rect 4672 11092 4678 11144
rect 4246 11024 4252 11076
rect 4304 11024 4310 11076
rect 4430 11024 4436 11076
rect 4488 11024 4494 11076
rect 4540 10996 4568 11092
rect 4724 11064 4752 11172
rect 4792 11169 4804 11172
rect 4838 11169 4850 11203
rect 4890 11194 4896 11246
rect 4948 11194 4954 11246
rect 6264 11237 6276 11271
rect 6310 11268 6322 11271
rect 6362 11268 6368 11280
rect 6310 11240 6368 11268
rect 6310 11237 6322 11240
rect 6264 11231 6322 11237
rect 6362 11228 6368 11240
rect 6420 11228 6426 11280
rect 9674 11268 9680 11280
rect 8312 11240 9680 11268
rect 8312 11212 8340 11240
rect 5169 11203 5227 11209
rect 4792 11163 4850 11169
rect 5169 11169 5181 11203
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11200 5503 11203
rect 5534 11200 5540 11212
rect 5491 11172 5540 11200
rect 5491 11169 5503 11172
rect 5445 11163 5503 11169
rect 4982 11092 4988 11144
rect 5040 11132 5046 11144
rect 5184 11132 5212 11163
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 8294 11160 8300 11212
rect 8352 11160 8358 11212
rect 8938 11160 8944 11212
rect 8996 11160 9002 11212
rect 9232 11209 9260 11240
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 9217 11203 9275 11209
rect 9217 11169 9229 11203
rect 9263 11169 9275 11203
rect 9217 11163 9275 11169
rect 9309 11203 9367 11209
rect 9309 11169 9321 11203
rect 9355 11200 9367 11203
rect 9398 11200 9404 11212
rect 9355 11172 9404 11200
rect 9355 11169 9367 11172
rect 9309 11163 9367 11169
rect 9398 11160 9404 11172
rect 9456 11160 9462 11212
rect 9784 11209 9812 11308
rect 10965 11305 10977 11308
rect 11011 11305 11023 11339
rect 10965 11299 11023 11305
rect 12710 11296 12716 11348
rect 12768 11336 12774 11348
rect 12768 11308 13124 11336
rect 12768 11296 12774 11308
rect 10686 11228 10692 11280
rect 10744 11228 10750 11280
rect 12437 11271 12495 11277
rect 12437 11237 12449 11271
rect 12483 11268 12495 11271
rect 12483 11240 12756 11268
rect 12483 11237 12495 11240
rect 12437 11231 12495 11237
rect 9769 11203 9827 11209
rect 9769 11169 9781 11203
rect 9815 11169 9827 11203
rect 9769 11163 9827 11169
rect 9950 11160 9956 11212
rect 10008 11160 10014 11212
rect 10042 11160 10048 11212
rect 10100 11160 10106 11212
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11200 10379 11203
rect 10704 11200 10732 11228
rect 10367 11172 10732 11200
rect 10367 11169 10379 11172
rect 10321 11163 10379 11169
rect 11146 11160 11152 11212
rect 11204 11160 11210 11212
rect 11517 11203 11575 11209
rect 11517 11169 11529 11203
rect 11563 11169 11575 11203
rect 11517 11163 11575 11169
rect 5040 11104 5212 11132
rect 5040 11092 5046 11104
rect 5718 11092 5724 11144
rect 5776 11132 5782 11144
rect 5997 11135 6055 11141
rect 5997 11132 6009 11135
rect 5776 11104 6009 11132
rect 5776 11092 5782 11104
rect 5997 11101 6009 11104
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 9030 11092 9036 11144
rect 9088 11092 9094 11144
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11132 10839 11135
rect 10870 11132 10876 11144
rect 10827 11104 10876 11132
rect 10827 11101 10839 11104
rect 10781 11095 10839 11101
rect 10870 11092 10876 11104
rect 10928 11132 10934 11144
rect 11532 11132 11560 11163
rect 11974 11160 11980 11212
rect 12032 11160 12038 11212
rect 12345 11203 12403 11209
rect 12345 11169 12357 11203
rect 12391 11169 12403 11203
rect 12345 11163 12403 11169
rect 12529 11203 12587 11209
rect 12529 11169 12541 11203
rect 12575 11169 12587 11203
rect 12529 11163 12587 11169
rect 10928 11104 11560 11132
rect 10928 11092 10934 11104
rect 11882 11092 11888 11144
rect 11940 11092 11946 11144
rect 12360 11132 12388 11163
rect 12434 11132 12440 11144
rect 12360 11104 12440 11132
rect 12434 11092 12440 11104
rect 12492 11092 12498 11144
rect 12544 11132 12572 11163
rect 12618 11160 12624 11212
rect 12676 11160 12682 11212
rect 12728 11209 12756 11240
rect 12714 11203 12772 11209
rect 12714 11169 12726 11203
rect 12760 11169 12772 11203
rect 12714 11163 12772 11169
rect 12894 11160 12900 11212
rect 12952 11160 12958 11212
rect 12986 11160 12992 11212
rect 13044 11160 13050 11212
rect 13096 11209 13124 11308
rect 13086 11203 13144 11209
rect 13086 11169 13098 11203
rect 13132 11169 13144 11203
rect 13086 11163 13144 11169
rect 13262 11160 13268 11212
rect 13320 11200 13326 11212
rect 13357 11203 13415 11209
rect 13357 11200 13369 11203
rect 13320 11172 13369 11200
rect 13320 11160 13326 11172
rect 13357 11169 13369 11172
rect 13403 11169 13415 11203
rect 14274 11200 14280 11212
rect 13357 11163 13415 11169
rect 13464 11172 14280 11200
rect 13464 11132 13492 11172
rect 14274 11160 14280 11172
rect 14332 11160 14338 11212
rect 12544 11104 13492 11132
rect 13630 11092 13636 11144
rect 13688 11092 13694 11144
rect 9493 11067 9551 11073
rect 4724 11036 4936 11064
rect 4028 10968 4568 10996
rect 4908 10996 4936 11036
rect 9493 11033 9505 11067
rect 9539 11064 9551 11067
rect 9861 11067 9919 11073
rect 9861 11064 9873 11067
rect 9539 11036 9873 11064
rect 9539 11033 9551 11036
rect 9493 11027 9551 11033
rect 9861 11033 9873 11036
rect 9907 11033 9919 11067
rect 9861 11027 9919 11033
rect 5350 10996 5356 11008
rect 4908 10968 5356 10996
rect 4028 10956 4034 10968
rect 5350 10956 5356 10968
rect 5408 10956 5414 11008
rect 5810 10956 5816 11008
rect 5868 10996 5874 11008
rect 6914 10996 6920 11008
rect 5868 10968 6920 10996
rect 5868 10956 5874 10968
rect 6914 10956 6920 10968
rect 6972 10996 6978 11008
rect 7377 10999 7435 11005
rect 7377 10996 7389 10999
rect 6972 10968 7389 10996
rect 6972 10956 6978 10968
rect 7377 10965 7389 10968
rect 7423 10965 7435 10999
rect 7377 10959 7435 10965
rect 9306 10956 9312 11008
rect 9364 10996 9370 11008
rect 9585 10999 9643 11005
rect 9585 10996 9597 10999
rect 9364 10968 9597 10996
rect 9364 10956 9370 10968
rect 9585 10965 9597 10968
rect 9631 10965 9643 10999
rect 9585 10959 9643 10965
rect 10594 10956 10600 11008
rect 10652 10956 10658 11008
rect 11054 10956 11060 11008
rect 11112 10996 11118 11008
rect 11149 10999 11207 11005
rect 11149 10996 11161 10999
rect 11112 10968 11161 10996
rect 11112 10956 11118 10968
rect 11149 10965 11161 10968
rect 11195 10996 11207 10999
rect 11609 10999 11667 11005
rect 11609 10996 11621 10999
rect 11195 10968 11621 10996
rect 11195 10965 11207 10968
rect 11149 10959 11207 10965
rect 11609 10965 11621 10968
rect 11655 10965 11667 10999
rect 11609 10959 11667 10965
rect 13265 10999 13323 11005
rect 13265 10965 13277 10999
rect 13311 10996 13323 10999
rect 13998 10996 14004 11008
rect 13311 10968 14004 10996
rect 13311 10965 13323 10968
rect 13265 10959 13323 10965
rect 13998 10956 14004 10968
rect 14056 10956 14062 11008
rect 14918 10956 14924 11008
rect 14976 10956 14982 11008
rect 552 10906 15364 10928
rect 552 10854 2249 10906
rect 2301 10854 2313 10906
rect 2365 10854 2377 10906
rect 2429 10854 2441 10906
rect 2493 10854 2505 10906
rect 2557 10854 5951 10906
rect 6003 10854 6015 10906
rect 6067 10854 6079 10906
rect 6131 10854 6143 10906
rect 6195 10854 6207 10906
rect 6259 10854 9653 10906
rect 9705 10854 9717 10906
rect 9769 10854 9781 10906
rect 9833 10854 9845 10906
rect 9897 10854 9909 10906
rect 9961 10854 13355 10906
rect 13407 10854 13419 10906
rect 13471 10854 13483 10906
rect 13535 10854 13547 10906
rect 13599 10854 13611 10906
rect 13663 10854 15364 10906
rect 552 10832 15364 10854
rect 2130 10752 2136 10804
rect 2188 10792 2194 10804
rect 2317 10795 2375 10801
rect 2317 10792 2329 10795
rect 2188 10764 2329 10792
rect 2188 10752 2194 10764
rect 2317 10761 2329 10764
rect 2363 10761 2375 10795
rect 3234 10792 3240 10804
rect 2317 10755 2375 10761
rect 2746 10764 3240 10792
rect 2746 10656 2774 10764
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 3697 10795 3755 10801
rect 3697 10792 3709 10795
rect 3384 10764 3709 10792
rect 3384 10752 3390 10764
rect 3697 10761 3709 10764
rect 3743 10792 3755 10795
rect 3743 10764 4384 10792
rect 3743 10761 3755 10764
rect 3697 10755 3755 10761
rect 3786 10684 3792 10736
rect 3844 10724 3850 10736
rect 4246 10724 4252 10736
rect 3844 10696 4252 10724
rect 3844 10684 3850 10696
rect 4246 10684 4252 10696
rect 4304 10684 4310 10736
rect 4356 10724 4384 10764
rect 4430 10752 4436 10804
rect 4488 10792 4494 10804
rect 5077 10795 5135 10801
rect 5077 10792 5089 10795
rect 4488 10764 5089 10792
rect 4488 10752 4494 10764
rect 5077 10761 5089 10764
rect 5123 10761 5135 10795
rect 5718 10792 5724 10804
rect 5077 10755 5135 10761
rect 5184 10764 5724 10792
rect 5184 10724 5212 10764
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 6365 10795 6423 10801
rect 6365 10761 6377 10795
rect 6411 10792 6423 10795
rect 6546 10792 6552 10804
rect 6411 10764 6552 10792
rect 6411 10761 6423 10764
rect 6365 10755 6423 10761
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 8113 10795 8171 10801
rect 7208 10764 8064 10792
rect 4356 10696 5212 10724
rect 5258 10684 5264 10736
rect 5316 10724 5322 10736
rect 5442 10724 5448 10736
rect 5316 10696 5448 10724
rect 5316 10684 5322 10696
rect 5442 10684 5448 10696
rect 5500 10724 5506 10736
rect 5810 10724 5816 10736
rect 5500 10696 5816 10724
rect 5500 10684 5506 10696
rect 5810 10684 5816 10696
rect 5868 10684 5874 10736
rect 7208 10724 7236 10764
rect 6012 10696 7236 10724
rect 2608 10628 2774 10656
rect 2608 10597 2636 10628
rect 3694 10616 3700 10668
rect 3752 10656 3758 10668
rect 4614 10656 4620 10668
rect 3752 10628 4620 10656
rect 3752 10616 3758 10628
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 6012 10656 6040 10696
rect 6362 10656 6368 10668
rect 5000 10628 6040 10656
rect 6104 10628 6368 10656
rect 5000 10600 5028 10628
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10557 2651 10591
rect 2593 10551 2651 10557
rect 2682 10548 2688 10600
rect 2740 10548 2746 10600
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 2869 10591 2927 10597
rect 2869 10588 2881 10591
rect 2832 10560 2881 10588
rect 2832 10548 2838 10560
rect 2869 10557 2881 10560
rect 2915 10557 2927 10591
rect 2869 10551 2927 10557
rect 4982 10548 4988 10600
rect 5040 10548 5046 10600
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10557 5319 10591
rect 5261 10551 5319 10557
rect 2317 10523 2375 10529
rect 2317 10489 2329 10523
rect 2363 10520 2375 10523
rect 3142 10520 3148 10532
rect 2363 10492 3148 10520
rect 2363 10489 2375 10492
rect 2317 10483 2375 10489
rect 3142 10480 3148 10492
rect 3200 10480 3206 10532
rect 5276 10520 5304 10551
rect 5350 10548 5356 10600
rect 5408 10548 5414 10600
rect 5810 10588 5816 10600
rect 5736 10560 5816 10588
rect 5276 10492 5396 10520
rect 5368 10464 5396 10492
rect 5442 10480 5448 10532
rect 5500 10520 5506 10532
rect 5736 10529 5764 10560
rect 5810 10548 5816 10560
rect 5868 10548 5874 10600
rect 6104 10597 6132 10628
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 8036 10656 8064 10764
rect 8113 10761 8125 10795
rect 8159 10792 8171 10795
rect 8294 10792 8300 10804
rect 8159 10764 8300 10792
rect 8159 10761 8171 10764
rect 8113 10755 8171 10761
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 9861 10795 9919 10801
rect 9861 10761 9873 10795
rect 9907 10792 9919 10795
rect 10318 10792 10324 10804
rect 9907 10764 10324 10792
rect 9907 10761 9919 10764
rect 9861 10755 9919 10761
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 12894 10752 12900 10804
rect 12952 10752 12958 10804
rect 13541 10795 13599 10801
rect 13541 10761 13553 10795
rect 13587 10792 13599 10795
rect 13722 10792 13728 10804
rect 13587 10764 13728 10792
rect 13587 10761 13599 10764
rect 13541 10755 13599 10761
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 14274 10752 14280 10804
rect 14332 10752 14338 10804
rect 14461 10795 14519 10801
rect 14461 10761 14473 10795
rect 14507 10792 14519 10795
rect 14550 10792 14556 10804
rect 14507 10764 14556 10792
rect 14507 10761 14519 10764
rect 14461 10755 14519 10761
rect 10042 10684 10048 10736
rect 10100 10724 10106 10736
rect 10505 10727 10563 10733
rect 10505 10724 10517 10727
rect 10100 10696 10517 10724
rect 10100 10684 10106 10696
rect 10505 10693 10517 10696
rect 10551 10693 10563 10727
rect 11609 10727 11667 10733
rect 11609 10724 11621 10727
rect 10505 10687 10563 10693
rect 10612 10696 11621 10724
rect 8036 10628 8432 10656
rect 8404 10600 8432 10628
rect 8846 10616 8852 10668
rect 8904 10656 8910 10668
rect 10612 10656 10640 10696
rect 11609 10693 11621 10696
rect 11655 10724 11667 10727
rect 14090 10724 14096 10736
rect 11655 10696 14096 10724
rect 11655 10693 11667 10696
rect 11609 10687 11667 10693
rect 14090 10684 14096 10696
rect 14148 10684 14154 10736
rect 11054 10656 11060 10668
rect 8904 10628 10640 10656
rect 10796 10628 11060 10656
rect 8904 10616 8910 10628
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10557 6147 10591
rect 6089 10551 6147 10557
rect 6181 10591 6239 10597
rect 6181 10557 6193 10591
rect 6227 10588 6239 10591
rect 6457 10591 6515 10597
rect 6457 10588 6469 10591
rect 6227 10560 6469 10588
rect 6227 10557 6239 10560
rect 6181 10551 6239 10557
rect 6457 10557 6469 10560
rect 6503 10557 6515 10591
rect 6457 10551 6515 10557
rect 6638 10548 6644 10600
rect 6696 10548 6702 10600
rect 6914 10548 6920 10600
rect 6972 10597 6978 10600
rect 6972 10591 7001 10597
rect 6989 10557 7001 10591
rect 6972 10551 7001 10557
rect 7101 10591 7159 10597
rect 7101 10557 7113 10591
rect 7147 10588 7159 10591
rect 7466 10588 7472 10600
rect 7147 10560 7472 10588
rect 7147 10557 7159 10560
rect 7101 10551 7159 10557
rect 6972 10548 6978 10551
rect 7466 10548 7472 10560
rect 7524 10548 7530 10600
rect 8205 10591 8263 10597
rect 8205 10557 8217 10591
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 5537 10523 5595 10529
rect 5537 10520 5549 10523
rect 5500 10492 5549 10520
rect 5500 10480 5506 10492
rect 5537 10489 5549 10492
rect 5583 10489 5595 10523
rect 5537 10483 5595 10489
rect 5721 10523 5779 10529
rect 5721 10489 5733 10523
rect 5767 10489 5779 10523
rect 5721 10483 5779 10489
rect 5905 10523 5963 10529
rect 5905 10489 5917 10523
rect 5951 10520 5963 10523
rect 6733 10523 6791 10529
rect 6733 10520 6745 10523
rect 5951 10492 6745 10520
rect 5951 10489 5963 10492
rect 5905 10483 5963 10489
rect 6733 10489 6745 10492
rect 6779 10489 6791 10523
rect 6733 10483 6791 10489
rect 6822 10480 6828 10532
rect 6880 10480 6886 10532
rect 8220 10464 8248 10551
rect 8386 10548 8392 10600
rect 8444 10548 8450 10600
rect 10796 10597 10824 10628
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 14476 10656 14504 10755
rect 14550 10752 14556 10764
rect 14608 10752 14614 10804
rect 13280 10628 14504 10656
rect 10781 10591 10839 10597
rect 10781 10557 10793 10591
rect 10827 10557 10839 10591
rect 10781 10551 10839 10557
rect 10870 10548 10876 10600
rect 10928 10548 10934 10600
rect 10965 10591 11023 10597
rect 10965 10557 10977 10591
rect 11011 10557 11023 10591
rect 10965 10551 11023 10557
rect 11149 10591 11207 10597
rect 11149 10557 11161 10591
rect 11195 10588 11207 10591
rect 11422 10588 11428 10600
rect 11195 10560 11428 10588
rect 11195 10557 11207 10560
rect 11149 10551 11207 10557
rect 10980 10520 11008 10551
rect 11422 10548 11428 10560
rect 11480 10548 11486 10600
rect 13280 10597 13308 10628
rect 13081 10591 13139 10597
rect 13081 10557 13093 10591
rect 13127 10557 13139 10591
rect 13081 10551 13139 10557
rect 13265 10591 13323 10597
rect 13265 10557 13277 10591
rect 13311 10557 13323 10591
rect 13265 10551 13323 10557
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10588 13415 10591
rect 13722 10588 13728 10600
rect 13403 10560 13728 10588
rect 13403 10557 13415 10560
rect 13357 10551 13415 10557
rect 11330 10520 11336 10532
rect 10980 10492 11336 10520
rect 11330 10480 11336 10492
rect 11388 10480 11394 10532
rect 13096 10520 13124 10551
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 13832 10520 13860 10551
rect 13906 10548 13912 10600
rect 13964 10548 13970 10600
rect 13998 10548 14004 10600
rect 14056 10548 14062 10600
rect 14182 10548 14188 10600
rect 14240 10548 14246 10600
rect 14645 10523 14703 10529
rect 14645 10520 14657 10523
rect 13096 10492 14657 10520
rect 14645 10489 14657 10492
rect 14691 10520 14703 10523
rect 14918 10520 14924 10532
rect 14691 10492 14924 10520
rect 14691 10489 14703 10492
rect 14645 10483 14703 10489
rect 14918 10480 14924 10492
rect 14976 10480 14982 10532
rect 2501 10455 2559 10461
rect 2501 10421 2513 10455
rect 2547 10452 2559 10455
rect 2777 10455 2835 10461
rect 2777 10452 2789 10455
rect 2547 10424 2789 10452
rect 2547 10421 2559 10424
rect 2501 10415 2559 10421
rect 2777 10421 2789 10424
rect 2823 10421 2835 10455
rect 2777 10415 2835 10421
rect 5350 10412 5356 10464
rect 5408 10412 5414 10464
rect 8202 10412 8208 10464
rect 8260 10412 8266 10464
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 14274 10452 14280 10464
rect 13780 10424 14280 10452
rect 13780 10412 13786 10424
rect 14274 10412 14280 10424
rect 14332 10452 14338 10464
rect 14435 10455 14493 10461
rect 14435 10452 14447 10455
rect 14332 10424 14447 10452
rect 14332 10412 14338 10424
rect 14435 10421 14447 10424
rect 14481 10421 14493 10455
rect 14435 10415 14493 10421
rect 552 10362 15520 10384
rect 552 10310 4100 10362
rect 4152 10310 4164 10362
rect 4216 10310 4228 10362
rect 4280 10310 4292 10362
rect 4344 10310 4356 10362
rect 4408 10310 7802 10362
rect 7854 10310 7866 10362
rect 7918 10310 7930 10362
rect 7982 10310 7994 10362
rect 8046 10310 8058 10362
rect 8110 10310 11504 10362
rect 11556 10310 11568 10362
rect 11620 10310 11632 10362
rect 11684 10310 11696 10362
rect 11748 10310 11760 10362
rect 11812 10310 15206 10362
rect 15258 10310 15270 10362
rect 15322 10310 15334 10362
rect 15386 10310 15398 10362
rect 15450 10310 15462 10362
rect 15514 10310 15520 10362
rect 552 10288 15520 10310
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 4341 10251 4399 10257
rect 4341 10248 4353 10251
rect 4028 10220 4353 10248
rect 4028 10208 4034 10220
rect 4341 10217 4353 10220
rect 4387 10217 4399 10251
rect 4341 10211 4399 10217
rect 5258 10208 5264 10260
rect 5316 10208 5322 10260
rect 5350 10208 5356 10260
rect 5408 10248 5414 10260
rect 6638 10248 6644 10260
rect 5408 10220 6644 10248
rect 5408 10208 5414 10220
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 9122 10208 9128 10260
rect 9180 10208 9186 10260
rect 9306 10208 9312 10260
rect 9364 10208 9370 10260
rect 4509 10183 4567 10189
rect 4509 10149 4521 10183
rect 4555 10180 4567 10183
rect 4555 10152 4660 10180
rect 4555 10149 4567 10152
rect 4509 10143 4567 10149
rect 4632 10056 4660 10152
rect 4706 10140 4712 10192
rect 4764 10140 4770 10192
rect 5074 10072 5080 10124
rect 5132 10112 5138 10124
rect 5276 10121 5304 10208
rect 5261 10115 5319 10121
rect 5261 10112 5273 10115
rect 5132 10084 5273 10112
rect 5132 10072 5138 10084
rect 5261 10081 5273 10084
rect 5307 10081 5319 10115
rect 5261 10075 5319 10081
rect 5442 10072 5448 10124
rect 5500 10072 5506 10124
rect 8757 10115 8815 10121
rect 8757 10081 8769 10115
rect 8803 10081 8815 10115
rect 8757 10075 8815 10081
rect 8941 10115 8999 10121
rect 8941 10081 8953 10115
rect 8987 10112 8999 10115
rect 9033 10115 9091 10121
rect 9033 10112 9045 10115
rect 8987 10084 9045 10112
rect 8987 10081 8999 10084
rect 8941 10075 8999 10081
rect 9033 10081 9045 10084
rect 9079 10112 9091 10115
rect 9140 10112 9168 10208
rect 9079 10084 9168 10112
rect 9217 10115 9275 10121
rect 9079 10081 9091 10084
rect 9033 10075 9091 10081
rect 9217 10081 9229 10115
rect 9263 10112 9275 10115
rect 9324 10112 9352 10208
rect 9263 10084 9352 10112
rect 9401 10115 9459 10121
rect 9263 10081 9275 10084
rect 9217 10075 9275 10081
rect 9401 10081 9413 10115
rect 9447 10081 9459 10115
rect 9401 10075 9459 10081
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 5460 10044 5488 10072
rect 4672 10016 5488 10044
rect 8772 10044 8800 10075
rect 9232 10044 9260 10075
rect 9416 10044 9444 10075
rect 10686 10072 10692 10124
rect 10744 10072 10750 10124
rect 11241 10115 11299 10121
rect 11241 10081 11253 10115
rect 11287 10112 11299 10115
rect 11974 10112 11980 10124
rect 11287 10084 11980 10112
rect 11287 10081 11299 10084
rect 11241 10075 11299 10081
rect 11974 10072 11980 10084
rect 12032 10112 12038 10124
rect 12434 10112 12440 10124
rect 12032 10084 12440 10112
rect 12032 10072 12038 10084
rect 12434 10072 12440 10084
rect 12492 10072 12498 10124
rect 12618 10072 12624 10124
rect 12676 10072 12682 10124
rect 8772 10016 9260 10044
rect 9324 10016 9444 10044
rect 10704 10044 10732 10072
rect 11333 10047 11391 10053
rect 10704 10016 11054 10044
rect 4672 10004 4678 10016
rect 5276 9920 5304 10016
rect 6822 9936 6828 9988
rect 6880 9976 6886 9988
rect 8573 9979 8631 9985
rect 8573 9976 8585 9979
rect 6880 9948 8585 9976
rect 6880 9936 6886 9948
rect 8573 9945 8585 9948
rect 8619 9976 8631 9979
rect 9324 9976 9352 10016
rect 8619 9948 9352 9976
rect 11026 9976 11054 10016
rect 11333 10013 11345 10047
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 11348 9976 11376 10007
rect 11026 9948 11376 9976
rect 11440 9976 11468 10007
rect 11514 10004 11520 10056
rect 11572 10004 11578 10056
rect 12636 9976 12664 10072
rect 11440 9948 12664 9976
rect 8619 9945 8631 9948
rect 8573 9939 8631 9945
rect 4525 9911 4583 9917
rect 4525 9877 4537 9911
rect 4571 9908 4583 9911
rect 5074 9908 5080 9920
rect 4571 9880 5080 9908
rect 4571 9877 4583 9880
rect 4525 9871 4583 9877
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 5258 9868 5264 9920
rect 5316 9868 5322 9920
rect 5626 9868 5632 9920
rect 5684 9908 5690 9920
rect 9122 9908 9128 9920
rect 5684 9880 9128 9908
rect 5684 9868 5690 9880
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 9306 9868 9312 9920
rect 9364 9908 9370 9920
rect 9677 9911 9735 9917
rect 9677 9908 9689 9911
rect 9364 9880 9689 9908
rect 9364 9868 9370 9880
rect 9677 9877 9689 9880
rect 9723 9908 9735 9911
rect 11440 9908 11468 9948
rect 9723 9880 11468 9908
rect 11701 9911 11759 9917
rect 9723 9877 9735 9880
rect 9677 9871 9735 9877
rect 11701 9877 11713 9911
rect 11747 9908 11759 9911
rect 11974 9908 11980 9920
rect 11747 9880 11980 9908
rect 11747 9877 11759 9880
rect 11701 9871 11759 9877
rect 11974 9868 11980 9880
rect 12032 9868 12038 9920
rect 552 9818 15364 9840
rect 552 9766 2249 9818
rect 2301 9766 2313 9818
rect 2365 9766 2377 9818
rect 2429 9766 2441 9818
rect 2493 9766 2505 9818
rect 2557 9766 5951 9818
rect 6003 9766 6015 9818
rect 6067 9766 6079 9818
rect 6131 9766 6143 9818
rect 6195 9766 6207 9818
rect 6259 9766 9653 9818
rect 9705 9766 9717 9818
rect 9769 9766 9781 9818
rect 9833 9766 9845 9818
rect 9897 9766 9909 9818
rect 9961 9766 13355 9818
rect 13407 9766 13419 9818
rect 13471 9766 13483 9818
rect 13535 9766 13547 9818
rect 13599 9766 13611 9818
rect 13663 9766 15364 9818
rect 552 9744 15364 9766
rect 4430 9664 4436 9716
rect 4488 9704 4494 9716
rect 4893 9707 4951 9713
rect 4893 9704 4905 9707
rect 4488 9676 4905 9704
rect 4488 9664 4494 9676
rect 4893 9673 4905 9676
rect 4939 9673 4951 9707
rect 4893 9667 4951 9673
rect 5077 9707 5135 9713
rect 5077 9673 5089 9707
rect 5123 9673 5135 9707
rect 5077 9667 5135 9673
rect 3053 9639 3111 9645
rect 3053 9605 3065 9639
rect 3099 9605 3111 9639
rect 3053 9599 3111 9605
rect 3068 9568 3096 9599
rect 3510 9596 3516 9648
rect 3568 9596 3574 9648
rect 4614 9636 4620 9648
rect 3620 9608 4620 9636
rect 3068 9540 3556 9568
rect 1486 9460 1492 9512
rect 1544 9500 1550 9512
rect 1673 9503 1731 9509
rect 1673 9500 1685 9503
rect 1544 9472 1685 9500
rect 1544 9460 1550 9472
rect 1673 9469 1685 9472
rect 1719 9469 1731 9503
rect 1673 9463 1731 9469
rect 3421 9503 3479 9509
rect 3421 9469 3433 9503
rect 3467 9469 3479 9503
rect 3421 9463 3479 9469
rect 1940 9435 1998 9441
rect 1940 9401 1952 9435
rect 1986 9432 1998 9435
rect 3326 9432 3332 9444
rect 1986 9404 3332 9432
rect 1986 9401 1998 9404
rect 1940 9395 1998 9401
rect 3326 9392 3332 9404
rect 3384 9392 3390 9444
rect 3234 9324 3240 9376
rect 3292 9324 3298 9376
rect 3436 9364 3464 9463
rect 3528 9432 3556 9540
rect 3620 9509 3648 9608
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 5092 9580 5120 9667
rect 7926 9664 7932 9716
rect 7984 9704 7990 9716
rect 8202 9704 8208 9716
rect 7984 9676 8208 9704
rect 7984 9664 7990 9676
rect 8202 9664 8208 9676
rect 8260 9704 8266 9716
rect 8573 9707 8631 9713
rect 8573 9704 8585 9707
rect 8260 9676 8585 9704
rect 8260 9664 8266 9676
rect 8573 9673 8585 9676
rect 8619 9704 8631 9707
rect 9030 9704 9036 9716
rect 8619 9676 9036 9704
rect 8619 9673 8631 9676
rect 8573 9667 8631 9673
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 12529 9707 12587 9713
rect 12529 9704 12541 9707
rect 11026 9676 12541 9704
rect 5629 9639 5687 9645
rect 5629 9605 5641 9639
rect 5675 9636 5687 9639
rect 5675 9608 8156 9636
rect 5675 9605 5687 9608
rect 5629 9599 5687 9605
rect 3694 9528 3700 9580
rect 3752 9528 3758 9580
rect 4890 9568 4896 9580
rect 3896 9540 4896 9568
rect 3896 9509 3924 9540
rect 4890 9528 4896 9540
rect 4948 9528 4954 9580
rect 5074 9568 5080 9580
rect 5000 9540 5080 9568
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9469 3663 9503
rect 3605 9463 3663 9469
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 4065 9503 4123 9509
rect 4065 9469 4077 9503
rect 4111 9469 4123 9503
rect 4065 9463 4123 9469
rect 3970 9432 3976 9444
rect 3528 9404 3976 9432
rect 3970 9392 3976 9404
rect 4028 9432 4034 9444
rect 4080 9432 4108 9463
rect 4522 9460 4528 9512
rect 4580 9500 4586 9512
rect 5000 9500 5028 9540
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 8021 9571 8079 9577
rect 8021 9568 8033 9571
rect 6932 9540 8033 9568
rect 4580 9472 5028 9500
rect 4580 9460 4586 9472
rect 5258 9460 5264 9512
rect 5316 9460 5322 9512
rect 5445 9503 5503 9509
rect 5445 9469 5457 9503
rect 5491 9469 5503 9503
rect 5445 9463 5503 9469
rect 4709 9435 4767 9441
rect 4709 9432 4721 9435
rect 4028 9404 4721 9432
rect 4028 9392 4034 9404
rect 4709 9401 4721 9404
rect 4755 9401 4767 9435
rect 4709 9395 4767 9401
rect 4798 9392 4804 9444
rect 4856 9392 4862 9444
rect 3786 9364 3792 9376
rect 3436 9336 3792 9364
rect 3786 9324 3792 9336
rect 3844 9324 3850 9376
rect 4614 9324 4620 9376
rect 4672 9324 4678 9376
rect 4816 9364 4844 9392
rect 4909 9367 4967 9373
rect 4909 9364 4921 9367
rect 4816 9336 4921 9364
rect 4909 9333 4921 9336
rect 4955 9364 4967 9367
rect 5460 9364 5488 9463
rect 5626 9460 5632 9512
rect 5684 9500 5690 9512
rect 5721 9503 5779 9509
rect 5721 9500 5733 9503
rect 5684 9472 5733 9500
rect 5684 9460 5690 9472
rect 5721 9469 5733 9472
rect 5767 9469 5779 9503
rect 5721 9463 5779 9469
rect 6454 9460 6460 9512
rect 6512 9460 6518 9512
rect 6932 9509 6960 9540
rect 8021 9537 8033 9540
rect 8067 9537 8079 9571
rect 8021 9531 8079 9537
rect 6917 9503 6975 9509
rect 6917 9469 6929 9503
rect 6963 9469 6975 9503
rect 6917 9463 6975 9469
rect 7098 9460 7104 9512
rect 7156 9460 7162 9512
rect 7377 9503 7435 9509
rect 7377 9469 7389 9503
rect 7423 9500 7435 9503
rect 7466 9500 7472 9512
rect 7423 9472 7472 9500
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 7558 9460 7564 9512
rect 7616 9500 7622 9512
rect 7837 9503 7895 9509
rect 7837 9500 7849 9503
rect 7616 9472 7849 9500
rect 7616 9460 7622 9472
rect 7837 9469 7849 9472
rect 7883 9469 7895 9503
rect 7837 9463 7895 9469
rect 7926 9460 7932 9512
rect 7984 9460 7990 9512
rect 8128 9509 8156 9608
rect 8754 9596 8760 9648
rect 8812 9636 8818 9648
rect 8812 9608 10824 9636
rect 8812 9596 8818 9608
rect 9122 9528 9128 9580
rect 9180 9528 9186 9580
rect 8113 9503 8171 9509
rect 8113 9469 8125 9503
rect 8159 9500 8171 9503
rect 9140 9500 9168 9528
rect 9401 9503 9459 9509
rect 9401 9500 9413 9503
rect 8159 9472 8984 9500
rect 9140 9472 9413 9500
rect 8159 9469 8171 9472
rect 8113 9463 8171 9469
rect 7009 9435 7067 9441
rect 7009 9401 7021 9435
rect 7055 9401 7067 9435
rect 7009 9395 7067 9401
rect 4955 9336 5488 9364
rect 4955 9333 4967 9336
rect 4909 9327 4967 9333
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 5905 9367 5963 9373
rect 5905 9364 5917 9367
rect 5592 9336 5917 9364
rect 5592 9324 5598 9336
rect 5905 9333 5917 9336
rect 5951 9333 5963 9367
rect 5905 9327 5963 9333
rect 6270 9324 6276 9376
rect 6328 9324 6334 9376
rect 6546 9324 6552 9376
rect 6604 9364 6610 9376
rect 6733 9367 6791 9373
rect 6733 9364 6745 9367
rect 6604 9336 6745 9364
rect 6604 9324 6610 9336
rect 6733 9333 6745 9336
rect 6779 9333 6791 9367
rect 7024 9364 7052 9395
rect 7190 9392 7196 9444
rect 7248 9441 7254 9444
rect 7248 9435 7297 9441
rect 7248 9401 7251 9435
rect 7285 9432 7297 9435
rect 7650 9432 7656 9444
rect 7285 9404 7656 9432
rect 7285 9401 7297 9404
rect 7248 9395 7297 9401
rect 7248 9392 7254 9395
rect 7650 9392 7656 9404
rect 7708 9392 7714 9444
rect 8389 9435 8447 9441
rect 8389 9401 8401 9435
rect 8435 9432 8447 9435
rect 8849 9435 8907 9441
rect 8849 9432 8861 9435
rect 8435 9404 8861 9432
rect 8435 9401 8447 9404
rect 8389 9395 8447 9401
rect 8849 9401 8861 9404
rect 8895 9401 8907 9435
rect 8956 9432 8984 9472
rect 9401 9469 9413 9472
rect 9447 9469 9459 9503
rect 9401 9463 9459 9469
rect 9490 9460 9496 9512
rect 9548 9460 9554 9512
rect 9049 9435 9107 9441
rect 9049 9432 9061 9435
rect 8956 9404 9061 9432
rect 8849 9395 8907 9401
rect 9049 9401 9061 9404
rect 9095 9401 9107 9435
rect 9508 9432 9536 9460
rect 10796 9444 10824 9608
rect 11026 9568 11054 9676
rect 12529 9673 12541 9676
rect 12575 9673 12587 9707
rect 12529 9667 12587 9673
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 12492 9608 13124 9636
rect 12492 9596 12498 9608
rect 13096 9577 13124 9608
rect 10980 9540 11054 9568
rect 13081 9571 13139 9577
rect 10980 9509 11008 9540
rect 13081 9537 13093 9571
rect 13127 9537 13139 9571
rect 13081 9531 13139 9537
rect 14090 9528 14096 9580
rect 14148 9528 14154 9580
rect 10965 9503 11023 9509
rect 10965 9469 10977 9503
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 11057 9503 11115 9509
rect 11057 9469 11069 9503
rect 11103 9500 11115 9503
rect 12986 9500 12992 9512
rect 11103 9472 12992 9500
rect 11103 9469 11115 9472
rect 11057 9463 11115 9469
rect 12986 9460 12992 9472
rect 13044 9460 13050 9512
rect 14369 9503 14427 9509
rect 14369 9469 14381 9503
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 9049 9395 9107 9401
rect 9140 9404 9536 9432
rect 7469 9367 7527 9373
rect 7469 9364 7481 9367
rect 7024 9336 7481 9364
rect 6733 9327 6791 9333
rect 7469 9333 7481 9336
rect 7515 9333 7527 9367
rect 7469 9327 7527 9333
rect 7558 9324 7564 9376
rect 7616 9364 7622 9376
rect 8589 9367 8647 9373
rect 8589 9364 8601 9367
rect 7616 9336 8601 9364
rect 7616 9324 7622 9336
rect 8589 9333 8601 9336
rect 8635 9333 8647 9367
rect 8864 9364 8892 9395
rect 9140 9364 9168 9404
rect 10778 9392 10784 9444
rect 10836 9432 10842 9444
rect 11324 9435 11382 9441
rect 10836 9404 11008 9432
rect 10836 9392 10842 9404
rect 8864 9336 9168 9364
rect 8589 9327 8647 9333
rect 9214 9324 9220 9376
rect 9272 9324 9278 9376
rect 9677 9367 9735 9373
rect 9677 9333 9689 9367
rect 9723 9364 9735 9367
rect 10594 9364 10600 9376
rect 9723 9336 10600 9364
rect 9723 9333 9735 9336
rect 9677 9327 9735 9333
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 10870 9324 10876 9376
rect 10928 9324 10934 9376
rect 10980 9364 11008 9404
rect 11324 9401 11336 9435
rect 11370 9432 11382 9435
rect 11422 9432 11428 9444
rect 11370 9404 11428 9432
rect 11370 9401 11382 9404
rect 11324 9395 11382 9401
rect 11422 9392 11428 9404
rect 11480 9392 11486 9444
rect 12250 9392 12256 9444
rect 12308 9432 12314 9444
rect 13909 9435 13967 9441
rect 13909 9432 13921 9435
rect 12308 9404 13921 9432
rect 12308 9392 12314 9404
rect 13909 9401 13921 9404
rect 13955 9401 13967 9435
rect 13909 9395 13967 9401
rect 14274 9392 14280 9444
rect 14332 9432 14338 9444
rect 14384 9432 14412 9463
rect 14550 9460 14556 9512
rect 14608 9460 14614 9512
rect 14332 9404 14412 9432
rect 14568 9432 14596 9460
rect 15010 9432 15016 9444
rect 14568 9404 15016 9432
rect 14332 9392 14338 9404
rect 15010 9392 15016 9404
rect 15068 9392 15074 9444
rect 11514 9364 11520 9376
rect 10980 9336 11520 9364
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 13541 9367 13599 9373
rect 13541 9364 13553 9367
rect 13136 9336 13553 9364
rect 13136 9324 13142 9336
rect 13541 9333 13553 9336
rect 13587 9333 13599 9367
rect 13541 9327 13599 9333
rect 14001 9367 14059 9373
rect 14001 9333 14013 9367
rect 14047 9364 14059 9367
rect 14461 9367 14519 9373
rect 14461 9364 14473 9367
rect 14047 9336 14473 9364
rect 14047 9333 14059 9336
rect 14001 9327 14059 9333
rect 14461 9333 14473 9336
rect 14507 9333 14519 9367
rect 14461 9327 14519 9333
rect 552 9274 15520 9296
rect 552 9222 4100 9274
rect 4152 9222 4164 9274
rect 4216 9222 4228 9274
rect 4280 9222 4292 9274
rect 4344 9222 4356 9274
rect 4408 9222 7802 9274
rect 7854 9222 7866 9274
rect 7918 9222 7930 9274
rect 7982 9222 7994 9274
rect 8046 9222 8058 9274
rect 8110 9222 11504 9274
rect 11556 9222 11568 9274
rect 11620 9222 11632 9274
rect 11684 9222 11696 9274
rect 11748 9222 11760 9274
rect 11812 9222 15206 9274
rect 15258 9222 15270 9274
rect 15322 9222 15334 9274
rect 15386 9222 15398 9274
rect 15450 9222 15462 9274
rect 15514 9222 15520 9274
rect 552 9200 15520 9222
rect 3234 9120 3240 9172
rect 3292 9120 3298 9172
rect 3326 9120 3332 9172
rect 3384 9120 3390 9172
rect 3510 9120 3516 9172
rect 3568 9160 3574 9172
rect 3973 9163 4031 9169
rect 3973 9160 3985 9163
rect 3568 9132 3985 9160
rect 3568 9120 3574 9132
rect 3973 9129 3985 9132
rect 4019 9129 4031 9163
rect 3973 9123 4031 9129
rect 4614 9120 4620 9172
rect 4672 9120 4678 9172
rect 4890 9120 4896 9172
rect 4948 9120 4954 9172
rect 7190 9120 7196 9172
rect 7248 9120 7254 9172
rect 8386 9120 8392 9172
rect 8444 9160 8450 9172
rect 8573 9163 8631 9169
rect 8573 9160 8585 9163
rect 8444 9132 8585 9160
rect 8444 9120 8450 9132
rect 8573 9129 8585 9132
rect 8619 9129 8631 9163
rect 8573 9123 8631 9129
rect 9214 9120 9220 9172
rect 9272 9120 9278 9172
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 10042 9160 10048 9172
rect 9364 9132 10048 9160
rect 9364 9120 9370 9132
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 10597 9163 10655 9169
rect 10597 9129 10609 9163
rect 10643 9160 10655 9163
rect 10686 9160 10692 9172
rect 10643 9132 10692 9160
rect 10643 9129 10655 9132
rect 10597 9123 10655 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 11422 9120 11428 9172
rect 11480 9160 11486 9172
rect 11701 9163 11759 9169
rect 11701 9160 11713 9163
rect 11480 9132 11713 9160
rect 11480 9120 11486 9132
rect 11701 9129 11713 9132
rect 11747 9129 11759 9163
rect 12894 9160 12900 9172
rect 11701 9123 11759 9129
rect 12268 9132 12900 9160
rect 3252 9033 3280 9120
rect 3237 9027 3295 9033
rect 3237 8993 3249 9027
rect 3283 8993 3295 9027
rect 3237 8987 3295 8993
rect 3421 9027 3479 9033
rect 3421 8993 3433 9027
rect 3467 9024 3479 9027
rect 3602 9024 3608 9036
rect 3467 8996 3608 9024
rect 3467 8993 3479 8996
rect 3421 8987 3479 8993
rect 3602 8984 3608 8996
rect 3660 8984 3666 9036
rect 3881 9027 3939 9033
rect 3881 8993 3893 9027
rect 3927 9024 3939 9027
rect 3970 9024 3976 9036
rect 3927 8996 3976 9024
rect 3927 8993 3939 8996
rect 3881 8987 3939 8993
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 9024 4123 9027
rect 4430 9024 4436 9036
rect 4111 8996 4436 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 4632 9024 4660 9120
rect 5534 9092 5540 9104
rect 4908 9064 5540 9092
rect 4801 9027 4859 9033
rect 4801 9024 4813 9027
rect 4632 8996 4813 9024
rect 4801 8993 4813 8996
rect 4847 8993 4859 9027
rect 4801 8987 4859 8993
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8956 2651 8959
rect 2866 8956 2872 8968
rect 2639 8928 2872 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3786 8916 3792 8968
rect 3844 8956 3850 8968
rect 4908 8956 4936 9064
rect 5534 9052 5540 9064
rect 5592 9052 5598 9104
rect 6080 9095 6138 9101
rect 6080 9061 6092 9095
rect 6126 9092 6138 9095
rect 6270 9092 6276 9104
rect 6126 9064 6276 9092
rect 6126 9061 6138 9064
rect 6080 9055 6138 9061
rect 6270 9052 6276 9064
rect 6328 9052 6334 9104
rect 7282 9052 7288 9104
rect 7340 9052 7346 9104
rect 9232 9092 9260 9120
rect 9140 9064 9260 9092
rect 9140 9033 9168 9064
rect 9125 9027 9183 9033
rect 9125 8993 9137 9027
rect 9171 8993 9183 9027
rect 9125 8987 9183 8993
rect 9217 9027 9275 9033
rect 9217 8993 9229 9027
rect 9263 9024 9275 9027
rect 9324 9024 9352 9120
rect 9585 9095 9643 9101
rect 9585 9061 9597 9095
rect 9631 9092 9643 9095
rect 10226 9092 10232 9104
rect 9631 9064 9904 9092
rect 9631 9061 9643 9064
rect 9585 9055 9643 9061
rect 9263 8996 9352 9024
rect 9401 9027 9459 9033
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 9401 8993 9413 9027
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 3844 8928 4936 8956
rect 3844 8916 3850 8928
rect 5810 8916 5816 8968
rect 5868 8916 5874 8968
rect 9416 8956 9444 8987
rect 9674 8984 9680 9036
rect 9732 8984 9738 9036
rect 9876 9033 9904 9064
rect 10060 9064 10232 9092
rect 9861 9027 9919 9033
rect 9861 8993 9873 9027
rect 9907 8993 9919 9027
rect 9861 8987 9919 8993
rect 9950 8984 9956 9036
rect 10008 8984 10014 9036
rect 10060 9033 10088 9064
rect 10226 9052 10232 9064
rect 10284 9092 10290 9104
rect 12268 9092 12296 9132
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 13078 9120 13084 9172
rect 13136 9120 13142 9172
rect 14550 9160 14556 9172
rect 13188 9132 14556 9160
rect 13096 9092 13124 9120
rect 10284 9064 12296 9092
rect 10284 9052 10290 9064
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 10413 9027 10471 9033
rect 10413 8993 10425 9027
rect 10459 9024 10471 9027
rect 10594 9024 10600 9036
rect 10459 8996 10600 9024
rect 10459 8993 10471 8996
rect 10413 8987 10471 8993
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 10689 9027 10747 9033
rect 10689 8993 10701 9027
rect 10735 9024 10747 9027
rect 10778 9024 10784 9036
rect 10735 8996 10784 9024
rect 10735 8993 10747 8996
rect 10689 8987 10747 8993
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 11885 9027 11943 9033
rect 11885 9024 11897 9027
rect 10928 8996 11897 9024
rect 10928 8984 10934 8996
rect 11885 8993 11897 8996
rect 11931 8993 11943 9027
rect 11885 8987 11943 8993
rect 11974 8984 11980 9036
rect 12032 9024 12038 9036
rect 12161 9027 12219 9033
rect 12161 9024 12173 9027
rect 12032 8996 12173 9024
rect 12032 8984 12038 8996
rect 12161 8993 12173 8996
rect 12207 8993 12219 9027
rect 12161 8987 12219 8993
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 9324 8928 9444 8956
rect 9784 8928 10977 8956
rect 3694 8848 3700 8900
rect 3752 8888 3758 8900
rect 5718 8888 5724 8900
rect 3752 8860 5724 8888
rect 3752 8848 3758 8860
rect 5718 8848 5724 8860
rect 5776 8848 5782 8900
rect 1946 8780 1952 8832
rect 2004 8780 2010 8832
rect 5074 8780 5080 8832
rect 5132 8820 5138 8832
rect 7558 8820 7564 8832
rect 5132 8792 7564 8820
rect 5132 8780 5138 8792
rect 7558 8780 7564 8792
rect 7616 8820 7622 8832
rect 9122 8820 9128 8832
rect 7616 8792 9128 8820
rect 7616 8780 7622 8792
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 9324 8820 9352 8928
rect 9784 8820 9812 8928
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8925 11575 8959
rect 12268 8956 12296 9064
rect 12728 9064 13124 9092
rect 12345 9027 12403 9033
rect 12345 8993 12357 9027
rect 12391 9024 12403 9027
rect 12434 9024 12440 9036
rect 12391 8996 12440 9024
rect 12391 8993 12403 8996
rect 12345 8987 12403 8993
rect 12434 8984 12440 8996
rect 12492 9024 12498 9036
rect 12529 9027 12587 9033
rect 12529 9024 12541 9027
rect 12492 8996 12541 9024
rect 12492 8984 12498 8996
rect 12529 8993 12541 8996
rect 12575 8993 12587 9027
rect 12529 8987 12587 8993
rect 11517 8919 11575 8925
rect 11992 8928 12296 8956
rect 9950 8848 9956 8900
rect 10008 8888 10014 8900
rect 10008 8860 10456 8888
rect 10008 8848 10014 8860
rect 9324 8792 9812 8820
rect 10134 8780 10140 8832
rect 10192 8820 10198 8832
rect 10428 8829 10456 8860
rect 10686 8848 10692 8900
rect 10744 8888 10750 8900
rect 11238 8888 11244 8900
rect 10744 8860 11244 8888
rect 10744 8848 10750 8860
rect 11238 8848 11244 8860
rect 11296 8888 11302 8900
rect 11532 8888 11560 8919
rect 11992 8897 12020 8928
rect 11296 8860 11560 8888
rect 11977 8891 12035 8897
rect 11296 8848 11302 8860
rect 11977 8857 11989 8891
rect 12023 8857 12035 8891
rect 11977 8851 12035 8857
rect 12069 8891 12127 8897
rect 12069 8857 12081 8891
rect 12115 8857 12127 8891
rect 12069 8851 12127 8857
rect 10321 8823 10379 8829
rect 10321 8820 10333 8823
rect 10192 8792 10333 8820
rect 10192 8780 10198 8792
rect 10321 8789 10333 8792
rect 10367 8789 10379 8823
rect 10321 8783 10379 8789
rect 10413 8823 10471 8829
rect 10413 8789 10425 8823
rect 10459 8820 10471 8823
rect 12084 8820 12112 8851
rect 10459 8792 12112 8820
rect 12544 8820 12572 8987
rect 12618 8984 12624 9036
rect 12676 8984 12682 9036
rect 12728 9033 12756 9064
rect 12713 9027 12771 9033
rect 12713 8993 12725 9027
rect 12759 8993 12771 9027
rect 12713 8987 12771 8993
rect 13081 9027 13139 9033
rect 13081 8993 13093 9027
rect 13127 9024 13139 9027
rect 13188 9024 13216 9132
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 13127 8996 13216 9024
rect 13265 9027 13323 9033
rect 13127 8993 13139 8996
rect 13081 8987 13139 8993
rect 13265 8993 13277 9027
rect 13311 9024 13323 9027
rect 13633 9027 13691 9033
rect 13633 9024 13645 9027
rect 13311 8996 13645 9024
rect 13311 8993 13323 8996
rect 13265 8987 13323 8993
rect 13633 8993 13645 8996
rect 13679 8993 13691 9027
rect 13633 8987 13691 8993
rect 12636 8956 12664 8984
rect 12805 8959 12863 8965
rect 12805 8956 12817 8959
rect 12636 8928 12817 8956
rect 12805 8925 12817 8928
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 12894 8916 12900 8968
rect 12952 8916 12958 8968
rect 12986 8916 12992 8968
rect 13044 8956 13050 8968
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 13044 8928 13369 8956
rect 13044 8916 13050 8928
rect 13357 8925 13369 8928
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 14090 8820 14096 8832
rect 12544 8792 14096 8820
rect 10459 8789 10471 8792
rect 10413 8783 10471 8789
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 14921 8823 14979 8829
rect 14921 8789 14933 8823
rect 14967 8820 14979 8823
rect 15010 8820 15016 8832
rect 14967 8792 15016 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15010 8780 15016 8792
rect 15068 8780 15074 8832
rect 552 8730 15364 8752
rect 552 8678 2249 8730
rect 2301 8678 2313 8730
rect 2365 8678 2377 8730
rect 2429 8678 2441 8730
rect 2493 8678 2505 8730
rect 2557 8678 5951 8730
rect 6003 8678 6015 8730
rect 6067 8678 6079 8730
rect 6131 8678 6143 8730
rect 6195 8678 6207 8730
rect 6259 8678 9653 8730
rect 9705 8678 9717 8730
rect 9769 8678 9781 8730
rect 9833 8678 9845 8730
rect 9897 8678 9909 8730
rect 9961 8678 13355 8730
rect 13407 8678 13419 8730
rect 13471 8678 13483 8730
rect 13535 8678 13547 8730
rect 13599 8678 13611 8730
rect 13663 8678 15364 8730
rect 552 8656 15364 8678
rect 2866 8576 2872 8628
rect 2924 8576 2930 8628
rect 4433 8619 4491 8625
rect 4433 8585 4445 8619
rect 4479 8616 4491 8619
rect 5169 8619 5227 8625
rect 4479 8588 5120 8616
rect 4479 8585 4491 8588
rect 4433 8579 4491 8585
rect 3237 8551 3295 8557
rect 3237 8517 3249 8551
rect 3283 8517 3295 8551
rect 3237 8511 3295 8517
rect 3973 8551 4031 8557
rect 3973 8517 3985 8551
rect 4019 8517 4031 8551
rect 3973 8511 4031 8517
rect 1486 8372 1492 8424
rect 1544 8412 1550 8424
rect 2682 8412 2688 8424
rect 1544 8384 2688 8412
rect 1544 8372 1550 8384
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 3252 8412 3280 8511
rect 2976 8384 3280 8412
rect 3513 8415 3571 8421
rect 1756 8347 1814 8353
rect 1756 8313 1768 8347
rect 1802 8344 1814 8347
rect 2976 8344 3004 8384
rect 3513 8381 3525 8415
rect 3559 8412 3571 8415
rect 3988 8412 4016 8511
rect 4062 8508 4068 8560
rect 4120 8548 4126 8560
rect 4617 8551 4675 8557
rect 4617 8548 4629 8551
rect 4120 8520 4629 8548
rect 4120 8508 4126 8520
rect 4617 8517 4629 8520
rect 4663 8517 4675 8551
rect 5092 8548 5120 8588
rect 5169 8585 5181 8619
rect 5215 8616 5227 8619
rect 5258 8616 5264 8628
rect 5215 8588 5264 8616
rect 5215 8585 5227 8588
rect 5169 8579 5227 8585
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 6273 8619 6331 8625
rect 6273 8585 6285 8619
rect 6319 8616 6331 8619
rect 6454 8616 6460 8628
rect 6319 8588 6460 8616
rect 6319 8585 6331 8588
rect 6273 8579 6331 8585
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 11238 8576 11244 8628
rect 11296 8576 11302 8628
rect 12894 8576 12900 8628
rect 12952 8616 12958 8628
rect 13173 8619 13231 8625
rect 13173 8616 13185 8619
rect 12952 8588 13185 8616
rect 12952 8576 12958 8588
rect 13173 8585 13185 8588
rect 13219 8585 13231 8619
rect 13173 8579 13231 8585
rect 5626 8548 5632 8560
rect 5092 8520 5632 8548
rect 4617 8511 4675 8517
rect 5626 8508 5632 8520
rect 5684 8508 5690 8560
rect 8665 8551 8723 8557
rect 8665 8517 8677 8551
rect 8711 8548 8723 8551
rect 9401 8551 9459 8557
rect 9401 8548 9413 8551
rect 8711 8520 9413 8548
rect 8711 8517 8723 8520
rect 8665 8511 8723 8517
rect 9401 8517 9413 8520
rect 9447 8517 9459 8551
rect 9401 8511 9459 8517
rect 12342 8508 12348 8560
rect 12400 8548 12406 8560
rect 12400 8520 13768 8548
rect 12400 8508 12406 8520
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8480 4307 8483
rect 4430 8480 4436 8492
rect 4295 8452 4436 8480
rect 4295 8449 4307 8452
rect 4249 8443 4307 8449
rect 4430 8440 4436 8452
rect 4488 8440 4494 8492
rect 6362 8440 6368 8492
rect 6420 8480 6426 8492
rect 6641 8483 6699 8489
rect 6641 8480 6653 8483
rect 6420 8452 6653 8480
rect 6420 8440 6426 8452
rect 6641 8449 6653 8452
rect 6687 8449 6699 8483
rect 9214 8480 9220 8492
rect 6641 8443 6699 8449
rect 7392 8452 9220 8480
rect 7392 8424 7420 8452
rect 9214 8440 9220 8452
rect 9272 8480 9278 8492
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 9272 8452 9873 8480
rect 9272 8440 9278 8452
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 13633 8483 13691 8489
rect 13633 8480 13645 8483
rect 9861 8443 9919 8449
rect 13188 8452 13645 8480
rect 13188 8424 13216 8452
rect 13633 8449 13645 8452
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 3559 8384 4016 8412
rect 3559 8381 3571 8384
rect 3513 8375 3571 8381
rect 4522 8372 4528 8424
rect 4580 8372 4586 8424
rect 4798 8372 4804 8424
rect 4856 8412 4862 8424
rect 4985 8415 5043 8421
rect 4985 8412 4997 8415
rect 4856 8384 4997 8412
rect 4856 8372 4862 8384
rect 4985 8381 4997 8384
rect 5031 8381 5043 8415
rect 4985 8375 5043 8381
rect 5166 8372 5172 8424
rect 5224 8412 5230 8424
rect 5445 8415 5503 8421
rect 5445 8412 5457 8415
rect 5224 8384 5457 8412
rect 5224 8372 5230 8384
rect 5445 8381 5457 8384
rect 5491 8381 5503 8415
rect 5445 8375 5503 8381
rect 6457 8415 6515 8421
rect 6457 8381 6469 8415
rect 6503 8412 6515 8415
rect 6546 8412 6552 8424
rect 6503 8384 6552 8412
rect 6503 8381 6515 8384
rect 6457 8375 6515 8381
rect 6546 8372 6552 8384
rect 6604 8372 6610 8424
rect 7374 8372 7380 8424
rect 7432 8372 7438 8424
rect 8573 8415 8631 8421
rect 8573 8412 8585 8415
rect 8496 8384 8585 8412
rect 1802 8316 3004 8344
rect 1802 8313 1814 8316
rect 1756 8307 1814 8313
rect 3142 8304 3148 8356
rect 3200 8344 3206 8356
rect 3237 8347 3295 8353
rect 3237 8344 3249 8347
rect 3200 8316 3249 8344
rect 3200 8304 3206 8316
rect 3237 8313 3249 8316
rect 3283 8344 3295 8347
rect 3694 8344 3700 8356
rect 3283 8316 3700 8344
rect 3283 8313 3295 8316
rect 3237 8307 3295 8313
rect 3694 8304 3700 8316
rect 3752 8304 3758 8356
rect 3786 8304 3792 8356
rect 3844 8344 3850 8356
rect 3844 8316 5534 8344
rect 3844 8304 3850 8316
rect 3418 8236 3424 8288
rect 3476 8236 3482 8288
rect 4706 8236 4712 8288
rect 4764 8276 4770 8288
rect 4801 8279 4859 8285
rect 4801 8276 4813 8279
rect 4764 8248 4813 8276
rect 4764 8236 4770 8248
rect 4801 8245 4813 8248
rect 4847 8245 4859 8279
rect 4801 8239 4859 8245
rect 4890 8236 4896 8288
rect 4948 8236 4954 8288
rect 5506 8276 5534 8316
rect 8496 8288 8524 8384
rect 8573 8381 8585 8384
rect 8619 8381 8631 8415
rect 8573 8375 8631 8381
rect 8754 8372 8760 8424
rect 8812 8372 8818 8424
rect 8846 8372 8852 8424
rect 8904 8372 8910 8424
rect 8938 8372 8944 8424
rect 8996 8412 9002 8424
rect 9033 8415 9091 8421
rect 9033 8412 9045 8415
rect 8996 8384 9045 8412
rect 8996 8372 9002 8384
rect 9033 8381 9045 8384
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 9048 8344 9076 8375
rect 9122 8372 9128 8424
rect 9180 8372 9186 8424
rect 10134 8421 10140 8424
rect 9585 8415 9643 8421
rect 9585 8412 9597 8415
rect 9232 8384 9597 8412
rect 9232 8344 9260 8384
rect 9585 8381 9597 8384
rect 9631 8381 9643 8415
rect 9585 8375 9643 8381
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8381 9735 8415
rect 10128 8412 10140 8421
rect 10095 8384 10140 8412
rect 9677 8375 9735 8381
rect 10128 8375 10140 8384
rect 9048 8316 9260 8344
rect 9401 8347 9459 8353
rect 9401 8313 9413 8347
rect 9447 8344 9459 8347
rect 9490 8344 9496 8356
rect 9447 8316 9496 8344
rect 9447 8313 9459 8316
rect 9401 8307 9459 8313
rect 9490 8304 9496 8316
rect 9548 8344 9554 8356
rect 9692 8344 9720 8375
rect 10134 8372 10140 8375
rect 10192 8372 10198 8424
rect 12618 8372 12624 8424
rect 12676 8372 12682 8424
rect 13170 8372 13176 8424
rect 13228 8372 13234 8424
rect 13740 8421 13768 8520
rect 13357 8415 13415 8421
rect 13357 8381 13369 8415
rect 13403 8381 13415 8415
rect 13357 8375 13415 8381
rect 13541 8415 13599 8421
rect 13541 8381 13553 8415
rect 13587 8381 13599 8415
rect 13541 8375 13599 8381
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 9548 8316 9720 8344
rect 12636 8344 12664 8372
rect 13372 8344 13400 8375
rect 12636 8316 13400 8344
rect 13556 8344 13584 8375
rect 14274 8372 14280 8424
rect 14332 8372 14338 8424
rect 14292 8344 14320 8372
rect 13556 8316 14320 8344
rect 9548 8304 9554 8316
rect 5626 8276 5632 8288
rect 5506 8248 5632 8276
rect 5626 8236 5632 8248
rect 5684 8236 5690 8288
rect 8202 8236 8208 8288
rect 8260 8276 8266 8288
rect 8389 8279 8447 8285
rect 8389 8276 8401 8279
rect 8260 8248 8401 8276
rect 8260 8236 8266 8248
rect 8389 8245 8401 8248
rect 8435 8245 8447 8279
rect 8389 8239 8447 8245
rect 8478 8236 8484 8288
rect 8536 8236 8542 8288
rect 9030 8236 9036 8288
rect 9088 8276 9094 8288
rect 9217 8279 9275 8285
rect 9217 8276 9229 8279
rect 9088 8248 9229 8276
rect 9088 8236 9094 8248
rect 9217 8245 9229 8248
rect 9263 8245 9275 8279
rect 9217 8239 9275 8245
rect 11974 8236 11980 8288
rect 12032 8276 12038 8288
rect 13906 8276 13912 8288
rect 12032 8248 13912 8276
rect 12032 8236 12038 8248
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 552 8186 15520 8208
rect 552 8134 4100 8186
rect 4152 8134 4164 8186
rect 4216 8134 4228 8186
rect 4280 8134 4292 8186
rect 4344 8134 4356 8186
rect 4408 8134 7802 8186
rect 7854 8134 7866 8186
rect 7918 8134 7930 8186
rect 7982 8134 7994 8186
rect 8046 8134 8058 8186
rect 8110 8134 11504 8186
rect 11556 8134 11568 8186
rect 11620 8134 11632 8186
rect 11684 8134 11696 8186
rect 11748 8134 11760 8186
rect 11812 8134 15206 8186
rect 15258 8134 15270 8186
rect 15322 8134 15334 8186
rect 15386 8134 15398 8186
rect 15450 8134 15462 8186
rect 15514 8134 15520 8186
rect 552 8112 15520 8134
rect 1946 8032 1952 8084
rect 2004 8032 2010 8084
rect 2501 8075 2559 8081
rect 2501 8041 2513 8075
rect 2547 8072 2559 8075
rect 3418 8072 3424 8084
rect 2547 8044 3424 8072
rect 2547 8041 2559 8044
rect 2501 8035 2559 8041
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 9490 8072 9496 8084
rect 8803 8044 9496 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 10226 8032 10232 8084
rect 10284 8032 10290 8084
rect 10410 8032 10416 8084
rect 10468 8072 10474 8084
rect 10468 8044 13400 8072
rect 10468 8032 10474 8044
rect 1964 7936 1992 8032
rect 2774 8004 2780 8016
rect 2516 7976 2780 8004
rect 2516 7945 2544 7976
rect 2774 7964 2780 7976
rect 2832 7964 2838 8016
rect 4341 8007 4399 8013
rect 4341 7973 4353 8007
rect 4387 8004 4399 8007
rect 4982 8004 4988 8016
rect 4387 7976 4988 8004
rect 4387 7973 4399 7976
rect 4341 7967 4399 7973
rect 4982 7964 4988 7976
rect 5040 7964 5046 8016
rect 5626 7964 5632 8016
rect 5684 8004 5690 8016
rect 5684 7976 9076 8004
rect 5684 7964 5690 7976
rect 9048 7948 9076 7976
rect 2317 7939 2375 7945
rect 2317 7936 2329 7939
rect 1964 7908 2329 7936
rect 2317 7905 2329 7908
rect 2363 7905 2375 7939
rect 2317 7899 2375 7905
rect 2501 7939 2559 7945
rect 2501 7905 2513 7939
rect 2547 7905 2559 7939
rect 2501 7899 2559 7905
rect 4706 7896 4712 7948
rect 4764 7896 4770 7948
rect 7374 7896 7380 7948
rect 7432 7896 7438 7948
rect 7650 7945 7656 7948
rect 7644 7899 7656 7945
rect 7650 7896 7656 7899
rect 7708 7896 7714 7948
rect 8570 7896 8576 7948
rect 8628 7936 8634 7948
rect 8849 7939 8907 7945
rect 8849 7936 8861 7939
rect 8628 7908 8861 7936
rect 8628 7896 8634 7908
rect 8849 7905 8861 7908
rect 8895 7905 8907 7939
rect 8849 7899 8907 7905
rect 9030 7896 9036 7948
rect 9088 7936 9094 7948
rect 10244 7936 10272 8032
rect 12066 7964 12072 8016
rect 12124 7964 12130 8016
rect 12618 7964 12624 8016
rect 12676 8004 12682 8016
rect 12676 7976 12940 8004
rect 12676 7964 12682 7976
rect 9088 7908 10272 7936
rect 9088 7896 9094 7908
rect 10594 7896 10600 7948
rect 10652 7936 10658 7948
rect 11330 7936 11336 7948
rect 10652 7908 11336 7936
rect 10652 7896 10658 7908
rect 11330 7896 11336 7908
rect 11388 7936 11394 7948
rect 11974 7936 11980 7948
rect 11388 7908 11980 7936
rect 11388 7896 11394 7908
rect 11974 7896 11980 7908
rect 12032 7896 12038 7948
rect 12084 7936 12112 7964
rect 12084 7908 12388 7936
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 4525 7871 4583 7877
rect 4525 7868 4537 7871
rect 4120 7840 4537 7868
rect 4120 7828 4126 7840
rect 4525 7837 4537 7840
rect 4571 7837 4583 7871
rect 4525 7831 4583 7837
rect 4614 7828 4620 7880
rect 4672 7828 4678 7880
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7868 4859 7871
rect 4890 7868 4896 7880
rect 4847 7840 4896 7868
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 11882 7828 11888 7880
rect 11940 7828 11946 7880
rect 12069 7871 12127 7877
rect 12069 7837 12081 7871
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 12161 7871 12219 7877
rect 12161 7837 12173 7871
rect 12207 7837 12219 7871
rect 12360 7868 12388 7908
rect 12526 7896 12532 7948
rect 12584 7936 12590 7948
rect 12912 7945 12940 7976
rect 13170 7964 13176 8016
rect 13228 7964 13234 8016
rect 13078 7945 13084 7948
rect 12805 7939 12863 7945
rect 12805 7936 12817 7939
rect 12584 7908 12817 7936
rect 12584 7896 12590 7908
rect 12805 7905 12817 7908
rect 12851 7905 12863 7939
rect 12805 7899 12863 7905
rect 12897 7939 12955 7945
rect 12897 7905 12909 7939
rect 12943 7905 12955 7939
rect 12897 7899 12955 7905
rect 13045 7939 13084 7945
rect 13045 7905 13057 7939
rect 13045 7899 13084 7905
rect 13078 7896 13084 7899
rect 13136 7896 13142 7948
rect 13372 7945 13400 8044
rect 13265 7939 13323 7945
rect 13265 7905 13277 7939
rect 13311 7905 13323 7939
rect 13265 7899 13323 7905
rect 13362 7939 13420 7945
rect 13362 7905 13374 7939
rect 13408 7905 13420 7939
rect 13362 7899 13420 7905
rect 12710 7868 12716 7880
rect 12360 7840 12716 7868
rect 12161 7831 12219 7837
rect 2682 7760 2688 7812
rect 2740 7800 2746 7812
rect 3053 7803 3111 7809
rect 3053 7800 3065 7803
rect 2740 7772 3065 7800
rect 2740 7760 2746 7772
rect 3053 7769 3065 7772
rect 3099 7800 3111 7803
rect 3326 7800 3332 7812
rect 3099 7772 3332 7800
rect 3099 7769 3111 7772
rect 3053 7763 3111 7769
rect 3326 7760 3332 7772
rect 3384 7800 3390 7812
rect 5810 7800 5816 7812
rect 3384 7772 5816 7800
rect 3384 7760 3390 7772
rect 5810 7760 5816 7772
rect 5868 7760 5874 7812
rect 8941 7803 8999 7809
rect 8941 7769 8953 7803
rect 8987 7800 8999 7803
rect 12084 7800 12112 7831
rect 8987 7772 12112 7800
rect 12176 7800 12204 7831
rect 12710 7828 12716 7840
rect 12768 7828 12774 7880
rect 13280 7868 13308 7899
rect 12820 7840 13308 7868
rect 12820 7812 12848 7840
rect 12437 7803 12495 7809
rect 12437 7800 12449 7803
rect 12176 7772 12449 7800
rect 8987 7769 8999 7772
rect 8941 7763 8999 7769
rect 12437 7769 12449 7772
rect 12483 7769 12495 7803
rect 12437 7763 12495 7769
rect 12802 7760 12808 7812
rect 12860 7760 12866 7812
rect 4522 7692 4528 7744
rect 4580 7732 4586 7744
rect 4985 7735 5043 7741
rect 4985 7732 4997 7735
rect 4580 7704 4997 7732
rect 4580 7692 4586 7704
rect 4985 7701 4997 7704
rect 5031 7701 5043 7735
rect 4985 7695 5043 7701
rect 9306 7692 9312 7744
rect 9364 7732 9370 7744
rect 10226 7732 10232 7744
rect 9364 7704 10232 7732
rect 9364 7692 9370 7704
rect 10226 7692 10232 7704
rect 10284 7692 10290 7744
rect 12342 7692 12348 7744
rect 12400 7692 12406 7744
rect 12618 7692 12624 7744
rect 12676 7692 12682 7744
rect 13541 7735 13599 7741
rect 13541 7701 13553 7735
rect 13587 7732 13599 7735
rect 13998 7732 14004 7744
rect 13587 7704 14004 7732
rect 13587 7701 13599 7704
rect 13541 7695 13599 7701
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 552 7642 15364 7664
rect 552 7590 2249 7642
rect 2301 7590 2313 7642
rect 2365 7590 2377 7642
rect 2429 7590 2441 7642
rect 2493 7590 2505 7642
rect 2557 7590 5951 7642
rect 6003 7590 6015 7642
rect 6067 7590 6079 7642
rect 6131 7590 6143 7642
rect 6195 7590 6207 7642
rect 6259 7590 9653 7642
rect 9705 7590 9717 7642
rect 9769 7590 9781 7642
rect 9833 7590 9845 7642
rect 9897 7590 9909 7642
rect 9961 7590 13355 7642
rect 13407 7590 13419 7642
rect 13471 7590 13483 7642
rect 13535 7590 13547 7642
rect 13599 7590 13611 7642
rect 13663 7590 15364 7642
rect 552 7568 15364 7590
rect 4341 7531 4399 7537
rect 4341 7497 4353 7531
rect 4387 7528 4399 7531
rect 4430 7528 4436 7540
rect 4387 7500 4436 7528
rect 4387 7497 4399 7500
rect 4341 7491 4399 7497
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 4798 7488 4804 7540
rect 4856 7488 4862 7540
rect 7650 7488 7656 7540
rect 7708 7528 7714 7540
rect 7837 7531 7895 7537
rect 7837 7528 7849 7531
rect 7708 7500 7849 7528
rect 7708 7488 7714 7500
rect 7837 7497 7849 7500
rect 7883 7497 7895 7531
rect 10962 7528 10968 7540
rect 7837 7491 7895 7497
rect 9600 7500 10968 7528
rect 2866 7420 2872 7472
rect 2924 7460 2930 7472
rect 3789 7463 3847 7469
rect 3789 7460 3801 7463
rect 2924 7432 3801 7460
rect 2924 7420 2930 7432
rect 3789 7429 3801 7432
rect 3835 7429 3847 7463
rect 3789 7423 3847 7429
rect 3804 7392 3832 7423
rect 6362 7420 6368 7472
rect 6420 7460 6426 7472
rect 6420 7432 6868 7460
rect 6420 7420 6426 7432
rect 4062 7392 4068 7404
rect 3804 7364 4068 7392
rect 4062 7352 4068 7364
rect 4120 7392 4126 7404
rect 6840 7401 6868 7432
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 4120 7364 4445 7392
rect 4120 7352 4126 7364
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 7469 7395 7527 7401
rect 7469 7361 7481 7395
rect 7515 7392 7527 7395
rect 9600 7392 9628 7500
rect 10962 7488 10968 7500
rect 11020 7528 11026 7540
rect 11425 7531 11483 7537
rect 11425 7528 11437 7531
rect 11020 7500 11437 7528
rect 11020 7488 11026 7500
rect 11425 7497 11437 7500
rect 11471 7497 11483 7531
rect 11425 7491 11483 7497
rect 12161 7531 12219 7537
rect 12161 7497 12173 7531
rect 12207 7528 12219 7531
rect 12250 7528 12256 7540
rect 12207 7500 12256 7528
rect 12207 7497 12219 7500
rect 12161 7491 12219 7497
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 13078 7488 13084 7540
rect 13136 7528 13142 7540
rect 13265 7531 13323 7537
rect 13265 7528 13277 7531
rect 13136 7500 13277 7528
rect 13136 7488 13142 7500
rect 13265 7497 13277 7500
rect 13311 7497 13323 7531
rect 13265 7491 13323 7497
rect 9677 7463 9735 7469
rect 9677 7429 9689 7463
rect 9723 7460 9735 7463
rect 9861 7463 9919 7469
rect 9861 7460 9873 7463
rect 9723 7432 9873 7460
rect 9723 7429 9735 7432
rect 9677 7423 9735 7429
rect 9861 7429 9873 7432
rect 9907 7429 9919 7463
rect 9861 7423 9919 7429
rect 7515 7364 7972 7392
rect 9600 7364 9720 7392
rect 7515 7361 7527 7364
rect 7469 7355 7527 7361
rect 4614 7324 4620 7336
rect 3988 7296 4620 7324
rect 2866 7148 2872 7200
rect 2924 7188 2930 7200
rect 3878 7188 3884 7200
rect 2924 7160 3884 7188
rect 2924 7148 2930 7160
rect 3878 7148 3884 7160
rect 3936 7188 3942 7200
rect 3988 7197 4016 7296
rect 4614 7284 4620 7296
rect 4672 7284 4678 7336
rect 4706 7284 4712 7336
rect 4764 7284 4770 7336
rect 4985 7327 5043 7333
rect 4985 7293 4997 7327
rect 5031 7324 5043 7327
rect 5810 7324 5816 7336
rect 5031 7296 5816 7324
rect 5031 7293 5043 7296
rect 4985 7287 5043 7293
rect 5810 7284 5816 7296
rect 5868 7284 5874 7336
rect 7653 7327 7711 7333
rect 7653 7293 7665 7327
rect 7699 7324 7711 7327
rect 7742 7324 7748 7336
rect 7699 7296 7748 7324
rect 7699 7293 7711 7296
rect 7653 7287 7711 7293
rect 4065 7259 4123 7265
rect 4065 7225 4077 7259
rect 4111 7256 4123 7259
rect 4724 7256 4752 7284
rect 4111 7228 4752 7256
rect 5252 7259 5310 7265
rect 4111 7225 4123 7228
rect 4065 7219 4123 7225
rect 5252 7225 5264 7259
rect 5298 7256 5310 7259
rect 5350 7256 5356 7268
rect 5298 7228 5356 7256
rect 5298 7225 5310 7228
rect 5252 7219 5310 7225
rect 5350 7216 5356 7228
rect 5408 7216 5414 7268
rect 7466 7216 7472 7268
rect 7524 7256 7530 7268
rect 7668 7256 7696 7287
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 7944 7333 7972 7364
rect 7837 7327 7895 7333
rect 7837 7293 7849 7327
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7293 7987 7327
rect 7929 7287 7987 7293
rect 7524 7228 7696 7256
rect 7852 7256 7880 7287
rect 8202 7284 8208 7336
rect 8260 7284 8266 7336
rect 9398 7284 9404 7336
rect 9456 7284 9462 7336
rect 9692 7333 9720 7364
rect 9677 7327 9735 7333
rect 9677 7293 9689 7327
rect 9723 7293 9735 7327
rect 9677 7287 9735 7293
rect 9769 7327 9827 7333
rect 9769 7293 9781 7327
rect 9815 7293 9827 7327
rect 9876 7324 9904 7423
rect 10134 7420 10140 7472
rect 10192 7420 10198 7472
rect 10226 7420 10232 7472
rect 10284 7420 10290 7472
rect 12268 7460 12296 7488
rect 11164 7432 11744 7460
rect 12268 7432 12664 7460
rect 10045 7395 10103 7401
rect 10045 7361 10057 7395
rect 10091 7392 10103 7395
rect 10244 7392 10272 7420
rect 10091 7364 10272 7392
rect 10091 7361 10103 7364
rect 10045 7355 10103 7361
rect 10413 7327 10471 7333
rect 10413 7324 10425 7327
rect 9876 7296 10425 7324
rect 9769 7287 9827 7293
rect 10413 7293 10425 7296
rect 10459 7293 10471 7327
rect 10413 7287 10471 7293
rect 8220 7256 8248 7284
rect 7852 7228 8248 7256
rect 7524 7216 7530 7228
rect 3973 7191 4031 7197
rect 3973 7188 3985 7191
rect 3936 7160 3985 7188
rect 3936 7148 3942 7160
rect 3973 7157 3985 7160
rect 4019 7157 4031 7191
rect 3973 7151 4031 7157
rect 4157 7191 4215 7197
rect 4157 7157 4169 7191
rect 4203 7188 4215 7191
rect 4522 7188 4528 7200
rect 4203 7160 4528 7188
rect 4203 7157 4215 7160
rect 4157 7151 4215 7157
rect 4522 7148 4528 7160
rect 4580 7188 4586 7200
rect 4890 7188 4896 7200
rect 4580 7160 4896 7188
rect 4580 7148 4586 7160
rect 4890 7148 4896 7160
rect 4948 7148 4954 7200
rect 7558 7148 7564 7200
rect 7616 7188 7622 7200
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 7616 7160 8033 7188
rect 7616 7148 7622 7160
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 8021 7151 8079 7157
rect 9490 7148 9496 7200
rect 9548 7148 9554 7200
rect 9784 7188 9812 7287
rect 10502 7284 10508 7336
rect 10560 7324 10566 7336
rect 11164 7333 11192 7432
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 10560 7296 10977 7324
rect 10560 7284 10566 7296
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 10965 7287 11023 7293
rect 11149 7327 11207 7333
rect 11149 7293 11161 7327
rect 11195 7293 11207 7327
rect 11149 7287 11207 7293
rect 11333 7327 11391 7333
rect 11333 7293 11345 7327
rect 11379 7324 11391 7327
rect 11422 7324 11428 7336
rect 11379 7296 11428 7324
rect 11379 7293 11391 7296
rect 11333 7287 11391 7293
rect 11422 7284 11428 7296
rect 11480 7284 11486 7336
rect 11609 7327 11667 7333
rect 11609 7293 11621 7327
rect 11655 7293 11667 7327
rect 11716 7324 11744 7432
rect 12529 7395 12587 7401
rect 12529 7392 12541 7395
rect 12084 7364 12541 7392
rect 12084 7324 12112 7364
rect 12529 7361 12541 7364
rect 12575 7361 12587 7395
rect 12529 7355 12587 7361
rect 11716 7296 12112 7324
rect 12253 7327 12311 7333
rect 11609 7287 11667 7293
rect 12253 7293 12265 7327
rect 12299 7324 12311 7327
rect 12299 7296 12388 7324
rect 12299 7293 12311 7296
rect 12253 7287 12311 7293
rect 10045 7259 10103 7265
rect 10045 7225 10057 7259
rect 10091 7256 10103 7259
rect 10137 7259 10195 7265
rect 10137 7256 10149 7259
rect 10091 7228 10149 7256
rect 10091 7225 10103 7228
rect 10045 7219 10103 7225
rect 10137 7225 10149 7228
rect 10183 7225 10195 7259
rect 10137 7219 10195 7225
rect 10321 7259 10379 7265
rect 10321 7225 10333 7259
rect 10367 7256 10379 7259
rect 10594 7256 10600 7268
rect 10367 7228 10600 7256
rect 10367 7225 10379 7228
rect 10321 7219 10379 7225
rect 10336 7188 10364 7219
rect 10594 7216 10600 7228
rect 10652 7216 10658 7268
rect 11054 7216 11060 7268
rect 11112 7256 11118 7268
rect 11624 7256 11652 7287
rect 11112 7228 12296 7256
rect 11112 7216 11118 7228
rect 12268 7200 12296 7228
rect 9784 7160 10364 7188
rect 10781 7191 10839 7197
rect 10781 7157 10793 7191
rect 10827 7188 10839 7191
rect 11238 7188 11244 7200
rect 10827 7160 11244 7188
rect 10827 7157 10839 7160
rect 10781 7151 10839 7157
rect 11238 7148 11244 7160
rect 11296 7148 11302 7200
rect 12250 7148 12256 7200
rect 12308 7148 12314 7200
rect 12360 7188 12388 7296
rect 12434 7284 12440 7336
rect 12492 7284 12498 7336
rect 12636 7333 12664 7432
rect 13832 7364 15056 7392
rect 13832 7333 13860 7364
rect 15028 7336 15056 7364
rect 12621 7327 12679 7333
rect 12621 7293 12633 7327
rect 12667 7293 12679 7327
rect 12621 7287 12679 7293
rect 13081 7327 13139 7333
rect 13081 7293 13093 7327
rect 13127 7324 13139 7327
rect 13817 7327 13875 7333
rect 13817 7324 13829 7327
rect 13127 7296 13829 7324
rect 13127 7293 13139 7296
rect 13081 7287 13139 7293
rect 13817 7293 13829 7296
rect 13863 7293 13875 7327
rect 13817 7287 13875 7293
rect 13906 7284 13912 7336
rect 13964 7284 13970 7336
rect 13998 7284 14004 7336
rect 14056 7284 14062 7336
rect 14182 7284 14188 7336
rect 14240 7284 14246 7336
rect 15010 7284 15016 7336
rect 15068 7284 15074 7336
rect 12526 7216 12532 7268
rect 12584 7256 12590 7268
rect 12897 7259 12955 7265
rect 12897 7256 12909 7259
rect 12584 7228 12909 7256
rect 12584 7216 12590 7228
rect 12897 7225 12909 7228
rect 12943 7225 12955 7259
rect 12897 7219 12955 7225
rect 12710 7188 12716 7200
rect 12360 7160 12716 7188
rect 12710 7148 12716 7160
rect 12768 7148 12774 7200
rect 13541 7191 13599 7197
rect 13541 7157 13553 7191
rect 13587 7188 13599 7191
rect 13630 7188 13636 7200
rect 13587 7160 13636 7188
rect 13587 7157 13599 7160
rect 13541 7151 13599 7157
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 552 7098 15520 7120
rect 552 7046 4100 7098
rect 4152 7046 4164 7098
rect 4216 7046 4228 7098
rect 4280 7046 4292 7098
rect 4344 7046 4356 7098
rect 4408 7046 7802 7098
rect 7854 7046 7866 7098
rect 7918 7046 7930 7098
rect 7982 7046 7994 7098
rect 8046 7046 8058 7098
rect 8110 7046 11504 7098
rect 11556 7046 11568 7098
rect 11620 7046 11632 7098
rect 11684 7046 11696 7098
rect 11748 7046 11760 7098
rect 11812 7046 15206 7098
rect 15258 7046 15270 7098
rect 15322 7046 15334 7098
rect 15386 7046 15398 7098
rect 15450 7046 15462 7098
rect 15514 7046 15520 7098
rect 552 7024 15520 7046
rect 2961 6987 3019 6993
rect 2961 6984 2973 6987
rect 2884 6956 2973 6984
rect 2884 6928 2912 6956
rect 2961 6953 2973 6956
rect 3007 6953 3019 6987
rect 2961 6947 3019 6953
rect 3602 6944 3608 6996
rect 3660 6984 3666 6996
rect 3660 6956 4844 6984
rect 3660 6944 3666 6956
rect 2866 6876 2872 6928
rect 2924 6876 2930 6928
rect 4706 6916 4712 6928
rect 4172 6888 4712 6916
rect 2774 6808 2780 6860
rect 2832 6848 2838 6860
rect 2958 6851 3016 6857
rect 2958 6848 2970 6851
rect 2832 6820 2970 6848
rect 2832 6808 2838 6820
rect 2958 6817 2970 6820
rect 3004 6848 3016 6851
rect 3786 6848 3792 6860
rect 3004 6820 3792 6848
rect 3004 6817 3016 6820
rect 2958 6811 3016 6817
rect 3786 6808 3792 6820
rect 3844 6808 3850 6860
rect 3878 6808 3884 6860
rect 3936 6857 3942 6860
rect 4172 6857 4200 6888
rect 4706 6876 4712 6888
rect 4764 6876 4770 6928
rect 3936 6848 3946 6857
rect 4157 6851 4215 6857
rect 3936 6820 3977 6848
rect 3936 6811 3946 6820
rect 4157 6817 4169 6851
rect 4203 6817 4215 6851
rect 4157 6811 4215 6817
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6848 4399 6851
rect 4816 6848 4844 6956
rect 5350 6944 5356 6996
rect 5408 6944 5414 6996
rect 7558 6944 7564 6996
rect 7616 6944 7622 6996
rect 7650 6944 7656 6996
rect 7708 6984 7714 6996
rect 9490 6984 9496 6996
rect 7708 6956 9496 6984
rect 7708 6944 7714 6956
rect 9490 6944 9496 6956
rect 9548 6984 9554 6996
rect 11054 6984 11060 6996
rect 9548 6956 11060 6984
rect 9548 6944 9554 6956
rect 11054 6944 11060 6956
rect 11112 6944 11118 6996
rect 12069 6987 12127 6993
rect 12069 6953 12081 6987
rect 12115 6984 12127 6987
rect 12434 6984 12440 6996
rect 12115 6956 12440 6984
rect 12115 6953 12127 6956
rect 12069 6947 12127 6953
rect 12434 6944 12440 6956
rect 12492 6944 12498 6996
rect 12526 6944 12532 6996
rect 12584 6944 12590 6996
rect 12912 6956 14504 6984
rect 5261 6851 5319 6857
rect 5261 6848 5273 6851
rect 4387 6820 4568 6848
rect 4816 6820 5273 6848
rect 4387 6817 4399 6820
rect 4341 6811 4399 6817
rect 3936 6808 3942 6811
rect 4540 6792 4568 6820
rect 5261 6817 5273 6820
rect 5307 6817 5319 6851
rect 5261 6811 5319 6817
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6817 5503 6851
rect 5445 6811 5503 6817
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6780 4031 6783
rect 4019 6752 4292 6780
rect 4019 6749 4031 6752
rect 3973 6743 4031 6749
rect 3436 6712 3464 6743
rect 3436 6684 4200 6712
rect 4172 6656 4200 6684
rect 2774 6604 2780 6656
rect 2832 6604 2838 6656
rect 3329 6647 3387 6653
rect 3329 6613 3341 6647
rect 3375 6644 3387 6647
rect 3513 6647 3571 6653
rect 3513 6644 3525 6647
rect 3375 6616 3525 6644
rect 3375 6613 3387 6616
rect 3329 6607 3387 6613
rect 3513 6613 3525 6616
rect 3559 6613 3571 6647
rect 3513 6607 3571 6613
rect 4154 6604 4160 6656
rect 4212 6604 4218 6656
rect 4264 6653 4292 6752
rect 4522 6740 4528 6792
rect 4580 6740 4586 6792
rect 5460 6712 5488 6811
rect 5810 6808 5816 6860
rect 5868 6848 5874 6860
rect 6181 6851 6239 6857
rect 6181 6848 6193 6851
rect 5868 6820 6193 6848
rect 5868 6808 5874 6820
rect 6181 6817 6193 6820
rect 6227 6817 6239 6851
rect 6181 6811 6239 6817
rect 6362 6808 6368 6860
rect 6420 6808 6426 6860
rect 6638 6808 6644 6860
rect 6696 6848 6702 6860
rect 7101 6851 7159 6857
rect 6696 6820 7052 6848
rect 6696 6808 6702 6820
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6780 6331 6783
rect 6825 6783 6883 6789
rect 6825 6780 6837 6783
rect 6319 6752 6837 6780
rect 6319 6749 6331 6752
rect 6273 6743 6331 6749
rect 6825 6749 6837 6752
rect 6871 6749 6883 6783
rect 6825 6743 6883 6749
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6749 6975 6783
rect 7024 6780 7052 6820
rect 7101 6817 7113 6851
rect 7147 6848 7159 6851
rect 7576 6848 7604 6944
rect 11422 6876 11428 6928
rect 11480 6916 11486 6928
rect 12912 6925 12940 6956
rect 14476 6928 14504 6956
rect 12681 6919 12739 6925
rect 12681 6916 12693 6919
rect 11480 6888 12693 6916
rect 11480 6876 11486 6888
rect 7147 6820 7604 6848
rect 7147 6817 7159 6820
rect 7101 6811 7159 6817
rect 8478 6808 8484 6860
rect 8536 6808 8542 6860
rect 11992 6857 12020 6888
rect 12681 6885 12693 6888
rect 12727 6885 12739 6919
rect 12681 6879 12739 6885
rect 12897 6919 12955 6925
rect 12897 6885 12909 6919
rect 12943 6885 12955 6919
rect 12897 6879 12955 6885
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 11935 6820 11989 6848
rect 11977 6817 11989 6820
rect 12023 6817 12035 6851
rect 11977 6811 12035 6817
rect 12253 6851 12311 6857
rect 12253 6817 12265 6851
rect 12299 6848 12311 6851
rect 12912 6848 12940 6879
rect 14458 6876 14464 6928
rect 14516 6876 14522 6928
rect 12299 6820 12940 6848
rect 12299 6817 12311 6820
rect 12253 6811 12311 6817
rect 8496 6780 8524 6808
rect 7024 6752 8524 6780
rect 11992 6780 12020 6811
rect 12986 6808 12992 6860
rect 13044 6848 13050 6860
rect 13357 6851 13415 6857
rect 13357 6848 13369 6851
rect 13044 6820 13369 6848
rect 13044 6808 13050 6820
rect 13357 6817 13369 6820
rect 13403 6817 13415 6851
rect 13357 6811 13415 6817
rect 13630 6808 13636 6860
rect 13688 6808 13694 6860
rect 15010 6808 15016 6860
rect 15068 6808 15074 6860
rect 11992 6752 12848 6780
rect 6917 6743 6975 6749
rect 6457 6715 6515 6721
rect 6457 6712 6469 6715
rect 5460 6684 6469 6712
rect 6457 6681 6469 6684
rect 6503 6681 6515 6715
rect 6457 6675 6515 6681
rect 6730 6672 6736 6724
rect 6788 6672 6794 6724
rect 6932 6712 6960 6743
rect 8846 6712 8852 6724
rect 6932 6684 8852 6712
rect 4249 6647 4307 6653
rect 4249 6613 4261 6647
rect 4295 6644 4307 6647
rect 4430 6644 4436 6656
rect 4295 6616 4436 6644
rect 4295 6613 4307 6616
rect 4249 6607 4307 6613
rect 4430 6604 4436 6616
rect 4488 6604 4494 6656
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 6270 6644 6276 6656
rect 5776 6616 6276 6644
rect 5776 6604 5782 6616
rect 6270 6604 6276 6616
rect 6328 6644 6334 6656
rect 6932 6644 6960 6684
rect 8846 6672 8852 6684
rect 8904 6672 8910 6724
rect 12253 6715 12311 6721
rect 12253 6681 12265 6715
rect 12299 6712 12311 6715
rect 12618 6712 12624 6724
rect 12299 6684 12624 6712
rect 12299 6681 12311 6684
rect 12253 6675 12311 6681
rect 12618 6672 12624 6684
rect 12676 6672 12682 6724
rect 12820 6656 12848 6752
rect 6328 6616 6960 6644
rect 6328 6604 6334 6616
rect 12710 6604 12716 6656
rect 12768 6604 12774 6656
rect 12802 6604 12808 6656
rect 12860 6604 12866 6656
rect 552 6554 15364 6576
rect 552 6502 2249 6554
rect 2301 6502 2313 6554
rect 2365 6502 2377 6554
rect 2429 6502 2441 6554
rect 2493 6502 2505 6554
rect 2557 6502 5951 6554
rect 6003 6502 6015 6554
rect 6067 6502 6079 6554
rect 6131 6502 6143 6554
rect 6195 6502 6207 6554
rect 6259 6502 9653 6554
rect 9705 6502 9717 6554
rect 9769 6502 9781 6554
rect 9833 6502 9845 6554
rect 9897 6502 9909 6554
rect 9961 6502 13355 6554
rect 13407 6502 13419 6554
rect 13471 6502 13483 6554
rect 13535 6502 13547 6554
rect 13599 6502 13611 6554
rect 13663 6502 15364 6554
rect 552 6480 15364 6502
rect 2774 6400 2780 6452
rect 2832 6400 2838 6452
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4341 6443 4399 6449
rect 4341 6440 4353 6443
rect 4212 6412 4353 6440
rect 4212 6400 4218 6412
rect 4341 6409 4353 6412
rect 4387 6409 4399 6443
rect 4341 6403 4399 6409
rect 1394 6264 1400 6316
rect 1452 6264 1458 6316
rect 2792 6236 2820 6400
rect 4356 6372 4384 6403
rect 4522 6400 4528 6452
rect 4580 6440 4586 6452
rect 6730 6440 6736 6452
rect 4580 6412 6736 6440
rect 4580 6400 4586 6412
rect 6730 6400 6736 6412
rect 6788 6440 6794 6452
rect 7009 6443 7067 6449
rect 7009 6440 7021 6443
rect 6788 6412 7021 6440
rect 6788 6400 6794 6412
rect 7009 6409 7021 6412
rect 7055 6409 7067 6443
rect 7009 6403 7067 6409
rect 9677 6443 9735 6449
rect 9677 6409 9689 6443
rect 9723 6440 9735 6443
rect 10042 6440 10048 6452
rect 9723 6412 10048 6440
rect 9723 6409 9735 6412
rect 9677 6403 9735 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10962 6400 10968 6452
rect 11020 6400 11026 6452
rect 14274 6400 14280 6452
rect 14332 6400 14338 6452
rect 5534 6372 5540 6384
rect 4356 6344 5540 6372
rect 5506 6332 5540 6344
rect 5592 6332 5598 6384
rect 6362 6332 6368 6384
rect 6420 6372 6426 6384
rect 6457 6375 6515 6381
rect 6457 6372 6469 6375
rect 6420 6344 6469 6372
rect 6420 6332 6426 6344
rect 6457 6341 6469 6344
rect 6503 6341 6515 6375
rect 6457 6335 6515 6341
rect 6638 6332 6644 6384
rect 6696 6332 6702 6384
rect 8113 6375 8171 6381
rect 8113 6341 8125 6375
rect 8159 6372 8171 6375
rect 8481 6375 8539 6381
rect 8481 6372 8493 6375
rect 8159 6344 8493 6372
rect 8159 6341 8171 6344
rect 8113 6335 8171 6341
rect 8481 6341 8493 6344
rect 8527 6341 8539 6375
rect 8481 6335 8539 6341
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 9861 6375 9919 6381
rect 9861 6372 9873 6375
rect 9824 6344 9873 6372
rect 9824 6332 9830 6344
rect 9861 6341 9873 6344
rect 9907 6341 9919 6375
rect 9861 6335 9919 6341
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4617 6307 4675 6313
rect 4617 6304 4629 6307
rect 4203 6276 4629 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 4617 6273 4629 6276
rect 4663 6273 4675 6307
rect 5506 6304 5534 6332
rect 6656 6304 6684 6332
rect 5506 6276 6684 6304
rect 4617 6267 4675 6273
rect 2869 6239 2927 6245
rect 2869 6236 2881 6239
rect 2792 6208 2881 6236
rect 2869 6205 2881 6208
rect 2915 6205 2927 6239
rect 2869 6199 2927 6205
rect 3053 6239 3111 6245
rect 3053 6205 3065 6239
rect 3099 6236 3111 6239
rect 3602 6236 3608 6248
rect 3099 6208 3608 6236
rect 3099 6205 3111 6208
rect 3053 6199 3111 6205
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 4430 6196 4436 6248
rect 4488 6196 4494 6248
rect 4522 6196 4528 6248
rect 4580 6196 4586 6248
rect 4706 6196 4712 6248
rect 4764 6196 4770 6248
rect 5920 6245 5948 6276
rect 7834 6264 7840 6316
rect 7892 6304 7898 6316
rect 10060 6304 10088 6400
rect 10226 6332 10232 6384
rect 10284 6372 10290 6384
rect 12066 6372 12072 6384
rect 10284 6344 12072 6372
rect 10284 6332 10290 6344
rect 12066 6332 12072 6344
rect 12124 6332 12130 6384
rect 12434 6332 12440 6384
rect 12492 6332 12498 6384
rect 14829 6375 14887 6381
rect 14829 6341 14841 6375
rect 14875 6372 14887 6375
rect 15010 6372 15016 6384
rect 14875 6344 15016 6372
rect 14875 6341 14887 6344
rect 14829 6335 14887 6341
rect 15010 6332 15016 6344
rect 15068 6332 15074 6384
rect 11149 6307 11207 6313
rect 7892 6276 9444 6304
rect 10060 6276 10916 6304
rect 7892 6264 7898 6276
rect 5905 6239 5963 6245
rect 5905 6205 5917 6239
rect 5951 6205 5963 6239
rect 5905 6199 5963 6205
rect 5994 6196 6000 6248
rect 6052 6196 6058 6248
rect 6086 6196 6092 6248
rect 6144 6196 6150 6248
rect 6181 6239 6239 6245
rect 6181 6205 6193 6239
rect 6227 6236 6239 6239
rect 6270 6236 6276 6248
rect 6227 6208 6276 6236
rect 6227 6205 6239 6208
rect 6181 6199 6239 6205
rect 6270 6196 6276 6208
rect 6328 6196 6334 6248
rect 6365 6239 6423 6245
rect 6365 6205 6377 6239
rect 6411 6236 6423 6239
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 6411 6208 7297 6236
rect 6411 6205 6423 6208
rect 6365 6199 6423 6205
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 7374 6196 7380 6248
rect 7432 6196 7438 6248
rect 7745 6239 7803 6245
rect 7745 6205 7757 6239
rect 7791 6205 7803 6239
rect 7745 6199 7803 6205
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 8478 6236 8484 6248
rect 8435 6208 8484 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 1664 6171 1722 6177
rect 1664 6137 1676 6171
rect 1710 6168 1722 6171
rect 2961 6171 3019 6177
rect 2961 6168 2973 6171
rect 1710 6140 2973 6168
rect 1710 6137 1722 6140
rect 1664 6131 1722 6137
rect 2961 6137 2973 6140
rect 3007 6137 3019 6171
rect 2961 6131 3019 6137
rect 6730 6128 6736 6180
rect 6788 6168 6794 6180
rect 7760 6168 7788 6199
rect 8478 6196 8484 6208
rect 8536 6196 8542 6248
rect 8908 6239 8966 6245
rect 8908 6205 8920 6239
rect 8954 6236 8966 6239
rect 9030 6236 9036 6248
rect 8954 6208 9036 6236
rect 8954 6205 8966 6208
rect 8908 6199 8966 6205
rect 9030 6196 9036 6208
rect 9088 6196 9094 6248
rect 6788 6140 8892 6168
rect 6788 6128 6794 6140
rect 2777 6103 2835 6109
rect 2777 6069 2789 6103
rect 2823 6100 2835 6103
rect 2866 6100 2872 6112
rect 2823 6072 2872 6100
rect 2823 6069 2835 6072
rect 2777 6063 2835 6069
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 3878 6060 3884 6112
rect 3936 6060 3942 6112
rect 5718 6060 5724 6112
rect 5776 6060 5782 6112
rect 6638 6060 6644 6112
rect 6696 6060 6702 6112
rect 6822 6060 6828 6112
rect 6880 6100 6886 6112
rect 7834 6100 7840 6112
rect 6880 6072 7840 6100
rect 6880 6060 6886 6072
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8864 6109 8892 6140
rect 8849 6103 8907 6109
rect 8849 6069 8861 6103
rect 8895 6069 8907 6103
rect 8849 6063 8907 6069
rect 9030 6060 9036 6112
rect 9088 6060 9094 6112
rect 9122 6060 9128 6112
rect 9180 6100 9186 6112
rect 9309 6103 9367 6109
rect 9309 6100 9321 6103
rect 9180 6072 9321 6100
rect 9180 6060 9186 6072
rect 9309 6069 9321 6072
rect 9355 6069 9367 6103
rect 9416 6100 9444 6276
rect 9493 6239 9551 6245
rect 9493 6205 9505 6239
rect 9539 6236 9551 6239
rect 9674 6236 9680 6248
rect 9539 6208 9680 6236
rect 9539 6205 9551 6208
rect 9493 6199 9551 6205
rect 9674 6196 9680 6208
rect 9732 6196 9738 6248
rect 9766 6196 9772 6248
rect 9824 6196 9830 6248
rect 10042 6196 10048 6248
rect 10100 6196 10106 6248
rect 10888 6245 10916 6276
rect 11149 6273 11161 6307
rect 11195 6304 11207 6307
rect 12452 6304 12480 6332
rect 11195 6276 12480 6304
rect 11195 6273 11207 6276
rect 11149 6267 11207 6273
rect 10137 6239 10195 6245
rect 10137 6205 10149 6239
rect 10183 6236 10195 6239
rect 10873 6239 10931 6245
rect 10183 6208 10364 6236
rect 10183 6205 10195 6208
rect 10137 6199 10195 6205
rect 9861 6171 9919 6177
rect 9861 6137 9873 6171
rect 9907 6168 9919 6171
rect 10226 6168 10232 6180
rect 9907 6140 10232 6168
rect 9907 6137 9919 6140
rect 9861 6131 9919 6137
rect 10226 6128 10232 6140
rect 10284 6128 10290 6180
rect 10336 6112 10364 6208
rect 10873 6205 10885 6239
rect 10919 6205 10931 6239
rect 10873 6199 10931 6205
rect 11238 6196 11244 6248
rect 11296 6196 11302 6248
rect 11422 6196 11428 6248
rect 11480 6196 11486 6248
rect 12342 6196 12348 6248
rect 12400 6236 12406 6248
rect 12713 6239 12771 6245
rect 12713 6236 12725 6239
rect 12400 6208 12725 6236
rect 12400 6196 12406 6208
rect 12713 6205 12725 6208
rect 12759 6205 12771 6239
rect 12713 6199 12771 6205
rect 12989 6239 13047 6245
rect 12989 6205 13001 6239
rect 13035 6205 13047 6239
rect 12989 6199 13047 6205
rect 13173 6239 13231 6245
rect 13173 6205 13185 6239
rect 13219 6236 13231 6239
rect 13541 6239 13599 6245
rect 13541 6236 13553 6239
rect 13219 6208 13553 6236
rect 13219 6205 13231 6208
rect 13173 6199 13231 6205
rect 13541 6205 13553 6208
rect 13587 6205 13599 6239
rect 13541 6199 13599 6205
rect 14185 6239 14243 6245
rect 14185 6205 14197 6239
rect 14231 6236 14243 6239
rect 14458 6236 14464 6248
rect 14231 6208 14464 6236
rect 14231 6205 14243 6208
rect 14185 6199 14243 6205
rect 11440 6168 11468 6196
rect 13004 6168 13032 6199
rect 14458 6196 14464 6208
rect 14516 6236 14522 6248
rect 14645 6239 14703 6245
rect 14645 6236 14657 6239
rect 14516 6208 14657 6236
rect 14516 6196 14522 6208
rect 14645 6205 14657 6208
rect 14691 6205 14703 6239
rect 14645 6199 14703 6205
rect 11440 6140 13032 6168
rect 10318 6100 10324 6112
rect 9416 6072 10324 6100
rect 9309 6063 9367 6069
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 11146 6060 11152 6112
rect 11204 6060 11210 6112
rect 11330 6060 11336 6112
rect 11388 6060 11394 6112
rect 12526 6060 12532 6112
rect 12584 6060 12590 6112
rect 12802 6060 12808 6112
rect 12860 6100 12866 6112
rect 14461 6103 14519 6109
rect 14461 6100 14473 6103
rect 12860 6072 14473 6100
rect 12860 6060 12866 6072
rect 14461 6069 14473 6072
rect 14507 6069 14519 6103
rect 14461 6063 14519 6069
rect 14550 6060 14556 6112
rect 14608 6060 14614 6112
rect 552 6010 15520 6032
rect 552 5958 4100 6010
rect 4152 5958 4164 6010
rect 4216 5958 4228 6010
rect 4280 5958 4292 6010
rect 4344 5958 4356 6010
rect 4408 5958 7802 6010
rect 7854 5958 7866 6010
rect 7918 5958 7930 6010
rect 7982 5958 7994 6010
rect 8046 5958 8058 6010
rect 8110 5958 11504 6010
rect 11556 5958 11568 6010
rect 11620 5958 11632 6010
rect 11684 5958 11696 6010
rect 11748 5958 11760 6010
rect 11812 5958 15206 6010
rect 15258 5958 15270 6010
rect 15322 5958 15334 6010
rect 15386 5958 15398 6010
rect 15450 5958 15462 6010
rect 15514 5958 15520 6010
rect 552 5936 15520 5958
rect 3878 5856 3884 5908
rect 3936 5856 3942 5908
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4028 5868 4108 5896
rect 4028 5856 4034 5868
rect 3694 5788 3700 5840
rect 3752 5788 3758 5840
rect 3896 5828 3924 5856
rect 3896 5800 4016 5828
rect 3602 5720 3608 5772
rect 3660 5720 3666 5772
rect 3988 5769 4016 5800
rect 4080 5769 4108 5868
rect 5994 5856 6000 5908
rect 6052 5896 6058 5908
rect 6546 5905 6552 5908
rect 6365 5899 6423 5905
rect 6365 5896 6377 5899
rect 6052 5868 6377 5896
rect 6052 5856 6058 5868
rect 6365 5865 6377 5868
rect 6411 5865 6423 5899
rect 6365 5859 6423 5865
rect 6528 5899 6552 5905
rect 6528 5865 6540 5899
rect 6604 5896 6610 5908
rect 6822 5896 6828 5908
rect 6604 5868 6828 5896
rect 6528 5859 6552 5865
rect 6546 5856 6552 5859
rect 6604 5856 6610 5868
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 7469 5899 7527 5905
rect 7469 5896 7481 5899
rect 7432 5868 7481 5896
rect 7432 5856 7438 5868
rect 7469 5865 7481 5868
rect 7515 5865 7527 5899
rect 7469 5859 7527 5865
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5896 9183 5899
rect 9214 5896 9220 5908
rect 9171 5868 9220 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 9766 5856 9772 5908
rect 9824 5896 9830 5908
rect 10045 5899 10103 5905
rect 10045 5896 10057 5899
rect 9824 5868 10057 5896
rect 9824 5856 9830 5868
rect 10045 5865 10057 5868
rect 10091 5865 10103 5899
rect 10045 5859 10103 5865
rect 11330 5856 11336 5908
rect 11388 5856 11394 5908
rect 12158 5856 12164 5908
rect 12216 5856 12222 5908
rect 6733 5831 6791 5837
rect 6012 5800 6500 5828
rect 6012 5772 6040 5800
rect 3881 5763 3939 5769
rect 3881 5729 3893 5763
rect 3927 5729 3939 5763
rect 3881 5723 3939 5729
rect 3973 5763 4031 5769
rect 3973 5729 3985 5763
rect 4019 5729 4031 5763
rect 3973 5723 4031 5729
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5729 4123 5763
rect 4065 5723 4123 5729
rect 4249 5763 4307 5769
rect 4249 5729 4261 5763
rect 4295 5760 4307 5763
rect 4525 5763 4583 5769
rect 4525 5760 4537 5763
rect 4295 5732 4537 5760
rect 4295 5729 4307 5732
rect 4249 5723 4307 5729
rect 4525 5729 4537 5732
rect 4571 5729 4583 5763
rect 4525 5723 4583 5729
rect 3620 5624 3648 5720
rect 3896 5692 3924 5723
rect 4706 5720 4712 5772
rect 4764 5760 4770 5772
rect 5077 5763 5135 5769
rect 5077 5760 5089 5763
rect 4764 5732 5089 5760
rect 4764 5720 4770 5732
rect 5077 5729 5089 5732
rect 5123 5729 5135 5763
rect 5261 5763 5319 5769
rect 5261 5760 5273 5763
rect 5077 5723 5135 5729
rect 5184 5732 5273 5760
rect 4157 5695 4215 5701
rect 4157 5692 4169 5695
rect 3896 5664 4169 5692
rect 4157 5661 4169 5664
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 5184 5624 5212 5732
rect 5261 5729 5273 5732
rect 5307 5729 5319 5763
rect 5261 5723 5319 5729
rect 5445 5763 5503 5769
rect 5445 5729 5457 5763
rect 5491 5760 5503 5763
rect 5718 5760 5724 5772
rect 5491 5732 5724 5760
rect 5491 5729 5503 5732
rect 5445 5723 5503 5729
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 5994 5720 6000 5772
rect 6052 5720 6058 5772
rect 6181 5763 6239 5769
rect 6181 5729 6193 5763
rect 6227 5729 6239 5763
rect 6181 5723 6239 5729
rect 6273 5763 6331 5769
rect 6273 5729 6285 5763
rect 6319 5760 6331 5763
rect 6362 5760 6368 5772
rect 6319 5732 6368 5760
rect 6319 5729 6331 5732
rect 6273 5723 6331 5729
rect 6086 5652 6092 5704
rect 6144 5652 6150 5704
rect 6196 5692 6224 5723
rect 6362 5720 6368 5732
rect 6420 5720 6426 5772
rect 6472 5760 6500 5800
rect 6733 5797 6745 5831
rect 6779 5797 6791 5831
rect 6733 5791 6791 5797
rect 7837 5831 7895 5837
rect 7837 5797 7849 5831
rect 7883 5828 7895 5831
rect 8386 5828 8392 5840
rect 7883 5800 8392 5828
rect 7883 5797 7895 5800
rect 7837 5791 7895 5797
rect 6638 5760 6644 5772
rect 6472 5732 6644 5760
rect 6638 5720 6644 5732
rect 6696 5760 6702 5772
rect 6748 5760 6776 5791
rect 8386 5788 8392 5800
rect 8444 5788 8450 5840
rect 11348 5828 11376 5856
rect 11256 5800 11376 5828
rect 11517 5831 11575 5837
rect 6825 5763 6883 5769
rect 6825 5760 6837 5763
rect 6696 5732 6837 5760
rect 6696 5720 6702 5732
rect 6825 5729 6837 5732
rect 6871 5729 6883 5763
rect 6825 5723 6883 5729
rect 7466 5720 7472 5772
rect 7524 5760 7530 5772
rect 7561 5763 7619 5769
rect 7561 5760 7573 5763
rect 7524 5732 7573 5760
rect 7524 5720 7530 5732
rect 7561 5729 7573 5732
rect 7607 5729 7619 5763
rect 7561 5723 7619 5729
rect 7745 5763 7803 5769
rect 7745 5729 7757 5763
rect 7791 5760 7803 5763
rect 9030 5760 9036 5772
rect 7791 5732 9036 5760
rect 7791 5729 7803 5732
rect 7745 5723 7803 5729
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 11256 5769 11284 5800
rect 11517 5797 11529 5831
rect 11563 5828 11575 5831
rect 12176 5828 12204 5856
rect 11563 5800 12204 5828
rect 11563 5797 11575 5800
rect 11517 5791 11575 5797
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5729 11299 5763
rect 11241 5723 11299 5729
rect 11333 5763 11391 5769
rect 11333 5729 11345 5763
rect 11379 5729 11391 5763
rect 11333 5723 11391 5729
rect 6730 5692 6736 5704
rect 6196 5664 6736 5692
rect 6730 5652 6736 5664
rect 6788 5652 6794 5704
rect 5997 5627 6055 5633
rect 3620 5596 5948 5624
rect 3694 5516 3700 5568
rect 3752 5516 3758 5568
rect 5258 5516 5264 5568
rect 5316 5556 5322 5568
rect 5445 5559 5503 5565
rect 5445 5556 5457 5559
rect 5316 5528 5457 5556
rect 5316 5516 5322 5528
rect 5445 5525 5457 5528
rect 5491 5525 5503 5559
rect 5920 5556 5948 5596
rect 5997 5593 6009 5627
rect 6043 5624 6055 5627
rect 6104 5624 6132 5652
rect 7484 5624 7512 5720
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 10597 5695 10655 5701
rect 10597 5692 10609 5695
rect 10376 5664 10609 5692
rect 10376 5652 10382 5664
rect 10597 5661 10609 5664
rect 10643 5661 10655 5695
rect 10597 5655 10655 5661
rect 11146 5652 11152 5704
rect 11204 5692 11210 5704
rect 11348 5692 11376 5723
rect 12066 5720 12072 5772
rect 12124 5720 12130 5772
rect 12526 5720 12532 5772
rect 12584 5760 12590 5772
rect 13081 5763 13139 5769
rect 13081 5760 13093 5763
rect 12584 5732 13093 5760
rect 12584 5720 12590 5732
rect 13081 5729 13093 5732
rect 13127 5729 13139 5763
rect 13081 5723 13139 5729
rect 11204 5664 11376 5692
rect 12805 5695 12863 5701
rect 11204 5652 11210 5664
rect 12805 5661 12817 5695
rect 12851 5692 12863 5695
rect 12986 5692 12992 5704
rect 12851 5664 12992 5692
rect 12851 5661 12863 5664
rect 12805 5655 12863 5661
rect 12986 5652 12992 5664
rect 13044 5652 13050 5704
rect 6043 5596 6132 5624
rect 6196 5596 7512 5624
rect 6043 5593 6055 5596
rect 5997 5587 6055 5593
rect 6196 5556 6224 5596
rect 5920 5528 6224 5556
rect 6549 5559 6607 5565
rect 5445 5519 5503 5525
rect 6549 5525 6561 5559
rect 6595 5556 6607 5559
rect 6730 5556 6736 5568
rect 6595 5528 6736 5556
rect 6595 5525 6607 5528
rect 6549 5519 6607 5525
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 7742 5516 7748 5568
rect 7800 5516 7806 5568
rect 11517 5559 11575 5565
rect 11517 5525 11529 5559
rect 11563 5556 11575 5559
rect 11606 5556 11612 5568
rect 11563 5528 11612 5556
rect 11563 5525 11575 5528
rect 11517 5519 11575 5525
rect 11606 5516 11612 5528
rect 11664 5516 11670 5568
rect 14369 5559 14427 5565
rect 14369 5525 14381 5559
rect 14415 5556 14427 5559
rect 14458 5556 14464 5568
rect 14415 5528 14464 5556
rect 14415 5525 14427 5528
rect 14369 5519 14427 5525
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 552 5466 15364 5488
rect 552 5414 2249 5466
rect 2301 5414 2313 5466
rect 2365 5414 2377 5466
rect 2429 5414 2441 5466
rect 2493 5414 2505 5466
rect 2557 5414 5951 5466
rect 6003 5414 6015 5466
rect 6067 5414 6079 5466
rect 6131 5414 6143 5466
rect 6195 5414 6207 5466
rect 6259 5414 9653 5466
rect 9705 5414 9717 5466
rect 9769 5414 9781 5466
rect 9833 5414 9845 5466
rect 9897 5414 9909 5466
rect 9961 5414 13355 5466
rect 13407 5414 13419 5466
rect 13471 5414 13483 5466
rect 13535 5414 13547 5466
rect 13599 5414 13611 5466
rect 13663 5414 15364 5466
rect 552 5392 15364 5414
rect 4706 5312 4712 5364
rect 4764 5312 4770 5364
rect 6270 5312 6276 5364
rect 6328 5352 6334 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 6328 5324 6377 5352
rect 6328 5312 6334 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 6730 5312 6736 5364
rect 6788 5352 6794 5364
rect 6825 5355 6883 5361
rect 6825 5352 6837 5355
rect 6788 5324 6837 5352
rect 6788 5312 6794 5324
rect 6825 5321 6837 5324
rect 6871 5321 6883 5355
rect 6825 5315 6883 5321
rect 10318 5312 10324 5364
rect 10376 5312 10382 5364
rect 12710 5312 12716 5364
rect 12768 5352 12774 5364
rect 12897 5355 12955 5361
rect 12897 5352 12909 5355
rect 12768 5324 12909 5352
rect 12768 5312 12774 5324
rect 12897 5321 12909 5324
rect 12943 5352 12955 5355
rect 14550 5352 14556 5364
rect 12943 5324 14556 5352
rect 12943 5321 12955 5324
rect 12897 5315 12955 5321
rect 14550 5312 14556 5324
rect 14608 5312 14614 5364
rect 3326 5176 3332 5228
rect 3384 5176 3390 5228
rect 11333 5219 11391 5225
rect 11333 5216 11345 5219
rect 11026 5188 11345 5216
rect 3344 5148 3372 5176
rect 5258 5157 5264 5160
rect 4985 5151 5043 5157
rect 4985 5148 4997 5151
rect 3344 5120 4997 5148
rect 4985 5117 4997 5120
rect 5031 5117 5043 5151
rect 5252 5148 5264 5157
rect 5219 5120 5264 5148
rect 4985 5111 5043 5117
rect 5252 5111 5264 5120
rect 5258 5108 5264 5111
rect 5316 5108 5322 5160
rect 7926 5108 7932 5160
rect 7984 5157 7990 5160
rect 7984 5111 7996 5157
rect 8205 5151 8263 5157
rect 8205 5117 8217 5151
rect 8251 5148 8263 5151
rect 8941 5151 8999 5157
rect 8941 5148 8953 5151
rect 8251 5120 8953 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 8941 5117 8953 5120
rect 8987 5148 8999 5151
rect 9490 5148 9496 5160
rect 8987 5120 9496 5148
rect 8987 5117 8999 5120
rect 8941 5111 8999 5117
rect 7984 5108 7990 5111
rect 9490 5108 9496 5120
rect 9548 5148 9554 5160
rect 11026 5148 11054 5188
rect 11333 5185 11345 5188
rect 11379 5216 11391 5219
rect 12986 5216 12992 5228
rect 11379 5188 12992 5216
rect 11379 5185 11391 5188
rect 11333 5179 11391 5185
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 9548 5120 11054 5148
rect 9548 5108 9554 5120
rect 11606 5108 11612 5160
rect 11664 5108 11670 5160
rect 3596 5083 3654 5089
rect 3596 5049 3608 5083
rect 3642 5080 3654 5083
rect 3694 5080 3700 5092
rect 3642 5052 3700 5080
rect 3642 5049 3654 5052
rect 3596 5043 3654 5049
rect 3694 5040 3700 5052
rect 3752 5040 3758 5092
rect 9208 5083 9266 5089
rect 9208 5049 9220 5083
rect 9254 5080 9266 5083
rect 9306 5080 9312 5092
rect 9254 5052 9312 5080
rect 9254 5049 9266 5052
rect 9208 5043 9266 5049
rect 9306 5040 9312 5052
rect 9364 5040 9370 5092
rect 552 4922 15520 4944
rect 552 4870 4100 4922
rect 4152 4870 4164 4922
rect 4216 4870 4228 4922
rect 4280 4870 4292 4922
rect 4344 4870 4356 4922
rect 4408 4870 7802 4922
rect 7854 4870 7866 4922
rect 7918 4870 7930 4922
rect 7982 4870 7994 4922
rect 8046 4870 8058 4922
rect 8110 4870 11504 4922
rect 11556 4870 11568 4922
rect 11620 4870 11632 4922
rect 11684 4870 11696 4922
rect 11748 4870 11760 4922
rect 11812 4870 15206 4922
rect 15258 4870 15270 4922
rect 15322 4870 15334 4922
rect 15386 4870 15398 4922
rect 15450 4870 15462 4922
rect 15514 4870 15520 4922
rect 552 4848 15520 4870
rect 552 4378 15364 4400
rect 552 4326 2249 4378
rect 2301 4326 2313 4378
rect 2365 4326 2377 4378
rect 2429 4326 2441 4378
rect 2493 4326 2505 4378
rect 2557 4326 5951 4378
rect 6003 4326 6015 4378
rect 6067 4326 6079 4378
rect 6131 4326 6143 4378
rect 6195 4326 6207 4378
rect 6259 4326 9653 4378
rect 9705 4326 9717 4378
rect 9769 4326 9781 4378
rect 9833 4326 9845 4378
rect 9897 4326 9909 4378
rect 9961 4326 13355 4378
rect 13407 4326 13419 4378
rect 13471 4326 13483 4378
rect 13535 4326 13547 4378
rect 13599 4326 13611 4378
rect 13663 4326 15364 4378
rect 552 4304 15364 4326
rect 11241 4267 11299 4273
rect 11241 4233 11253 4267
rect 11287 4264 11299 4267
rect 12342 4264 12348 4276
rect 11287 4236 12348 4264
rect 11287 4233 11299 4236
rect 11241 4227 11299 4233
rect 12342 4224 12348 4236
rect 12400 4264 12406 4276
rect 12802 4264 12808 4276
rect 12400 4236 12808 4264
rect 12400 4224 12406 4236
rect 12802 4224 12808 4236
rect 12860 4224 12866 4276
rect 9490 4088 9496 4140
rect 9548 4128 9554 4140
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 9548 4100 9689 4128
rect 9548 4088 9554 4100
rect 9677 4097 9689 4100
rect 9723 4097 9735 4131
rect 9677 4091 9735 4097
rect 9950 4088 9956 4140
rect 10008 4088 10014 4140
rect 552 3834 15520 3856
rect 552 3782 4100 3834
rect 4152 3782 4164 3834
rect 4216 3782 4228 3834
rect 4280 3782 4292 3834
rect 4344 3782 4356 3834
rect 4408 3782 7802 3834
rect 7854 3782 7866 3834
rect 7918 3782 7930 3834
rect 7982 3782 7994 3834
rect 8046 3782 8058 3834
rect 8110 3782 11504 3834
rect 11556 3782 11568 3834
rect 11620 3782 11632 3834
rect 11684 3782 11696 3834
rect 11748 3782 11760 3834
rect 11812 3782 15206 3834
rect 15258 3782 15270 3834
rect 15322 3782 15334 3834
rect 15386 3782 15398 3834
rect 15450 3782 15462 3834
rect 15514 3782 15520 3834
rect 552 3760 15520 3782
rect 552 3290 15364 3312
rect 552 3238 2249 3290
rect 2301 3238 2313 3290
rect 2365 3238 2377 3290
rect 2429 3238 2441 3290
rect 2493 3238 2505 3290
rect 2557 3238 5951 3290
rect 6003 3238 6015 3290
rect 6067 3238 6079 3290
rect 6131 3238 6143 3290
rect 6195 3238 6207 3290
rect 6259 3238 9653 3290
rect 9705 3238 9717 3290
rect 9769 3238 9781 3290
rect 9833 3238 9845 3290
rect 9897 3238 9909 3290
rect 9961 3238 13355 3290
rect 13407 3238 13419 3290
rect 13471 3238 13483 3290
rect 13535 3238 13547 3290
rect 13599 3238 13611 3290
rect 13663 3238 15364 3290
rect 552 3216 15364 3238
rect 552 2746 15520 2768
rect 552 2694 4100 2746
rect 4152 2694 4164 2746
rect 4216 2694 4228 2746
rect 4280 2694 4292 2746
rect 4344 2694 4356 2746
rect 4408 2694 7802 2746
rect 7854 2694 7866 2746
rect 7918 2694 7930 2746
rect 7982 2694 7994 2746
rect 8046 2694 8058 2746
rect 8110 2694 11504 2746
rect 11556 2694 11568 2746
rect 11620 2694 11632 2746
rect 11684 2694 11696 2746
rect 11748 2694 11760 2746
rect 11812 2694 15206 2746
rect 15258 2694 15270 2746
rect 15322 2694 15334 2746
rect 15386 2694 15398 2746
rect 15450 2694 15462 2746
rect 15514 2694 15520 2746
rect 552 2672 15520 2694
rect 552 2202 15364 2224
rect 552 2150 2249 2202
rect 2301 2150 2313 2202
rect 2365 2150 2377 2202
rect 2429 2150 2441 2202
rect 2493 2150 2505 2202
rect 2557 2150 5951 2202
rect 6003 2150 6015 2202
rect 6067 2150 6079 2202
rect 6131 2150 6143 2202
rect 6195 2150 6207 2202
rect 6259 2150 9653 2202
rect 9705 2150 9717 2202
rect 9769 2150 9781 2202
rect 9833 2150 9845 2202
rect 9897 2150 9909 2202
rect 9961 2150 13355 2202
rect 13407 2150 13419 2202
rect 13471 2150 13483 2202
rect 13535 2150 13547 2202
rect 13599 2150 13611 2202
rect 13663 2150 15364 2202
rect 552 2128 15364 2150
rect 552 1658 15520 1680
rect 552 1606 4100 1658
rect 4152 1606 4164 1658
rect 4216 1606 4228 1658
rect 4280 1606 4292 1658
rect 4344 1606 4356 1658
rect 4408 1606 7802 1658
rect 7854 1606 7866 1658
rect 7918 1606 7930 1658
rect 7982 1606 7994 1658
rect 8046 1606 8058 1658
rect 8110 1606 11504 1658
rect 11556 1606 11568 1658
rect 11620 1606 11632 1658
rect 11684 1606 11696 1658
rect 11748 1606 11760 1658
rect 11812 1606 15206 1658
rect 15258 1606 15270 1658
rect 15322 1606 15334 1658
rect 15386 1606 15398 1658
rect 15450 1606 15462 1658
rect 15514 1606 15520 1658
rect 552 1584 15520 1606
rect 552 1114 15364 1136
rect 552 1062 2249 1114
rect 2301 1062 2313 1114
rect 2365 1062 2377 1114
rect 2429 1062 2441 1114
rect 2493 1062 2505 1114
rect 2557 1062 5951 1114
rect 6003 1062 6015 1114
rect 6067 1062 6079 1114
rect 6131 1062 6143 1114
rect 6195 1062 6207 1114
rect 6259 1062 9653 1114
rect 9705 1062 9717 1114
rect 9769 1062 9781 1114
rect 9833 1062 9845 1114
rect 9897 1062 9909 1114
rect 9961 1062 13355 1114
rect 13407 1062 13419 1114
rect 13471 1062 13483 1114
rect 13535 1062 13547 1114
rect 13599 1062 13611 1114
rect 13663 1062 15364 1114
rect 552 1040 15364 1062
rect 552 570 15520 592
rect 552 518 4100 570
rect 4152 518 4164 570
rect 4216 518 4228 570
rect 4280 518 4292 570
rect 4344 518 4356 570
rect 4408 518 7802 570
rect 7854 518 7866 570
rect 7918 518 7930 570
rect 7982 518 7994 570
rect 8046 518 8058 570
rect 8110 518 11504 570
rect 11556 518 11568 570
rect 11620 518 11632 570
rect 11684 518 11696 570
rect 11748 518 11760 570
rect 11812 518 15206 570
rect 15258 518 15270 570
rect 15322 518 15334 570
rect 15386 518 15398 570
rect 15450 518 15462 570
rect 15514 518 15520 570
rect 552 496 15520 518
<< via1 >>
rect 4988 15308 5040 15360
rect 12164 15308 12216 15360
rect 2249 15206 2301 15258
rect 2313 15206 2365 15258
rect 2377 15206 2429 15258
rect 2441 15206 2493 15258
rect 2505 15206 2557 15258
rect 5951 15206 6003 15258
rect 6015 15206 6067 15258
rect 6079 15206 6131 15258
rect 6143 15206 6195 15258
rect 6207 15206 6259 15258
rect 9653 15206 9705 15258
rect 9717 15206 9769 15258
rect 9781 15206 9833 15258
rect 9845 15206 9897 15258
rect 9909 15206 9961 15258
rect 13355 15206 13407 15258
rect 13419 15206 13471 15258
rect 13483 15206 13535 15258
rect 13547 15206 13599 15258
rect 13611 15206 13663 15258
rect 6092 15147 6144 15156
rect 6092 15113 6101 15147
rect 6101 15113 6135 15147
rect 6135 15113 6144 15147
rect 6092 15104 6144 15113
rect 6276 15104 6328 15156
rect 6460 15104 6512 15156
rect 11428 15104 11480 15156
rect 10048 15036 10100 15088
rect 11152 15036 11204 15088
rect 2136 14900 2188 14952
rect 3424 14900 3476 14952
rect 4712 14900 4764 14952
rect 6000 14900 6052 14952
rect 6276 14900 6328 14952
rect 6368 14943 6420 14952
rect 6368 14909 6377 14943
rect 6377 14909 6411 14943
rect 6411 14909 6420 14943
rect 6368 14900 6420 14909
rect 7288 14900 7340 14952
rect 8392 14943 8444 14952
rect 8392 14909 8401 14943
rect 8401 14909 8435 14943
rect 8435 14909 8444 14943
rect 8392 14900 8444 14909
rect 4988 14832 5040 14884
rect 8576 14900 8628 14952
rect 2136 14807 2188 14816
rect 2136 14773 2145 14807
rect 2145 14773 2179 14807
rect 2179 14773 2188 14807
rect 2136 14764 2188 14773
rect 2596 14807 2648 14816
rect 2596 14773 2605 14807
rect 2605 14773 2639 14807
rect 2639 14773 2648 14807
rect 2596 14764 2648 14773
rect 5724 14764 5776 14816
rect 5816 14807 5868 14816
rect 5816 14773 5825 14807
rect 5825 14773 5859 14807
rect 5859 14773 5868 14807
rect 5816 14764 5868 14773
rect 8484 14832 8536 14884
rect 10140 14943 10192 14952
rect 10140 14909 10149 14943
rect 10149 14909 10183 14943
rect 10183 14909 10192 14943
rect 10140 14900 10192 14909
rect 12808 15036 12860 15088
rect 12440 14900 12492 14952
rect 13176 14943 13228 14952
rect 13176 14909 13185 14943
rect 13185 14909 13219 14943
rect 13219 14909 13228 14943
rect 13176 14900 13228 14909
rect 13728 14900 13780 14952
rect 15016 14943 15068 14952
rect 15016 14909 15025 14943
rect 15025 14909 15059 14943
rect 15059 14909 15068 14943
rect 15016 14900 15068 14909
rect 7564 14807 7616 14816
rect 7564 14773 7573 14807
rect 7573 14773 7607 14807
rect 7607 14773 7616 14807
rect 7564 14764 7616 14773
rect 8944 14807 8996 14816
rect 8944 14773 8953 14807
rect 8953 14773 8987 14807
rect 8987 14773 8996 14807
rect 8944 14764 8996 14773
rect 9036 14807 9088 14816
rect 9036 14773 9045 14807
rect 9045 14773 9079 14807
rect 9079 14773 9088 14807
rect 9036 14764 9088 14773
rect 9496 14764 9548 14816
rect 10416 14807 10468 14816
rect 10416 14773 10425 14807
rect 10425 14773 10459 14807
rect 10459 14773 10468 14807
rect 10416 14764 10468 14773
rect 11336 14807 11388 14816
rect 11336 14773 11345 14807
rect 11345 14773 11379 14807
rect 11379 14773 11388 14807
rect 11336 14764 11388 14773
rect 11980 14764 12032 14816
rect 12256 14764 12308 14816
rect 12716 14807 12768 14816
rect 12716 14773 12725 14807
rect 12725 14773 12759 14807
rect 12759 14773 12768 14807
rect 12716 14764 12768 14773
rect 13268 14807 13320 14816
rect 13268 14773 13277 14807
rect 13277 14773 13311 14807
rect 13311 14773 13320 14807
rect 13268 14764 13320 14773
rect 13820 14764 13872 14816
rect 14188 14764 14240 14816
rect 4100 14662 4152 14714
rect 4164 14662 4216 14714
rect 4228 14662 4280 14714
rect 4292 14662 4344 14714
rect 4356 14662 4408 14714
rect 7802 14662 7854 14714
rect 7866 14662 7918 14714
rect 7930 14662 7982 14714
rect 7994 14662 8046 14714
rect 8058 14662 8110 14714
rect 11504 14662 11556 14714
rect 11568 14662 11620 14714
rect 11632 14662 11684 14714
rect 11696 14662 11748 14714
rect 11760 14662 11812 14714
rect 15206 14662 15258 14714
rect 15270 14662 15322 14714
rect 15334 14662 15386 14714
rect 15398 14662 15450 14714
rect 15462 14662 15514 14714
rect 2136 14560 2188 14612
rect 2688 14492 2740 14544
rect 5816 14560 5868 14612
rect 7380 14560 7432 14612
rect 8392 14560 8444 14612
rect 9404 14560 9456 14612
rect 10140 14560 10192 14612
rect 11980 14560 12032 14612
rect 13176 14560 13228 14612
rect 6460 14492 6512 14544
rect 5540 14424 5592 14476
rect 6000 14424 6052 14476
rect 3332 14356 3384 14408
rect 6276 14399 6328 14408
rect 6276 14365 6285 14399
rect 6285 14365 6319 14399
rect 6319 14365 6328 14399
rect 6276 14356 6328 14365
rect 7564 14424 7616 14476
rect 8300 14424 8352 14476
rect 10232 14424 10284 14476
rect 10324 14467 10376 14476
rect 10324 14433 10333 14467
rect 10333 14433 10367 14467
rect 10367 14433 10376 14467
rect 10324 14424 10376 14433
rect 12072 14467 12124 14476
rect 12072 14433 12090 14467
rect 12090 14433 12124 14467
rect 12072 14424 12124 14433
rect 12808 14467 12860 14476
rect 12808 14433 12825 14467
rect 12825 14433 12860 14467
rect 12808 14424 12860 14433
rect 12900 14467 12952 14476
rect 12900 14433 12909 14467
rect 12909 14433 12943 14467
rect 12943 14433 12952 14467
rect 12900 14424 12952 14433
rect 12992 14467 13044 14476
rect 12992 14433 13001 14467
rect 13001 14433 13035 14467
rect 13035 14433 13044 14467
rect 12992 14424 13044 14433
rect 13084 14467 13136 14476
rect 13084 14433 13093 14467
rect 13093 14433 13127 14467
rect 13127 14433 13136 14467
rect 13084 14424 13136 14433
rect 15016 14467 15068 14476
rect 15016 14433 15025 14467
rect 15025 14433 15059 14467
rect 15059 14433 15068 14467
rect 15016 14424 15068 14433
rect 3884 14288 3936 14340
rect 3148 14220 3200 14272
rect 5816 14220 5868 14272
rect 6092 14220 6144 14272
rect 6276 14220 6328 14272
rect 6552 14263 6604 14272
rect 6552 14229 6561 14263
rect 6561 14229 6595 14263
rect 6595 14229 6604 14263
rect 6552 14220 6604 14229
rect 6920 14220 6972 14272
rect 12440 14220 12492 14272
rect 13728 14356 13780 14408
rect 14004 14220 14056 14272
rect 2249 14118 2301 14170
rect 2313 14118 2365 14170
rect 2377 14118 2429 14170
rect 2441 14118 2493 14170
rect 2505 14118 2557 14170
rect 5951 14118 6003 14170
rect 6015 14118 6067 14170
rect 6079 14118 6131 14170
rect 6143 14118 6195 14170
rect 6207 14118 6259 14170
rect 9653 14118 9705 14170
rect 9717 14118 9769 14170
rect 9781 14118 9833 14170
rect 9845 14118 9897 14170
rect 9909 14118 9961 14170
rect 13355 14118 13407 14170
rect 13419 14118 13471 14170
rect 13483 14118 13535 14170
rect 13547 14118 13599 14170
rect 13611 14118 13663 14170
rect 2596 14016 2648 14068
rect 2688 14016 2740 14068
rect 3884 14016 3936 14068
rect 6276 14016 6328 14068
rect 5632 13948 5684 14000
rect 6368 13948 6420 14000
rect 6552 13948 6604 14000
rect 8300 14016 8352 14068
rect 8576 14016 8628 14068
rect 10232 14059 10284 14068
rect 10232 14025 10241 14059
rect 10241 14025 10275 14059
rect 10275 14025 10284 14059
rect 10232 14016 10284 14025
rect 12072 14016 12124 14068
rect 13084 14016 13136 14068
rect 13728 14016 13780 14068
rect 3332 13812 3384 13864
rect 5540 13855 5592 13864
rect 5540 13821 5549 13855
rect 5549 13821 5583 13855
rect 5583 13821 5592 13855
rect 5540 13812 5592 13821
rect 5724 13855 5776 13864
rect 5724 13821 5733 13855
rect 5733 13821 5767 13855
rect 5767 13821 5776 13855
rect 5724 13812 5776 13821
rect 6920 13880 6972 13932
rect 8944 13880 8996 13932
rect 9496 13880 9548 13932
rect 12256 13948 12308 14000
rect 11336 13923 11388 13932
rect 11336 13889 11345 13923
rect 11345 13889 11379 13923
rect 11379 13889 11388 13923
rect 11336 13880 11388 13889
rect 12808 13880 12860 13932
rect 8668 13855 8720 13864
rect 8668 13821 8677 13855
rect 8677 13821 8711 13855
rect 8711 13821 8720 13855
rect 9956 13855 10008 13864
rect 8668 13812 8720 13821
rect 9956 13821 9965 13855
rect 9965 13821 9999 13855
rect 9999 13821 10008 13855
rect 9956 13812 10008 13821
rect 10416 13812 10468 13864
rect 11888 13812 11940 13864
rect 12164 13812 12216 13864
rect 15016 13880 15068 13932
rect 13268 13812 13320 13864
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 5816 13676 5868 13728
rect 7564 13676 7616 13728
rect 10508 13676 10560 13728
rect 13268 13676 13320 13728
rect 13360 13676 13412 13728
rect 4100 13574 4152 13626
rect 4164 13574 4216 13626
rect 4228 13574 4280 13626
rect 4292 13574 4344 13626
rect 4356 13574 4408 13626
rect 7802 13574 7854 13626
rect 7866 13574 7918 13626
rect 7930 13574 7982 13626
rect 7994 13574 8046 13626
rect 8058 13574 8110 13626
rect 11504 13574 11556 13626
rect 11568 13574 11620 13626
rect 11632 13574 11684 13626
rect 11696 13574 11748 13626
rect 11760 13574 11812 13626
rect 15206 13574 15258 13626
rect 15270 13574 15322 13626
rect 15334 13574 15386 13626
rect 15398 13574 15450 13626
rect 15462 13574 15514 13626
rect 6460 13379 6512 13388
rect 6460 13345 6469 13379
rect 6469 13345 6503 13379
rect 6503 13345 6512 13379
rect 6460 13336 6512 13345
rect 8668 13336 8720 13388
rect 8852 13379 8904 13388
rect 8852 13345 8861 13379
rect 8861 13345 8895 13379
rect 8895 13345 8904 13379
rect 8852 13336 8904 13345
rect 12716 13472 12768 13524
rect 13820 13472 13872 13524
rect 9956 13379 10008 13388
rect 9956 13345 9965 13379
rect 9965 13345 9999 13379
rect 9999 13345 10008 13379
rect 9956 13336 10008 13345
rect 11888 13336 11940 13388
rect 12624 13336 12676 13388
rect 13728 13404 13780 13456
rect 8484 13268 8536 13320
rect 10140 13268 10192 13320
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 9036 13200 9088 13252
rect 12348 13268 12400 13320
rect 13360 13268 13412 13320
rect 14004 13379 14056 13388
rect 14004 13345 14013 13379
rect 14013 13345 14047 13379
rect 14047 13345 14056 13379
rect 14004 13336 14056 13345
rect 14188 13379 14240 13388
rect 14188 13345 14197 13379
rect 14197 13345 14231 13379
rect 14231 13345 14240 13379
rect 14188 13336 14240 13345
rect 14464 13336 14516 13388
rect 13728 13268 13780 13320
rect 6460 13132 6512 13184
rect 7656 13132 7708 13184
rect 8576 13132 8628 13184
rect 8668 13132 8720 13184
rect 9496 13132 9548 13184
rect 10048 13132 10100 13184
rect 11888 13175 11940 13184
rect 11888 13141 11897 13175
rect 11897 13141 11931 13175
rect 11931 13141 11940 13175
rect 11888 13132 11940 13141
rect 12992 13175 13044 13184
rect 12992 13141 13001 13175
rect 13001 13141 13035 13175
rect 13035 13141 13044 13175
rect 12992 13132 13044 13141
rect 13912 13175 13964 13184
rect 13912 13141 13921 13175
rect 13921 13141 13955 13175
rect 13955 13141 13964 13175
rect 13912 13132 13964 13141
rect 14188 13132 14240 13184
rect 2249 13030 2301 13082
rect 2313 13030 2365 13082
rect 2377 13030 2429 13082
rect 2441 13030 2493 13082
rect 2505 13030 2557 13082
rect 5951 13030 6003 13082
rect 6015 13030 6067 13082
rect 6079 13030 6131 13082
rect 6143 13030 6195 13082
rect 6207 13030 6259 13082
rect 9653 13030 9705 13082
rect 9717 13030 9769 13082
rect 9781 13030 9833 13082
rect 9845 13030 9897 13082
rect 9909 13030 9961 13082
rect 13355 13030 13407 13082
rect 13419 13030 13471 13082
rect 13483 13030 13535 13082
rect 13547 13030 13599 13082
rect 13611 13030 13663 13082
rect 5632 12928 5684 12980
rect 5724 12928 5776 12980
rect 12992 12971 13044 12980
rect 12992 12937 13001 12971
rect 13001 12937 13035 12971
rect 13035 12937 13044 12971
rect 12992 12928 13044 12937
rect 13728 12928 13780 12980
rect 9312 12860 9364 12912
rect 12624 12860 12676 12912
rect 3332 12724 3384 12776
rect 3792 12656 3844 12708
rect 4712 12588 4764 12640
rect 7656 12767 7708 12776
rect 7656 12733 7674 12767
rect 7674 12733 7708 12767
rect 7656 12724 7708 12733
rect 10324 12835 10376 12844
rect 10324 12801 10333 12835
rect 10333 12801 10367 12835
rect 10367 12801 10376 12835
rect 10324 12792 10376 12801
rect 12164 12767 12216 12776
rect 5724 12631 5776 12640
rect 5724 12597 5733 12631
rect 5733 12597 5767 12631
rect 5767 12597 5776 12631
rect 5724 12588 5776 12597
rect 5908 12588 5960 12640
rect 7564 12588 7616 12640
rect 8760 12631 8812 12640
rect 8760 12597 8769 12631
rect 8769 12597 8803 12631
rect 8803 12597 8812 12631
rect 8760 12588 8812 12597
rect 12164 12733 12173 12767
rect 12173 12733 12207 12767
rect 12207 12733 12216 12767
rect 12164 12724 12216 12733
rect 12992 12724 13044 12776
rect 10048 12699 10100 12708
rect 10048 12665 10066 12699
rect 10066 12665 10100 12699
rect 10048 12656 10100 12665
rect 11888 12699 11940 12708
rect 11888 12665 11906 12699
rect 11906 12665 11940 12699
rect 11888 12656 11940 12665
rect 13084 12656 13136 12708
rect 13728 12767 13780 12776
rect 13728 12733 13737 12767
rect 13737 12733 13771 12767
rect 13771 12733 13780 12767
rect 13728 12724 13780 12733
rect 14188 12777 14240 12786
rect 14188 12743 14197 12777
rect 14197 12743 14231 12777
rect 14231 12743 14240 12777
rect 14188 12734 14240 12743
rect 13452 12656 13504 12708
rect 14280 12767 14332 12776
rect 14280 12733 14295 12767
rect 14295 12733 14329 12767
rect 14329 12733 14332 12767
rect 14280 12724 14332 12733
rect 14464 12767 14516 12776
rect 14464 12733 14473 12767
rect 14473 12733 14507 12767
rect 14507 12733 14516 12767
rect 14464 12724 14516 12733
rect 9036 12588 9088 12640
rect 10600 12588 10652 12640
rect 13544 12588 13596 12640
rect 15016 12656 15068 12708
rect 14004 12588 14056 12640
rect 14464 12588 14516 12640
rect 4100 12486 4152 12538
rect 4164 12486 4216 12538
rect 4228 12486 4280 12538
rect 4292 12486 4344 12538
rect 4356 12486 4408 12538
rect 7802 12486 7854 12538
rect 7866 12486 7918 12538
rect 7930 12486 7982 12538
rect 7994 12486 8046 12538
rect 8058 12486 8110 12538
rect 11504 12486 11556 12538
rect 11568 12486 11620 12538
rect 11632 12486 11684 12538
rect 11696 12486 11748 12538
rect 11760 12486 11812 12538
rect 15206 12486 15258 12538
rect 15270 12486 15322 12538
rect 15334 12486 15386 12538
rect 15398 12486 15450 12538
rect 15462 12486 15514 12538
rect 848 12384 900 12436
rect 7288 12384 7340 12436
rect 10140 12384 10192 12436
rect 11244 12384 11296 12436
rect 13084 12384 13136 12436
rect 14280 12384 14332 12436
rect 2596 12316 2648 12368
rect 3792 12359 3844 12368
rect 3792 12325 3801 12359
rect 3801 12325 3835 12359
rect 3835 12325 3844 12359
rect 3792 12316 3844 12325
rect 5724 12316 5776 12368
rect 3608 12248 3660 12300
rect 3884 12291 3936 12300
rect 3884 12257 3893 12291
rect 3893 12257 3927 12291
rect 3927 12257 3936 12291
rect 3884 12248 3936 12257
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 5908 12291 5960 12300
rect 5908 12257 5917 12291
rect 5917 12257 5951 12291
rect 5951 12257 5960 12291
rect 5908 12248 5960 12257
rect 4712 12180 4764 12232
rect 5632 12180 5684 12232
rect 6276 12291 6328 12300
rect 6276 12257 6285 12291
rect 6285 12257 6319 12291
rect 6319 12257 6328 12291
rect 6276 12248 6328 12257
rect 15016 12359 15068 12368
rect 15016 12325 15025 12359
rect 15025 12325 15059 12359
rect 15059 12325 15068 12359
rect 15016 12316 15068 12325
rect 3516 12155 3568 12164
rect 3516 12121 3525 12155
rect 3525 12121 3559 12155
rect 3559 12121 3568 12155
rect 3516 12112 3568 12121
rect 4344 12155 4396 12164
rect 4344 12121 4353 12155
rect 4353 12121 4387 12155
rect 4387 12121 4396 12155
rect 7472 12291 7524 12300
rect 7472 12257 7481 12291
rect 7481 12257 7515 12291
rect 7515 12257 7524 12291
rect 7472 12248 7524 12257
rect 7564 12291 7616 12300
rect 7564 12257 7573 12291
rect 7573 12257 7607 12291
rect 7607 12257 7616 12291
rect 7564 12248 7616 12257
rect 8852 12248 8904 12300
rect 9496 12291 9548 12300
rect 9496 12257 9505 12291
rect 9505 12257 9539 12291
rect 9539 12257 9548 12291
rect 9496 12248 9548 12257
rect 10232 12248 10284 12300
rect 10600 12248 10652 12300
rect 12164 12248 12216 12300
rect 13268 12248 13320 12300
rect 13912 12248 13964 12300
rect 8484 12180 8536 12232
rect 14096 12180 14148 12232
rect 14464 12180 14516 12232
rect 4344 12112 4396 12121
rect 7656 12112 7708 12164
rect 8116 12112 8168 12164
rect 9404 12112 9456 12164
rect 5540 12087 5592 12096
rect 5540 12053 5549 12087
rect 5549 12053 5583 12087
rect 5583 12053 5592 12087
rect 5540 12044 5592 12053
rect 7196 12044 7248 12096
rect 7380 12044 7432 12096
rect 8208 12044 8260 12096
rect 8760 12044 8812 12096
rect 9496 12087 9548 12096
rect 9496 12053 9505 12087
rect 9505 12053 9539 12087
rect 9539 12053 9548 12087
rect 9496 12044 9548 12053
rect 11428 12087 11480 12096
rect 11428 12053 11437 12087
rect 11437 12053 11471 12087
rect 11471 12053 11480 12087
rect 11428 12044 11480 12053
rect 2249 11942 2301 11994
rect 2313 11942 2365 11994
rect 2377 11942 2429 11994
rect 2441 11942 2493 11994
rect 2505 11942 2557 11994
rect 5951 11942 6003 11994
rect 6015 11942 6067 11994
rect 6079 11942 6131 11994
rect 6143 11942 6195 11994
rect 6207 11942 6259 11994
rect 9653 11942 9705 11994
rect 9717 11942 9769 11994
rect 9781 11942 9833 11994
rect 9845 11942 9897 11994
rect 9909 11942 9961 11994
rect 13355 11942 13407 11994
rect 13419 11942 13471 11994
rect 13483 11942 13535 11994
rect 13547 11942 13599 11994
rect 13611 11942 13663 11994
rect 2596 11840 2648 11892
rect 3516 11840 3568 11892
rect 3700 11772 3752 11824
rect 3976 11772 4028 11824
rect 5632 11883 5684 11892
rect 5632 11849 5641 11883
rect 5641 11849 5675 11883
rect 5675 11849 5684 11883
rect 5632 11840 5684 11849
rect 6276 11840 6328 11892
rect 7472 11840 7524 11892
rect 9036 11840 9088 11892
rect 4896 11772 4948 11824
rect 5724 11772 5776 11824
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 12072 11840 12124 11892
rect 10600 11772 10652 11824
rect 4068 11704 4120 11756
rect 3608 11636 3660 11688
rect 3792 11568 3844 11620
rect 3976 11679 4028 11688
rect 3976 11645 3985 11679
rect 3985 11645 4019 11679
rect 4019 11645 4028 11679
rect 3976 11636 4028 11645
rect 4344 11636 4396 11688
rect 4804 11636 4856 11688
rect 6552 11679 6604 11688
rect 6552 11645 6561 11679
rect 6561 11645 6595 11679
rect 6595 11645 6604 11679
rect 6552 11636 6604 11645
rect 7196 11636 7248 11688
rect 7380 11636 7432 11688
rect 7656 11679 7708 11688
rect 7656 11645 7666 11679
rect 7666 11645 7700 11679
rect 7700 11645 7708 11679
rect 7656 11636 7708 11645
rect 8116 11636 8168 11688
rect 8208 11636 8260 11688
rect 8668 11679 8720 11688
rect 8668 11645 8677 11679
rect 8677 11645 8711 11679
rect 8711 11645 8720 11679
rect 8668 11636 8720 11645
rect 9404 11747 9456 11756
rect 9404 11713 9413 11747
rect 9413 11713 9447 11747
rect 9447 11713 9456 11747
rect 9404 11704 9456 11713
rect 9588 11704 9640 11756
rect 4528 11500 4580 11552
rect 4620 11543 4672 11552
rect 4620 11509 4629 11543
rect 4629 11509 4663 11543
rect 4663 11509 4672 11543
rect 4620 11500 4672 11509
rect 4712 11543 4764 11552
rect 4712 11509 4721 11543
rect 4721 11509 4755 11543
rect 4755 11509 4764 11543
rect 4712 11500 4764 11509
rect 5448 11568 5500 11620
rect 6368 11543 6420 11552
rect 6368 11509 6377 11543
rect 6377 11509 6411 11543
rect 6411 11509 6420 11543
rect 6368 11500 6420 11509
rect 8300 11568 8352 11620
rect 9128 11543 9180 11552
rect 9128 11509 9137 11543
rect 9137 11509 9171 11543
rect 9171 11509 9180 11543
rect 9128 11500 9180 11509
rect 9680 11636 9732 11688
rect 9588 11568 9640 11620
rect 10692 11611 10744 11620
rect 10692 11577 10701 11611
rect 10701 11577 10735 11611
rect 10735 11577 10744 11611
rect 10692 11568 10744 11577
rect 9956 11543 10008 11552
rect 9956 11509 9965 11543
rect 9965 11509 9999 11543
rect 9999 11509 10008 11543
rect 9956 11500 10008 11509
rect 11152 11543 11204 11552
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 11152 11500 11204 11509
rect 11336 11543 11388 11552
rect 11336 11509 11345 11543
rect 11345 11509 11379 11543
rect 11379 11509 11388 11543
rect 11336 11500 11388 11509
rect 11428 11500 11480 11552
rect 11980 11500 12032 11552
rect 4100 11398 4152 11450
rect 4164 11398 4216 11450
rect 4228 11398 4280 11450
rect 4292 11398 4344 11450
rect 4356 11398 4408 11450
rect 7802 11398 7854 11450
rect 7866 11398 7918 11450
rect 7930 11398 7982 11450
rect 7994 11398 8046 11450
rect 8058 11398 8110 11450
rect 11504 11398 11556 11450
rect 11568 11398 11620 11450
rect 11632 11398 11684 11450
rect 11696 11398 11748 11450
rect 11760 11398 11812 11450
rect 15206 11398 15258 11450
rect 15270 11398 15322 11450
rect 15334 11398 15386 11450
rect 15398 11398 15450 11450
rect 15462 11398 15514 11450
rect 2136 11296 2188 11348
rect 2136 11203 2188 11212
rect 3884 11296 3936 11348
rect 2136 11169 2154 11203
rect 2154 11169 2188 11203
rect 2136 11160 2188 11169
rect 3332 11160 3384 11212
rect 3516 11203 3568 11212
rect 3516 11169 3525 11203
rect 3525 11169 3559 11203
rect 3559 11169 3568 11203
rect 3516 11160 3568 11169
rect 2688 10956 2740 11008
rect 3240 10999 3292 11008
rect 3240 10965 3249 10999
rect 3249 10965 3283 10999
rect 3283 10965 3292 10999
rect 3240 10956 3292 10965
rect 3792 11203 3844 11212
rect 3792 11169 3801 11203
rect 3801 11169 3835 11203
rect 3835 11169 3844 11203
rect 3792 11160 3844 11169
rect 3976 11228 4028 11280
rect 5264 11296 5316 11348
rect 8668 11296 8720 11348
rect 4068 11203 4120 11212
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 3976 10956 4028 11008
rect 4528 11135 4580 11144
rect 4528 11101 4537 11135
rect 4537 11101 4571 11135
rect 4571 11101 4580 11135
rect 4528 11092 4580 11101
rect 4620 11135 4672 11144
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 4252 11024 4304 11076
rect 4436 11067 4488 11076
rect 4436 11033 4445 11067
rect 4445 11033 4479 11067
rect 4479 11033 4488 11067
rect 4436 11024 4488 11033
rect 4896 11237 4948 11246
rect 4896 11203 4905 11237
rect 4905 11203 4939 11237
rect 4939 11203 4948 11237
rect 4896 11194 4948 11203
rect 6368 11228 6420 11280
rect 4988 11092 5040 11144
rect 5540 11160 5592 11212
rect 8300 11160 8352 11212
rect 8944 11203 8996 11212
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 9680 11228 9732 11280
rect 9404 11160 9456 11212
rect 12716 11296 12768 11348
rect 10692 11228 10744 11280
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 11152 11203 11204 11212
rect 11152 11169 11161 11203
rect 11161 11169 11195 11203
rect 11195 11169 11204 11203
rect 11152 11160 11204 11169
rect 5724 11092 5776 11144
rect 9036 11135 9088 11144
rect 9036 11101 9045 11135
rect 9045 11101 9079 11135
rect 9079 11101 9088 11135
rect 9036 11092 9088 11101
rect 10876 11092 10928 11144
rect 11980 11203 12032 11212
rect 11980 11169 11989 11203
rect 11989 11169 12023 11203
rect 12023 11169 12032 11203
rect 11980 11160 12032 11169
rect 11888 11135 11940 11144
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 12440 11092 12492 11144
rect 12624 11203 12676 11212
rect 12624 11169 12633 11203
rect 12633 11169 12667 11203
rect 12667 11169 12676 11203
rect 12624 11160 12676 11169
rect 12900 11203 12952 11212
rect 12900 11169 12909 11203
rect 12909 11169 12943 11203
rect 12943 11169 12952 11203
rect 12900 11160 12952 11169
rect 12992 11203 13044 11212
rect 12992 11169 13001 11203
rect 13001 11169 13035 11203
rect 13035 11169 13044 11203
rect 12992 11160 13044 11169
rect 13268 11160 13320 11212
rect 14280 11160 14332 11212
rect 13636 11135 13688 11144
rect 13636 11101 13645 11135
rect 13645 11101 13679 11135
rect 13679 11101 13688 11135
rect 13636 11092 13688 11101
rect 5356 10999 5408 11008
rect 5356 10965 5365 10999
rect 5365 10965 5399 10999
rect 5399 10965 5408 10999
rect 5356 10956 5408 10965
rect 5816 10956 5868 11008
rect 6920 10956 6972 11008
rect 9312 10956 9364 11008
rect 10600 10999 10652 11008
rect 10600 10965 10609 10999
rect 10609 10965 10643 10999
rect 10643 10965 10652 10999
rect 10600 10956 10652 10965
rect 11060 10956 11112 11008
rect 14004 10956 14056 11008
rect 14924 10999 14976 11008
rect 14924 10965 14933 10999
rect 14933 10965 14967 10999
rect 14967 10965 14976 10999
rect 14924 10956 14976 10965
rect 2249 10854 2301 10906
rect 2313 10854 2365 10906
rect 2377 10854 2429 10906
rect 2441 10854 2493 10906
rect 2505 10854 2557 10906
rect 5951 10854 6003 10906
rect 6015 10854 6067 10906
rect 6079 10854 6131 10906
rect 6143 10854 6195 10906
rect 6207 10854 6259 10906
rect 9653 10854 9705 10906
rect 9717 10854 9769 10906
rect 9781 10854 9833 10906
rect 9845 10854 9897 10906
rect 9909 10854 9961 10906
rect 13355 10854 13407 10906
rect 13419 10854 13471 10906
rect 13483 10854 13535 10906
rect 13547 10854 13599 10906
rect 13611 10854 13663 10906
rect 2136 10752 2188 10804
rect 3240 10752 3292 10804
rect 3332 10752 3384 10804
rect 3792 10684 3844 10736
rect 4252 10684 4304 10736
rect 4436 10752 4488 10804
rect 5724 10752 5776 10804
rect 6552 10752 6604 10804
rect 5264 10684 5316 10736
rect 5448 10684 5500 10736
rect 5816 10684 5868 10736
rect 3700 10616 3752 10668
rect 4620 10616 4672 10668
rect 2688 10591 2740 10600
rect 2688 10557 2697 10591
rect 2697 10557 2731 10591
rect 2731 10557 2740 10591
rect 2688 10548 2740 10557
rect 2780 10548 2832 10600
rect 4988 10591 5040 10600
rect 4988 10557 4997 10591
rect 4997 10557 5031 10591
rect 5031 10557 5040 10591
rect 4988 10548 5040 10557
rect 3148 10480 3200 10532
rect 5356 10591 5408 10600
rect 5356 10557 5365 10591
rect 5365 10557 5399 10591
rect 5399 10557 5408 10591
rect 5356 10548 5408 10557
rect 5448 10480 5500 10532
rect 5816 10548 5868 10600
rect 6368 10616 6420 10668
rect 8300 10752 8352 10804
rect 10324 10752 10376 10804
rect 12900 10795 12952 10804
rect 12900 10761 12909 10795
rect 12909 10761 12943 10795
rect 12943 10761 12952 10795
rect 12900 10752 12952 10761
rect 13728 10752 13780 10804
rect 14280 10795 14332 10804
rect 14280 10761 14289 10795
rect 14289 10761 14323 10795
rect 14323 10761 14332 10795
rect 14280 10752 14332 10761
rect 10048 10684 10100 10736
rect 8852 10616 8904 10668
rect 14096 10684 14148 10736
rect 6644 10591 6696 10600
rect 6644 10557 6653 10591
rect 6653 10557 6687 10591
rect 6687 10557 6696 10591
rect 6644 10548 6696 10557
rect 6920 10591 6972 10600
rect 6920 10557 6955 10591
rect 6955 10557 6972 10591
rect 6920 10548 6972 10557
rect 7472 10548 7524 10600
rect 6828 10523 6880 10532
rect 6828 10489 6837 10523
rect 6837 10489 6871 10523
rect 6871 10489 6880 10523
rect 6828 10480 6880 10489
rect 8392 10591 8444 10600
rect 8392 10557 8401 10591
rect 8401 10557 8435 10591
rect 8435 10557 8444 10591
rect 8392 10548 8444 10557
rect 11060 10616 11112 10668
rect 14556 10752 14608 10804
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 10876 10548 10928 10557
rect 11428 10548 11480 10600
rect 11336 10523 11388 10532
rect 11336 10489 11345 10523
rect 11345 10489 11379 10523
rect 11379 10489 11388 10523
rect 11336 10480 11388 10489
rect 13728 10548 13780 10600
rect 13912 10591 13964 10600
rect 13912 10557 13921 10591
rect 13921 10557 13955 10591
rect 13955 10557 13964 10591
rect 13912 10548 13964 10557
rect 14004 10591 14056 10600
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 14004 10548 14056 10557
rect 14188 10591 14240 10600
rect 14188 10557 14197 10591
rect 14197 10557 14231 10591
rect 14231 10557 14240 10591
rect 14188 10548 14240 10557
rect 14924 10480 14976 10532
rect 5356 10412 5408 10464
rect 8208 10412 8260 10464
rect 13728 10412 13780 10464
rect 14280 10412 14332 10464
rect 4100 10310 4152 10362
rect 4164 10310 4216 10362
rect 4228 10310 4280 10362
rect 4292 10310 4344 10362
rect 4356 10310 4408 10362
rect 7802 10310 7854 10362
rect 7866 10310 7918 10362
rect 7930 10310 7982 10362
rect 7994 10310 8046 10362
rect 8058 10310 8110 10362
rect 11504 10310 11556 10362
rect 11568 10310 11620 10362
rect 11632 10310 11684 10362
rect 11696 10310 11748 10362
rect 11760 10310 11812 10362
rect 15206 10310 15258 10362
rect 15270 10310 15322 10362
rect 15334 10310 15386 10362
rect 15398 10310 15450 10362
rect 15462 10310 15514 10362
rect 3976 10208 4028 10260
rect 5264 10208 5316 10260
rect 5356 10251 5408 10260
rect 5356 10217 5365 10251
rect 5365 10217 5399 10251
rect 5399 10217 5408 10251
rect 5356 10208 5408 10217
rect 6644 10208 6696 10260
rect 9128 10208 9180 10260
rect 9312 10208 9364 10260
rect 4712 10183 4764 10192
rect 4712 10149 4721 10183
rect 4721 10149 4755 10183
rect 4755 10149 4764 10183
rect 4712 10140 4764 10149
rect 5080 10072 5132 10124
rect 5448 10115 5500 10124
rect 5448 10081 5457 10115
rect 5457 10081 5491 10115
rect 5491 10081 5500 10115
rect 5448 10072 5500 10081
rect 4620 10004 4672 10056
rect 10692 10072 10744 10124
rect 11980 10072 12032 10124
rect 12440 10072 12492 10124
rect 12624 10072 12676 10124
rect 6828 9936 6880 9988
rect 11520 10047 11572 10056
rect 11520 10013 11529 10047
rect 11529 10013 11563 10047
rect 11563 10013 11572 10047
rect 11520 10004 11572 10013
rect 5080 9868 5132 9920
rect 5264 9868 5316 9920
rect 5632 9868 5684 9920
rect 9128 9911 9180 9920
rect 9128 9877 9137 9911
rect 9137 9877 9171 9911
rect 9171 9877 9180 9911
rect 9128 9868 9180 9877
rect 9312 9868 9364 9920
rect 11980 9868 12032 9920
rect 2249 9766 2301 9818
rect 2313 9766 2365 9818
rect 2377 9766 2429 9818
rect 2441 9766 2493 9818
rect 2505 9766 2557 9818
rect 5951 9766 6003 9818
rect 6015 9766 6067 9818
rect 6079 9766 6131 9818
rect 6143 9766 6195 9818
rect 6207 9766 6259 9818
rect 9653 9766 9705 9818
rect 9717 9766 9769 9818
rect 9781 9766 9833 9818
rect 9845 9766 9897 9818
rect 9909 9766 9961 9818
rect 13355 9766 13407 9818
rect 13419 9766 13471 9818
rect 13483 9766 13535 9818
rect 13547 9766 13599 9818
rect 13611 9766 13663 9818
rect 4436 9664 4488 9716
rect 3516 9639 3568 9648
rect 3516 9605 3525 9639
rect 3525 9605 3559 9639
rect 3559 9605 3568 9639
rect 3516 9596 3568 9605
rect 1492 9460 1544 9512
rect 3332 9392 3384 9444
rect 3240 9367 3292 9376
rect 3240 9333 3249 9367
rect 3249 9333 3283 9367
rect 3283 9333 3292 9367
rect 3240 9324 3292 9333
rect 4620 9596 4672 9648
rect 7932 9664 7984 9716
rect 8208 9664 8260 9716
rect 9036 9707 9088 9716
rect 9036 9673 9045 9707
rect 9045 9673 9079 9707
rect 9079 9673 9088 9707
rect 9036 9664 9088 9673
rect 3700 9571 3752 9580
rect 3700 9537 3709 9571
rect 3709 9537 3743 9571
rect 3743 9537 3752 9571
rect 3700 9528 3752 9537
rect 4896 9528 4948 9580
rect 3976 9392 4028 9444
rect 4528 9460 4580 9512
rect 5080 9528 5132 9580
rect 5264 9503 5316 9512
rect 5264 9469 5273 9503
rect 5273 9469 5307 9503
rect 5307 9469 5316 9503
rect 5264 9460 5316 9469
rect 4804 9392 4856 9444
rect 3792 9324 3844 9376
rect 4620 9367 4672 9376
rect 4620 9333 4629 9367
rect 4629 9333 4663 9367
rect 4663 9333 4672 9367
rect 4620 9324 4672 9333
rect 5632 9460 5684 9512
rect 6460 9503 6512 9512
rect 6460 9469 6469 9503
rect 6469 9469 6503 9503
rect 6503 9469 6512 9503
rect 6460 9460 6512 9469
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 7472 9460 7524 9512
rect 7564 9460 7616 9512
rect 7932 9503 7984 9512
rect 7932 9469 7941 9503
rect 7941 9469 7975 9503
rect 7975 9469 7984 9503
rect 7932 9460 7984 9469
rect 8760 9639 8812 9648
rect 8760 9605 8769 9639
rect 8769 9605 8803 9639
rect 8803 9605 8812 9639
rect 8760 9596 8812 9605
rect 9128 9528 9180 9580
rect 5540 9324 5592 9376
rect 6276 9367 6328 9376
rect 6276 9333 6285 9367
rect 6285 9333 6319 9367
rect 6319 9333 6328 9367
rect 6276 9324 6328 9333
rect 6552 9324 6604 9376
rect 7196 9392 7248 9444
rect 7656 9435 7708 9444
rect 7656 9401 7665 9435
rect 7665 9401 7699 9435
rect 7699 9401 7708 9435
rect 7656 9392 7708 9401
rect 9496 9460 9548 9512
rect 12440 9639 12492 9648
rect 12440 9605 12449 9639
rect 12449 9605 12483 9639
rect 12483 9605 12492 9639
rect 12440 9596 12492 9605
rect 14096 9571 14148 9580
rect 14096 9537 14105 9571
rect 14105 9537 14139 9571
rect 14139 9537 14148 9571
rect 14096 9528 14148 9537
rect 12992 9460 13044 9512
rect 7564 9324 7616 9376
rect 10784 9392 10836 9444
rect 9220 9367 9272 9376
rect 9220 9333 9229 9367
rect 9229 9333 9263 9367
rect 9263 9333 9272 9367
rect 9220 9324 9272 9333
rect 10600 9324 10652 9376
rect 10876 9367 10928 9376
rect 10876 9333 10885 9367
rect 10885 9333 10919 9367
rect 10919 9333 10928 9367
rect 10876 9324 10928 9333
rect 11428 9392 11480 9444
rect 12256 9392 12308 9444
rect 14280 9392 14332 9444
rect 14556 9503 14608 9512
rect 14556 9469 14565 9503
rect 14565 9469 14599 9503
rect 14599 9469 14608 9503
rect 14556 9460 14608 9469
rect 15016 9392 15068 9444
rect 11520 9324 11572 9376
rect 13084 9324 13136 9376
rect 4100 9222 4152 9274
rect 4164 9222 4216 9274
rect 4228 9222 4280 9274
rect 4292 9222 4344 9274
rect 4356 9222 4408 9274
rect 7802 9222 7854 9274
rect 7866 9222 7918 9274
rect 7930 9222 7982 9274
rect 7994 9222 8046 9274
rect 8058 9222 8110 9274
rect 11504 9222 11556 9274
rect 11568 9222 11620 9274
rect 11632 9222 11684 9274
rect 11696 9222 11748 9274
rect 11760 9222 11812 9274
rect 15206 9222 15258 9274
rect 15270 9222 15322 9274
rect 15334 9222 15386 9274
rect 15398 9222 15450 9274
rect 15462 9222 15514 9274
rect 3240 9120 3292 9172
rect 3332 9163 3384 9172
rect 3332 9129 3341 9163
rect 3341 9129 3375 9163
rect 3375 9129 3384 9163
rect 3332 9120 3384 9129
rect 3516 9120 3568 9172
rect 4620 9120 4672 9172
rect 4896 9163 4948 9172
rect 4896 9129 4905 9163
rect 4905 9129 4939 9163
rect 4939 9129 4948 9163
rect 4896 9120 4948 9129
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 7196 9120 7248 9129
rect 8392 9120 8444 9172
rect 9220 9120 9272 9172
rect 9312 9120 9364 9172
rect 10048 9120 10100 9172
rect 10692 9120 10744 9172
rect 11428 9120 11480 9172
rect 3608 8984 3660 9036
rect 3976 8984 4028 9036
rect 4436 8984 4488 9036
rect 2872 8916 2924 8968
rect 3792 8916 3844 8968
rect 5540 9052 5592 9104
rect 6276 9052 6328 9104
rect 7288 9095 7340 9104
rect 7288 9061 7297 9095
rect 7297 9061 7331 9095
rect 7331 9061 7340 9095
rect 7288 9052 7340 9061
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 9956 9027 10008 9036
rect 9956 8993 9965 9027
rect 9965 8993 9999 9027
rect 9999 8993 10008 9027
rect 9956 8984 10008 8993
rect 10232 9052 10284 9104
rect 12900 9120 12952 9172
rect 13084 9120 13136 9172
rect 10600 8984 10652 9036
rect 10784 8984 10836 9036
rect 10876 8984 10928 9036
rect 11980 8984 12032 9036
rect 3700 8848 3752 8900
rect 5724 8848 5776 8900
rect 1952 8823 2004 8832
rect 1952 8789 1961 8823
rect 1961 8789 1995 8823
rect 1995 8789 2004 8823
rect 1952 8780 2004 8789
rect 5080 8780 5132 8832
rect 7564 8780 7616 8832
rect 9128 8780 9180 8832
rect 12440 8984 12492 9036
rect 9956 8848 10008 8900
rect 10140 8780 10192 8832
rect 10692 8848 10744 8900
rect 11244 8848 11296 8900
rect 12624 8984 12676 9036
rect 14556 9120 14608 9172
rect 12900 8959 12952 8968
rect 12900 8925 12909 8959
rect 12909 8925 12943 8959
rect 12943 8925 12952 8959
rect 12900 8916 12952 8925
rect 12992 8916 13044 8968
rect 14096 8780 14148 8832
rect 15016 8780 15068 8832
rect 2249 8678 2301 8730
rect 2313 8678 2365 8730
rect 2377 8678 2429 8730
rect 2441 8678 2493 8730
rect 2505 8678 2557 8730
rect 5951 8678 6003 8730
rect 6015 8678 6067 8730
rect 6079 8678 6131 8730
rect 6143 8678 6195 8730
rect 6207 8678 6259 8730
rect 9653 8678 9705 8730
rect 9717 8678 9769 8730
rect 9781 8678 9833 8730
rect 9845 8678 9897 8730
rect 9909 8678 9961 8730
rect 13355 8678 13407 8730
rect 13419 8678 13471 8730
rect 13483 8678 13535 8730
rect 13547 8678 13599 8730
rect 13611 8678 13663 8730
rect 2872 8619 2924 8628
rect 2872 8585 2881 8619
rect 2881 8585 2915 8619
rect 2915 8585 2924 8619
rect 2872 8576 2924 8585
rect 1492 8415 1544 8424
rect 1492 8381 1501 8415
rect 1501 8381 1535 8415
rect 1535 8381 1544 8415
rect 1492 8372 1544 8381
rect 2688 8372 2740 8424
rect 4068 8508 4120 8560
rect 5264 8576 5316 8628
rect 6460 8576 6512 8628
rect 11244 8619 11296 8628
rect 11244 8585 11253 8619
rect 11253 8585 11287 8619
rect 11287 8585 11296 8619
rect 11244 8576 11296 8585
rect 12900 8576 12952 8628
rect 5632 8508 5684 8560
rect 12348 8508 12400 8560
rect 4436 8440 4488 8492
rect 6368 8440 6420 8492
rect 9220 8440 9272 8492
rect 4528 8415 4580 8424
rect 4528 8381 4537 8415
rect 4537 8381 4571 8415
rect 4571 8381 4580 8415
rect 4528 8372 4580 8381
rect 4804 8372 4856 8424
rect 5172 8372 5224 8424
rect 6552 8372 6604 8424
rect 7380 8372 7432 8424
rect 3148 8304 3200 8356
rect 3700 8304 3752 8356
rect 3792 8304 3844 8356
rect 3424 8279 3476 8288
rect 3424 8245 3433 8279
rect 3433 8245 3467 8279
rect 3467 8245 3476 8279
rect 3424 8236 3476 8245
rect 4712 8236 4764 8288
rect 4896 8279 4948 8288
rect 4896 8245 4905 8279
rect 4905 8245 4939 8279
rect 4939 8245 4948 8279
rect 4896 8236 4948 8245
rect 8760 8415 8812 8424
rect 8760 8381 8769 8415
rect 8769 8381 8803 8415
rect 8803 8381 8812 8415
rect 8760 8372 8812 8381
rect 8852 8415 8904 8424
rect 8852 8381 8861 8415
rect 8861 8381 8895 8415
rect 8895 8381 8904 8415
rect 8852 8372 8904 8381
rect 8944 8372 8996 8424
rect 9128 8415 9180 8424
rect 9128 8381 9137 8415
rect 9137 8381 9171 8415
rect 9171 8381 9180 8415
rect 9128 8372 9180 8381
rect 10140 8415 10192 8424
rect 10140 8381 10174 8415
rect 10174 8381 10192 8415
rect 9496 8304 9548 8356
rect 10140 8372 10192 8381
rect 12624 8372 12676 8424
rect 13176 8415 13228 8424
rect 13176 8381 13185 8415
rect 13185 8381 13219 8415
rect 13219 8381 13228 8415
rect 13176 8372 13228 8381
rect 14280 8372 14332 8424
rect 5632 8279 5684 8288
rect 5632 8245 5641 8279
rect 5641 8245 5675 8279
rect 5675 8245 5684 8279
rect 5632 8236 5684 8245
rect 8208 8236 8260 8288
rect 8484 8236 8536 8288
rect 9036 8236 9088 8288
rect 11980 8236 12032 8288
rect 13912 8236 13964 8288
rect 4100 8134 4152 8186
rect 4164 8134 4216 8186
rect 4228 8134 4280 8186
rect 4292 8134 4344 8186
rect 4356 8134 4408 8186
rect 7802 8134 7854 8186
rect 7866 8134 7918 8186
rect 7930 8134 7982 8186
rect 7994 8134 8046 8186
rect 8058 8134 8110 8186
rect 11504 8134 11556 8186
rect 11568 8134 11620 8186
rect 11632 8134 11684 8186
rect 11696 8134 11748 8186
rect 11760 8134 11812 8186
rect 15206 8134 15258 8186
rect 15270 8134 15322 8186
rect 15334 8134 15386 8186
rect 15398 8134 15450 8186
rect 15462 8134 15514 8186
rect 1952 8032 2004 8084
rect 3424 8032 3476 8084
rect 9496 8032 9548 8084
rect 10232 8032 10284 8084
rect 10416 8032 10468 8084
rect 2780 7964 2832 8016
rect 4988 7964 5040 8016
rect 5632 7964 5684 8016
rect 4712 7939 4764 7948
rect 4712 7905 4721 7939
rect 4721 7905 4755 7939
rect 4755 7905 4764 7939
rect 4712 7896 4764 7905
rect 7380 7939 7432 7948
rect 7380 7905 7389 7939
rect 7389 7905 7423 7939
rect 7423 7905 7432 7939
rect 7380 7896 7432 7905
rect 7656 7939 7708 7948
rect 7656 7905 7690 7939
rect 7690 7905 7708 7939
rect 7656 7896 7708 7905
rect 8576 7896 8628 7948
rect 9036 7939 9088 7948
rect 9036 7905 9045 7939
rect 9045 7905 9079 7939
rect 9079 7905 9088 7939
rect 12072 7964 12124 8016
rect 12624 7964 12676 8016
rect 9036 7896 9088 7905
rect 10600 7896 10652 7948
rect 11336 7896 11388 7948
rect 11980 7939 12032 7948
rect 11980 7905 11989 7939
rect 11989 7905 12023 7939
rect 12023 7905 12032 7939
rect 11980 7896 12032 7905
rect 4068 7828 4120 7880
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 4896 7828 4948 7880
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 12532 7896 12584 7948
rect 13176 8007 13228 8016
rect 13176 7973 13185 8007
rect 13185 7973 13219 8007
rect 13219 7973 13228 8007
rect 13176 7964 13228 7973
rect 13084 7939 13136 7948
rect 13084 7905 13091 7939
rect 13091 7905 13136 7939
rect 13084 7896 13136 7905
rect 12716 7871 12768 7880
rect 2688 7760 2740 7812
rect 3332 7760 3384 7812
rect 5816 7760 5868 7812
rect 12716 7837 12725 7871
rect 12725 7837 12759 7871
rect 12759 7837 12768 7871
rect 12716 7828 12768 7837
rect 12808 7760 12860 7812
rect 4528 7692 4580 7744
rect 9312 7692 9364 7744
rect 10232 7692 10284 7744
rect 12348 7735 12400 7744
rect 12348 7701 12357 7735
rect 12357 7701 12391 7735
rect 12391 7701 12400 7735
rect 12348 7692 12400 7701
rect 12624 7735 12676 7744
rect 12624 7701 12633 7735
rect 12633 7701 12667 7735
rect 12667 7701 12676 7735
rect 12624 7692 12676 7701
rect 14004 7692 14056 7744
rect 2249 7590 2301 7642
rect 2313 7590 2365 7642
rect 2377 7590 2429 7642
rect 2441 7590 2493 7642
rect 2505 7590 2557 7642
rect 5951 7590 6003 7642
rect 6015 7590 6067 7642
rect 6079 7590 6131 7642
rect 6143 7590 6195 7642
rect 6207 7590 6259 7642
rect 9653 7590 9705 7642
rect 9717 7590 9769 7642
rect 9781 7590 9833 7642
rect 9845 7590 9897 7642
rect 9909 7590 9961 7642
rect 13355 7590 13407 7642
rect 13419 7590 13471 7642
rect 13483 7590 13535 7642
rect 13547 7590 13599 7642
rect 13611 7590 13663 7642
rect 4436 7488 4488 7540
rect 4804 7531 4856 7540
rect 4804 7497 4813 7531
rect 4813 7497 4847 7531
rect 4847 7497 4856 7531
rect 4804 7488 4856 7497
rect 7656 7488 7708 7540
rect 2872 7420 2924 7472
rect 6368 7463 6420 7472
rect 6368 7429 6377 7463
rect 6377 7429 6411 7463
rect 6411 7429 6420 7463
rect 6368 7420 6420 7429
rect 4068 7352 4120 7404
rect 10968 7488 11020 7540
rect 12256 7488 12308 7540
rect 13084 7488 13136 7540
rect 4620 7327 4672 7336
rect 2872 7148 2924 7200
rect 3884 7148 3936 7200
rect 4620 7293 4629 7327
rect 4629 7293 4663 7327
rect 4663 7293 4672 7327
rect 4620 7284 4672 7293
rect 4712 7284 4764 7336
rect 5816 7284 5868 7336
rect 5356 7216 5408 7268
rect 7472 7216 7524 7268
rect 7748 7284 7800 7336
rect 8208 7284 8260 7336
rect 9404 7327 9456 7336
rect 9404 7293 9413 7327
rect 9413 7293 9447 7327
rect 9447 7293 9456 7327
rect 9404 7284 9456 7293
rect 10140 7463 10192 7472
rect 10140 7429 10149 7463
rect 10149 7429 10183 7463
rect 10183 7429 10192 7463
rect 10140 7420 10192 7429
rect 10232 7420 10284 7472
rect 4528 7148 4580 7200
rect 4896 7148 4948 7200
rect 7564 7148 7616 7200
rect 9496 7191 9548 7200
rect 9496 7157 9505 7191
rect 9505 7157 9539 7191
rect 9539 7157 9548 7191
rect 9496 7148 9548 7157
rect 10508 7284 10560 7336
rect 11428 7327 11480 7336
rect 11428 7293 11437 7327
rect 11437 7293 11471 7327
rect 11471 7293 11480 7327
rect 11428 7284 11480 7293
rect 10600 7216 10652 7268
rect 11060 7259 11112 7268
rect 11060 7225 11069 7259
rect 11069 7225 11103 7259
rect 11103 7225 11112 7259
rect 11060 7216 11112 7225
rect 11244 7148 11296 7200
rect 12256 7148 12308 7200
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 13912 7327 13964 7336
rect 13912 7293 13921 7327
rect 13921 7293 13955 7327
rect 13955 7293 13964 7327
rect 13912 7284 13964 7293
rect 14004 7327 14056 7336
rect 14004 7293 14013 7327
rect 14013 7293 14047 7327
rect 14047 7293 14056 7327
rect 14004 7284 14056 7293
rect 14188 7327 14240 7336
rect 14188 7293 14197 7327
rect 14197 7293 14231 7327
rect 14231 7293 14240 7327
rect 14188 7284 14240 7293
rect 15016 7284 15068 7336
rect 12532 7216 12584 7268
rect 12716 7148 12768 7200
rect 13636 7148 13688 7200
rect 4100 7046 4152 7098
rect 4164 7046 4216 7098
rect 4228 7046 4280 7098
rect 4292 7046 4344 7098
rect 4356 7046 4408 7098
rect 7802 7046 7854 7098
rect 7866 7046 7918 7098
rect 7930 7046 7982 7098
rect 7994 7046 8046 7098
rect 8058 7046 8110 7098
rect 11504 7046 11556 7098
rect 11568 7046 11620 7098
rect 11632 7046 11684 7098
rect 11696 7046 11748 7098
rect 11760 7046 11812 7098
rect 15206 7046 15258 7098
rect 15270 7046 15322 7098
rect 15334 7046 15386 7098
rect 15398 7046 15450 7098
rect 15462 7046 15514 7098
rect 3608 6944 3660 6996
rect 2872 6876 2924 6928
rect 2780 6808 2832 6860
rect 3792 6808 3844 6860
rect 3884 6851 3936 6860
rect 4712 6876 4764 6928
rect 3884 6817 3900 6851
rect 3900 6817 3934 6851
rect 3934 6817 3936 6851
rect 3884 6808 3936 6817
rect 5356 6987 5408 6996
rect 5356 6953 5365 6987
rect 5365 6953 5399 6987
rect 5399 6953 5408 6987
rect 5356 6944 5408 6953
rect 7564 6944 7616 6996
rect 7656 6944 7708 6996
rect 9496 6944 9548 6996
rect 11060 6944 11112 6996
rect 12440 6944 12492 6996
rect 12532 6987 12584 6996
rect 12532 6953 12541 6987
rect 12541 6953 12575 6987
rect 12575 6953 12584 6987
rect 12532 6944 12584 6953
rect 2780 6647 2832 6656
rect 2780 6613 2789 6647
rect 2789 6613 2823 6647
rect 2823 6613 2832 6647
rect 2780 6604 2832 6613
rect 4160 6604 4212 6656
rect 4528 6740 4580 6792
rect 5816 6808 5868 6860
rect 6368 6851 6420 6860
rect 6368 6817 6377 6851
rect 6377 6817 6411 6851
rect 6411 6817 6420 6851
rect 6368 6808 6420 6817
rect 6644 6851 6696 6860
rect 6644 6817 6653 6851
rect 6653 6817 6687 6851
rect 6687 6817 6696 6851
rect 6644 6808 6696 6817
rect 11428 6876 11480 6928
rect 8484 6808 8536 6860
rect 14464 6876 14516 6928
rect 12992 6808 13044 6860
rect 13636 6851 13688 6860
rect 13636 6817 13645 6851
rect 13645 6817 13679 6851
rect 13679 6817 13688 6851
rect 13636 6808 13688 6817
rect 15016 6851 15068 6860
rect 15016 6817 15025 6851
rect 15025 6817 15059 6851
rect 15059 6817 15068 6851
rect 15016 6808 15068 6817
rect 6736 6715 6788 6724
rect 6736 6681 6745 6715
rect 6745 6681 6779 6715
rect 6779 6681 6788 6715
rect 6736 6672 6788 6681
rect 4436 6604 4488 6656
rect 5724 6604 5776 6656
rect 6276 6604 6328 6656
rect 8852 6672 8904 6724
rect 12624 6672 12676 6724
rect 12716 6647 12768 6656
rect 12716 6613 12725 6647
rect 12725 6613 12759 6647
rect 12759 6613 12768 6647
rect 12716 6604 12768 6613
rect 12808 6604 12860 6656
rect 2249 6502 2301 6554
rect 2313 6502 2365 6554
rect 2377 6502 2429 6554
rect 2441 6502 2493 6554
rect 2505 6502 2557 6554
rect 5951 6502 6003 6554
rect 6015 6502 6067 6554
rect 6079 6502 6131 6554
rect 6143 6502 6195 6554
rect 6207 6502 6259 6554
rect 9653 6502 9705 6554
rect 9717 6502 9769 6554
rect 9781 6502 9833 6554
rect 9845 6502 9897 6554
rect 9909 6502 9961 6554
rect 13355 6502 13407 6554
rect 13419 6502 13471 6554
rect 13483 6502 13535 6554
rect 13547 6502 13599 6554
rect 13611 6502 13663 6554
rect 2780 6400 2832 6452
rect 4160 6400 4212 6452
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 4528 6400 4580 6452
rect 6736 6400 6788 6452
rect 10048 6400 10100 6452
rect 10968 6443 11020 6452
rect 10968 6409 10977 6443
rect 10977 6409 11011 6443
rect 11011 6409 11020 6443
rect 10968 6400 11020 6409
rect 14280 6443 14332 6452
rect 14280 6409 14289 6443
rect 14289 6409 14323 6443
rect 14323 6409 14332 6443
rect 14280 6400 14332 6409
rect 5540 6332 5592 6384
rect 6368 6332 6420 6384
rect 6644 6332 6696 6384
rect 9772 6332 9824 6384
rect 3608 6196 3660 6248
rect 4436 6239 4488 6248
rect 4436 6205 4445 6239
rect 4445 6205 4479 6239
rect 4479 6205 4488 6239
rect 4436 6196 4488 6205
rect 4528 6239 4580 6248
rect 4528 6205 4537 6239
rect 4537 6205 4571 6239
rect 4571 6205 4580 6239
rect 4528 6196 4580 6205
rect 4712 6239 4764 6248
rect 4712 6205 4721 6239
rect 4721 6205 4755 6239
rect 4755 6205 4764 6239
rect 4712 6196 4764 6205
rect 7840 6307 7892 6316
rect 7840 6273 7849 6307
rect 7849 6273 7883 6307
rect 7883 6273 7892 6307
rect 10232 6332 10284 6384
rect 12072 6332 12124 6384
rect 12440 6332 12492 6384
rect 15016 6332 15068 6384
rect 7840 6264 7892 6273
rect 6000 6239 6052 6248
rect 6000 6205 6009 6239
rect 6009 6205 6043 6239
rect 6043 6205 6052 6239
rect 6000 6196 6052 6205
rect 6092 6239 6144 6248
rect 6092 6205 6101 6239
rect 6101 6205 6135 6239
rect 6135 6205 6144 6239
rect 6092 6196 6144 6205
rect 6276 6196 6328 6248
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 6736 6171 6788 6180
rect 6736 6137 6745 6171
rect 6745 6137 6779 6171
rect 6779 6137 6788 6171
rect 8484 6196 8536 6248
rect 9036 6196 9088 6248
rect 6736 6128 6788 6137
rect 2872 6060 2924 6112
rect 3884 6103 3936 6112
rect 3884 6069 3893 6103
rect 3893 6069 3927 6103
rect 3927 6069 3936 6103
rect 3884 6060 3936 6069
rect 5724 6103 5776 6112
rect 5724 6069 5733 6103
rect 5733 6069 5767 6103
rect 5767 6069 5776 6103
rect 5724 6060 5776 6069
rect 6644 6103 6696 6112
rect 6644 6069 6653 6103
rect 6653 6069 6687 6103
rect 6687 6069 6696 6103
rect 6644 6060 6696 6069
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 7840 6060 7892 6112
rect 9036 6103 9088 6112
rect 9036 6069 9045 6103
rect 9045 6069 9079 6103
rect 9079 6069 9088 6103
rect 9036 6060 9088 6069
rect 9128 6060 9180 6112
rect 9680 6196 9732 6248
rect 9772 6239 9824 6248
rect 9772 6205 9781 6239
rect 9781 6205 9815 6239
rect 9815 6205 9824 6239
rect 9772 6196 9824 6205
rect 10048 6239 10100 6248
rect 10048 6205 10057 6239
rect 10057 6205 10091 6239
rect 10091 6205 10100 6239
rect 10048 6196 10100 6205
rect 10232 6128 10284 6180
rect 11244 6239 11296 6248
rect 11244 6205 11253 6239
rect 11253 6205 11287 6239
rect 11287 6205 11296 6239
rect 11244 6196 11296 6205
rect 11428 6239 11480 6248
rect 11428 6205 11437 6239
rect 11437 6205 11471 6239
rect 11471 6205 11480 6239
rect 11428 6196 11480 6205
rect 12348 6196 12400 6248
rect 14464 6196 14516 6248
rect 10324 6060 10376 6112
rect 11152 6103 11204 6112
rect 11152 6069 11161 6103
rect 11161 6069 11195 6103
rect 11195 6069 11204 6103
rect 11152 6060 11204 6069
rect 11336 6103 11388 6112
rect 11336 6069 11345 6103
rect 11345 6069 11379 6103
rect 11379 6069 11388 6103
rect 11336 6060 11388 6069
rect 12532 6103 12584 6112
rect 12532 6069 12541 6103
rect 12541 6069 12575 6103
rect 12575 6069 12584 6103
rect 12532 6060 12584 6069
rect 12808 6060 12860 6112
rect 14556 6103 14608 6112
rect 14556 6069 14565 6103
rect 14565 6069 14599 6103
rect 14599 6069 14608 6103
rect 14556 6060 14608 6069
rect 4100 5958 4152 6010
rect 4164 5958 4216 6010
rect 4228 5958 4280 6010
rect 4292 5958 4344 6010
rect 4356 5958 4408 6010
rect 7802 5958 7854 6010
rect 7866 5958 7918 6010
rect 7930 5958 7982 6010
rect 7994 5958 8046 6010
rect 8058 5958 8110 6010
rect 11504 5958 11556 6010
rect 11568 5958 11620 6010
rect 11632 5958 11684 6010
rect 11696 5958 11748 6010
rect 11760 5958 11812 6010
rect 15206 5958 15258 6010
rect 15270 5958 15322 6010
rect 15334 5958 15386 6010
rect 15398 5958 15450 6010
rect 15462 5958 15514 6010
rect 3884 5856 3936 5908
rect 3976 5856 4028 5908
rect 3700 5831 3752 5840
rect 3700 5797 3709 5831
rect 3709 5797 3743 5831
rect 3743 5797 3752 5831
rect 3700 5788 3752 5797
rect 3608 5720 3660 5772
rect 6000 5856 6052 5908
rect 6552 5899 6604 5908
rect 6552 5865 6574 5899
rect 6574 5865 6604 5899
rect 6552 5856 6604 5865
rect 6828 5856 6880 5908
rect 7380 5856 7432 5908
rect 9220 5856 9272 5908
rect 9772 5856 9824 5908
rect 11336 5856 11388 5908
rect 12164 5899 12216 5908
rect 12164 5865 12173 5899
rect 12173 5865 12207 5899
rect 12207 5865 12216 5899
rect 12164 5856 12216 5865
rect 4712 5720 4764 5772
rect 5724 5720 5776 5772
rect 6000 5763 6052 5772
rect 6000 5729 6009 5763
rect 6009 5729 6043 5763
rect 6043 5729 6052 5763
rect 6000 5720 6052 5729
rect 6092 5652 6144 5704
rect 6368 5720 6420 5772
rect 6644 5720 6696 5772
rect 8392 5788 8444 5840
rect 7472 5720 7524 5772
rect 9036 5720 9088 5772
rect 6736 5652 6788 5704
rect 3700 5559 3752 5568
rect 3700 5525 3709 5559
rect 3709 5525 3743 5559
rect 3743 5525 3752 5559
rect 3700 5516 3752 5525
rect 5264 5516 5316 5568
rect 10324 5652 10376 5704
rect 11152 5652 11204 5704
rect 12072 5763 12124 5772
rect 12072 5729 12081 5763
rect 12081 5729 12115 5763
rect 12115 5729 12124 5763
rect 12072 5720 12124 5729
rect 12532 5720 12584 5772
rect 12992 5652 13044 5704
rect 6736 5516 6788 5568
rect 7748 5559 7800 5568
rect 7748 5525 7757 5559
rect 7757 5525 7791 5559
rect 7791 5525 7800 5559
rect 7748 5516 7800 5525
rect 11612 5516 11664 5568
rect 14464 5516 14516 5568
rect 2249 5414 2301 5466
rect 2313 5414 2365 5466
rect 2377 5414 2429 5466
rect 2441 5414 2493 5466
rect 2505 5414 2557 5466
rect 5951 5414 6003 5466
rect 6015 5414 6067 5466
rect 6079 5414 6131 5466
rect 6143 5414 6195 5466
rect 6207 5414 6259 5466
rect 9653 5414 9705 5466
rect 9717 5414 9769 5466
rect 9781 5414 9833 5466
rect 9845 5414 9897 5466
rect 9909 5414 9961 5466
rect 13355 5414 13407 5466
rect 13419 5414 13471 5466
rect 13483 5414 13535 5466
rect 13547 5414 13599 5466
rect 13611 5414 13663 5466
rect 4712 5355 4764 5364
rect 4712 5321 4721 5355
rect 4721 5321 4755 5355
rect 4755 5321 4764 5355
rect 4712 5312 4764 5321
rect 6276 5312 6328 5364
rect 6736 5312 6788 5364
rect 10324 5355 10376 5364
rect 10324 5321 10333 5355
rect 10333 5321 10367 5355
rect 10367 5321 10376 5355
rect 10324 5312 10376 5321
rect 12716 5312 12768 5364
rect 14556 5312 14608 5364
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 5264 5151 5316 5160
rect 5264 5117 5298 5151
rect 5298 5117 5316 5151
rect 5264 5108 5316 5117
rect 7932 5151 7984 5160
rect 7932 5117 7950 5151
rect 7950 5117 7984 5151
rect 7932 5108 7984 5117
rect 9496 5108 9548 5160
rect 12992 5176 13044 5228
rect 11612 5151 11664 5160
rect 11612 5117 11621 5151
rect 11621 5117 11655 5151
rect 11655 5117 11664 5151
rect 11612 5108 11664 5117
rect 3700 5040 3752 5092
rect 9312 5040 9364 5092
rect 4100 4870 4152 4922
rect 4164 4870 4216 4922
rect 4228 4870 4280 4922
rect 4292 4870 4344 4922
rect 4356 4870 4408 4922
rect 7802 4870 7854 4922
rect 7866 4870 7918 4922
rect 7930 4870 7982 4922
rect 7994 4870 8046 4922
rect 8058 4870 8110 4922
rect 11504 4870 11556 4922
rect 11568 4870 11620 4922
rect 11632 4870 11684 4922
rect 11696 4870 11748 4922
rect 11760 4870 11812 4922
rect 15206 4870 15258 4922
rect 15270 4870 15322 4922
rect 15334 4870 15386 4922
rect 15398 4870 15450 4922
rect 15462 4870 15514 4922
rect 2249 4326 2301 4378
rect 2313 4326 2365 4378
rect 2377 4326 2429 4378
rect 2441 4326 2493 4378
rect 2505 4326 2557 4378
rect 5951 4326 6003 4378
rect 6015 4326 6067 4378
rect 6079 4326 6131 4378
rect 6143 4326 6195 4378
rect 6207 4326 6259 4378
rect 9653 4326 9705 4378
rect 9717 4326 9769 4378
rect 9781 4326 9833 4378
rect 9845 4326 9897 4378
rect 9909 4326 9961 4378
rect 13355 4326 13407 4378
rect 13419 4326 13471 4378
rect 13483 4326 13535 4378
rect 13547 4326 13599 4378
rect 13611 4326 13663 4378
rect 12348 4224 12400 4276
rect 12808 4224 12860 4276
rect 9496 4088 9548 4140
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 4100 3782 4152 3834
rect 4164 3782 4216 3834
rect 4228 3782 4280 3834
rect 4292 3782 4344 3834
rect 4356 3782 4408 3834
rect 7802 3782 7854 3834
rect 7866 3782 7918 3834
rect 7930 3782 7982 3834
rect 7994 3782 8046 3834
rect 8058 3782 8110 3834
rect 11504 3782 11556 3834
rect 11568 3782 11620 3834
rect 11632 3782 11684 3834
rect 11696 3782 11748 3834
rect 11760 3782 11812 3834
rect 15206 3782 15258 3834
rect 15270 3782 15322 3834
rect 15334 3782 15386 3834
rect 15398 3782 15450 3834
rect 15462 3782 15514 3834
rect 2249 3238 2301 3290
rect 2313 3238 2365 3290
rect 2377 3238 2429 3290
rect 2441 3238 2493 3290
rect 2505 3238 2557 3290
rect 5951 3238 6003 3290
rect 6015 3238 6067 3290
rect 6079 3238 6131 3290
rect 6143 3238 6195 3290
rect 6207 3238 6259 3290
rect 9653 3238 9705 3290
rect 9717 3238 9769 3290
rect 9781 3238 9833 3290
rect 9845 3238 9897 3290
rect 9909 3238 9961 3290
rect 13355 3238 13407 3290
rect 13419 3238 13471 3290
rect 13483 3238 13535 3290
rect 13547 3238 13599 3290
rect 13611 3238 13663 3290
rect 4100 2694 4152 2746
rect 4164 2694 4216 2746
rect 4228 2694 4280 2746
rect 4292 2694 4344 2746
rect 4356 2694 4408 2746
rect 7802 2694 7854 2746
rect 7866 2694 7918 2746
rect 7930 2694 7982 2746
rect 7994 2694 8046 2746
rect 8058 2694 8110 2746
rect 11504 2694 11556 2746
rect 11568 2694 11620 2746
rect 11632 2694 11684 2746
rect 11696 2694 11748 2746
rect 11760 2694 11812 2746
rect 15206 2694 15258 2746
rect 15270 2694 15322 2746
rect 15334 2694 15386 2746
rect 15398 2694 15450 2746
rect 15462 2694 15514 2746
rect 2249 2150 2301 2202
rect 2313 2150 2365 2202
rect 2377 2150 2429 2202
rect 2441 2150 2493 2202
rect 2505 2150 2557 2202
rect 5951 2150 6003 2202
rect 6015 2150 6067 2202
rect 6079 2150 6131 2202
rect 6143 2150 6195 2202
rect 6207 2150 6259 2202
rect 9653 2150 9705 2202
rect 9717 2150 9769 2202
rect 9781 2150 9833 2202
rect 9845 2150 9897 2202
rect 9909 2150 9961 2202
rect 13355 2150 13407 2202
rect 13419 2150 13471 2202
rect 13483 2150 13535 2202
rect 13547 2150 13599 2202
rect 13611 2150 13663 2202
rect 4100 1606 4152 1658
rect 4164 1606 4216 1658
rect 4228 1606 4280 1658
rect 4292 1606 4344 1658
rect 4356 1606 4408 1658
rect 7802 1606 7854 1658
rect 7866 1606 7918 1658
rect 7930 1606 7982 1658
rect 7994 1606 8046 1658
rect 8058 1606 8110 1658
rect 11504 1606 11556 1658
rect 11568 1606 11620 1658
rect 11632 1606 11684 1658
rect 11696 1606 11748 1658
rect 11760 1606 11812 1658
rect 15206 1606 15258 1658
rect 15270 1606 15322 1658
rect 15334 1606 15386 1658
rect 15398 1606 15450 1658
rect 15462 1606 15514 1658
rect 2249 1062 2301 1114
rect 2313 1062 2365 1114
rect 2377 1062 2429 1114
rect 2441 1062 2493 1114
rect 2505 1062 2557 1114
rect 5951 1062 6003 1114
rect 6015 1062 6067 1114
rect 6079 1062 6131 1114
rect 6143 1062 6195 1114
rect 6207 1062 6259 1114
rect 9653 1062 9705 1114
rect 9717 1062 9769 1114
rect 9781 1062 9833 1114
rect 9845 1062 9897 1114
rect 9909 1062 9961 1114
rect 13355 1062 13407 1114
rect 13419 1062 13471 1114
rect 13483 1062 13535 1114
rect 13547 1062 13599 1114
rect 13611 1062 13663 1114
rect 4100 518 4152 570
rect 4164 518 4216 570
rect 4228 518 4280 570
rect 4292 518 4344 570
rect 4356 518 4408 570
rect 7802 518 7854 570
rect 7866 518 7918 570
rect 7930 518 7982 570
rect 7994 518 8046 570
rect 8058 518 8110 570
rect 11504 518 11556 570
rect 11568 518 11620 570
rect 11632 518 11684 570
rect 11696 518 11748 570
rect 11760 518 11812 570
rect 15206 518 15258 570
rect 15270 518 15322 570
rect 15334 518 15386 570
rect 15398 518 15450 570
rect 15462 518 15514 570
<< metal2 >>
rect 846 15600 902 16000
rect 2134 15600 2190 16000
rect 3422 15600 3478 16000
rect 4710 15600 4766 16000
rect 5998 15600 6054 16000
rect 7286 15600 7342 16000
rect 8574 15600 8630 16000
rect 9862 15600 9918 16000
rect 11150 15600 11206 16000
rect 12438 15600 12494 16000
rect 13726 15600 13782 16000
rect 15014 15600 15070 16000
rect 860 12442 888 15600
rect 2148 14958 2176 15600
rect 2249 15260 2557 15269
rect 2249 15258 2255 15260
rect 2311 15258 2335 15260
rect 2391 15258 2415 15260
rect 2471 15258 2495 15260
rect 2551 15258 2557 15260
rect 2311 15206 2313 15258
rect 2493 15206 2495 15258
rect 2249 15204 2255 15206
rect 2311 15204 2335 15206
rect 2391 15204 2415 15206
rect 2471 15204 2495 15206
rect 2551 15204 2557 15206
rect 2249 15195 2557 15204
rect 3436 14958 3464 15600
rect 4724 14958 4752 15600
rect 6012 15450 6040 15600
rect 6012 15422 6316 15450
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 2136 14952 2188 14958
rect 2136 14894 2188 14900
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 5000 14890 5028 15302
rect 5951 15260 6259 15269
rect 5951 15258 5957 15260
rect 6013 15258 6037 15260
rect 6093 15258 6117 15260
rect 6173 15258 6197 15260
rect 6253 15258 6259 15260
rect 6013 15206 6015 15258
rect 6195 15206 6197 15258
rect 5951 15204 5957 15206
rect 6013 15204 6037 15206
rect 6093 15204 6117 15206
rect 6173 15204 6197 15206
rect 6253 15204 6259 15206
rect 5951 15195 6259 15204
rect 6288 15162 6316 15422
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6000 14952 6052 14958
rect 6000 14894 6052 14900
rect 4988 14884 5040 14890
rect 4988 14826 5040 14832
rect 2136 14816 2188 14822
rect 2136 14758 2188 14764
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2148 14618 2176 14758
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 2249 14172 2557 14181
rect 2249 14170 2255 14172
rect 2311 14170 2335 14172
rect 2391 14170 2415 14172
rect 2471 14170 2495 14172
rect 2551 14170 2557 14172
rect 2311 14118 2313 14170
rect 2493 14118 2495 14170
rect 2249 14116 2255 14118
rect 2311 14116 2335 14118
rect 2391 14116 2415 14118
rect 2471 14116 2495 14118
rect 2551 14116 2557 14118
rect 2249 14107 2557 14116
rect 2608 14074 2636 14758
rect 4100 14716 4408 14725
rect 4100 14714 4106 14716
rect 4162 14714 4186 14716
rect 4242 14714 4266 14716
rect 4322 14714 4346 14716
rect 4402 14714 4408 14716
rect 4162 14662 4164 14714
rect 4344 14662 4346 14714
rect 4100 14660 4106 14662
rect 4162 14660 4186 14662
rect 4242 14660 4266 14662
rect 4322 14660 4346 14662
rect 4402 14660 4408 14662
rect 4100 14651 4408 14660
rect 2688 14544 2740 14550
rect 2688 14486 2740 14492
rect 2700 14074 2728 14486
rect 3332 14408 3384 14414
rect 3332 14350 3384 14356
rect 3148 14272 3200 14278
rect 3148 14214 3200 14220
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2249 13084 2557 13093
rect 2249 13082 2255 13084
rect 2311 13082 2335 13084
rect 2391 13082 2415 13084
rect 2471 13082 2495 13084
rect 2551 13082 2557 13084
rect 2311 13030 2313 13082
rect 2493 13030 2495 13082
rect 2249 13028 2255 13030
rect 2311 13028 2335 13030
rect 2391 13028 2415 13030
rect 2471 13028 2495 13030
rect 2551 13028 2557 13030
rect 2249 13019 2557 13028
rect 848 12436 900 12442
rect 848 12378 900 12384
rect 2596 12368 2648 12374
rect 2596 12310 2648 12316
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2148 11354 2176 12174
rect 2249 11996 2557 12005
rect 2249 11994 2255 11996
rect 2311 11994 2335 11996
rect 2391 11994 2415 11996
rect 2471 11994 2495 11996
rect 2551 11994 2557 11996
rect 2311 11942 2313 11994
rect 2493 11942 2495 11994
rect 2249 11940 2255 11942
rect 2311 11940 2335 11942
rect 2391 11940 2415 11942
rect 2471 11940 2495 11942
rect 2551 11940 2557 11942
rect 2249 11931 2557 11940
rect 2608 11898 2636 12310
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2148 10810 2176 11154
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2249 10908 2557 10917
rect 2249 10906 2255 10908
rect 2311 10906 2335 10908
rect 2391 10906 2415 10908
rect 2471 10906 2495 10908
rect 2551 10906 2557 10908
rect 2311 10854 2313 10906
rect 2493 10854 2495 10906
rect 2249 10852 2255 10854
rect 2311 10852 2335 10854
rect 2391 10852 2415 10854
rect 2471 10852 2495 10854
rect 2551 10852 2557 10854
rect 2249 10843 2557 10852
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2700 10606 2728 10950
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2249 9820 2557 9829
rect 2249 9818 2255 9820
rect 2311 9818 2335 9820
rect 2391 9818 2415 9820
rect 2471 9818 2495 9820
rect 2551 9818 2557 9820
rect 2311 9766 2313 9818
rect 2493 9766 2495 9818
rect 2249 9764 2255 9766
rect 2311 9764 2335 9766
rect 2391 9764 2415 9766
rect 2471 9764 2495 9766
rect 2551 9764 2557 9766
rect 2249 9755 2557 9764
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1504 8430 1532 9454
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 1504 6914 1532 8366
rect 1964 8090 1992 8774
rect 2249 8732 2557 8741
rect 2249 8730 2255 8732
rect 2311 8730 2335 8732
rect 2391 8730 2415 8732
rect 2471 8730 2495 8732
rect 2551 8730 2557 8732
rect 2311 8678 2313 8730
rect 2493 8678 2495 8730
rect 2249 8676 2255 8678
rect 2311 8676 2335 8678
rect 2391 8676 2415 8678
rect 2471 8676 2495 8678
rect 2551 8676 2557 8678
rect 2249 8667 2557 8676
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 2700 7818 2728 8366
rect 2792 8022 2820 10542
rect 3160 10538 3188 14214
rect 3344 13870 3372 14350
rect 3884 14340 3936 14346
rect 3884 14282 3936 14288
rect 3896 14074 3924 14282
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3344 12782 3372 13806
rect 4100 13628 4408 13637
rect 4100 13626 4106 13628
rect 4162 13626 4186 13628
rect 4242 13626 4266 13628
rect 4322 13626 4346 13628
rect 4402 13626 4408 13628
rect 4162 13574 4164 13626
rect 4344 13574 4346 13626
rect 4100 13572 4106 13574
rect 4162 13572 4186 13574
rect 4242 13572 4266 13574
rect 4322 13572 4346 13574
rect 4402 13572 4408 13574
rect 4100 13563 4408 13572
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3344 11218 3372 12718
rect 3792 12708 3844 12714
rect 3792 12650 3844 12656
rect 3804 12374 3832 12650
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4100 12540 4408 12549
rect 4100 12538 4106 12540
rect 4162 12538 4186 12540
rect 4242 12538 4266 12540
rect 4322 12538 4346 12540
rect 4402 12538 4408 12540
rect 4162 12486 4164 12538
rect 4344 12486 4346 12538
rect 4100 12484 4106 12486
rect 4162 12484 4186 12486
rect 4242 12484 4266 12486
rect 4322 12484 4346 12486
rect 4402 12484 4408 12486
rect 4100 12475 4408 12484
rect 3792 12368 3844 12374
rect 3792 12310 3844 12316
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3528 11898 3556 12106
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3620 11694 3648 12242
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3514 11248 3570 11257
rect 3332 11212 3384 11218
rect 3514 11183 3516 11192
rect 3332 11154 3384 11160
rect 3568 11183 3570 11192
rect 3516 11154 3568 11160
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 3252 10810 3280 10950
rect 3344 10810 3372 11154
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3148 10532 3200 10538
rect 3148 10474 3200 10480
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 8634 2912 8910
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2249 7644 2557 7653
rect 2249 7642 2255 7644
rect 2311 7642 2335 7644
rect 2391 7642 2415 7644
rect 2471 7642 2495 7644
rect 2551 7642 2557 7644
rect 2311 7590 2313 7642
rect 2493 7590 2495 7642
rect 2249 7588 2255 7590
rect 2311 7588 2335 7590
rect 2391 7588 2415 7590
rect 2471 7588 2495 7590
rect 2551 7588 2557 7590
rect 2249 7579 2557 7588
rect 1412 6886 1532 6914
rect 1412 6322 1440 6886
rect 2792 6866 2820 7958
rect 2884 7478 2912 8570
rect 3160 8362 3188 10474
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3332 9444 3384 9450
rect 3332 9386 3384 9392
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 9178 3280 9318
rect 3344 9178 3372 9386
rect 3528 9178 3556 9590
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3620 9042 3648 11630
rect 3712 10674 3740 11766
rect 3792 11620 3844 11626
rect 3792 11562 3844 11568
rect 3804 11218 3832 11562
rect 3896 11354 3924 12242
rect 4724 12238 4752 12582
rect 5000 12434 5028 14826
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5552 13870 5580 14418
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5644 12986 5672 13942
rect 5736 13870 5764 14758
rect 5828 14618 5856 14758
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 6012 14482 6040 14894
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 6104 14278 6132 15098
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6288 14414 6316 14894
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 6092 14272 6144 14278
rect 6092 14214 6144 14220
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5736 12986 5764 13806
rect 5828 13734 5856 14214
rect 5951 14172 6259 14181
rect 5951 14170 5957 14172
rect 6013 14170 6037 14172
rect 6093 14170 6117 14172
rect 6173 14170 6197 14172
rect 6253 14170 6259 14172
rect 6013 14118 6015 14170
rect 6195 14118 6197 14170
rect 5951 14116 5957 14118
rect 6013 14116 6037 14118
rect 6093 14116 6117 14118
rect 6173 14116 6197 14118
rect 6253 14116 6259 14118
rect 5951 14107 6259 14116
rect 6288 14074 6316 14214
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6380 14006 6408 14894
rect 6472 14550 6500 15098
rect 7300 14958 7328 15600
rect 8588 14958 8616 15600
rect 9876 15450 9904 15600
rect 9876 15422 10088 15450
rect 9653 15260 9961 15269
rect 9653 15258 9659 15260
rect 9715 15258 9739 15260
rect 9795 15258 9819 15260
rect 9875 15258 9899 15260
rect 9955 15258 9961 15260
rect 9715 15206 9717 15258
rect 9897 15206 9899 15258
rect 9653 15204 9659 15206
rect 9715 15204 9739 15206
rect 9795 15204 9819 15206
rect 9875 15204 9899 15206
rect 9955 15204 9961 15206
rect 9653 15195 9961 15204
rect 10060 15094 10088 15422
rect 11164 15094 11192 15600
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 8392 14952 8444 14958
rect 8392 14894 8444 14900
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 6460 14544 6512 14550
rect 6460 14486 6512 14492
rect 6368 14000 6420 14006
rect 6368 13942 6420 13948
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5000 12406 5212 12434
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4344 12164 4396 12170
rect 4344 12106 4396 12112
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 3988 11694 4016 11766
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 4080 11540 4108 11698
rect 4356 11694 4384 12106
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4724 11558 4752 12174
rect 4896 11824 4948 11830
rect 4896 11766 4948 11772
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 3988 11512 4108 11540
rect 4528 11552 4580 11558
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3988 11286 4016 11512
rect 4528 11494 4580 11500
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4100 11452 4408 11461
rect 4100 11450 4106 11452
rect 4162 11450 4186 11452
rect 4242 11450 4266 11452
rect 4322 11450 4346 11452
rect 4402 11450 4408 11452
rect 4162 11398 4164 11450
rect 4344 11398 4346 11450
rect 4100 11396 4106 11398
rect 4162 11396 4186 11398
rect 4242 11396 4266 11398
rect 4322 11396 4346 11398
rect 4402 11396 4408 11398
rect 4100 11387 4408 11396
rect 3976 11280 4028 11286
rect 4540 11268 4568 11494
rect 3976 11222 4028 11228
rect 4066 11248 4122 11257
rect 3792 11212 3844 11218
rect 4066 11183 4068 11192
rect 3792 11154 3844 11160
rect 4120 11183 4122 11192
rect 4356 11240 4568 11268
rect 4632 11257 4660 11494
rect 4618 11248 4674 11257
rect 4068 11154 4120 11160
rect 3804 10742 3832 11154
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3712 9586 3740 10610
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 8090 3464 8230
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3332 7812 3384 7818
rect 3332 7754 3384 7760
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2884 6934 2912 7142
rect 2872 6928 2924 6934
rect 2872 6870 2924 6876
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2249 6556 2557 6565
rect 2249 6554 2255 6556
rect 2311 6554 2335 6556
rect 2391 6554 2415 6556
rect 2471 6554 2495 6556
rect 2551 6554 2557 6556
rect 2311 6502 2313 6554
rect 2493 6502 2495 6554
rect 2249 6500 2255 6502
rect 2311 6500 2335 6502
rect 2391 6500 2415 6502
rect 2471 6500 2495 6502
rect 2551 6500 2557 6502
rect 2249 6491 2557 6500
rect 2792 6458 2820 6598
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 2884 6118 2912 6870
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2249 5468 2557 5477
rect 2249 5466 2255 5468
rect 2311 5466 2335 5468
rect 2391 5466 2415 5468
rect 2471 5466 2495 5468
rect 2551 5466 2557 5468
rect 2311 5414 2313 5466
rect 2493 5414 2495 5466
rect 2249 5412 2255 5414
rect 2311 5412 2335 5414
rect 2391 5412 2415 5414
rect 2471 5412 2495 5414
rect 2551 5412 2557 5414
rect 2249 5403 2557 5412
rect 3344 5234 3372 7754
rect 3620 7002 3648 8978
rect 3712 8906 3740 9522
rect 3804 9382 3832 10678
rect 3988 10266 4016 10950
rect 4264 10742 4292 11018
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 4356 10554 4384 11240
rect 4618 11183 4674 11192
rect 4528 11144 4580 11150
rect 4526 11112 4528 11121
rect 4620 11144 4672 11150
rect 4580 11112 4582 11121
rect 4436 11076 4488 11082
rect 4620 11086 4672 11092
rect 4526 11047 4582 11056
rect 4436 11018 4488 11024
rect 4448 10810 4476 11018
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4632 10674 4660 11086
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4356 10526 4568 10554
rect 4100 10364 4408 10373
rect 4100 10362 4106 10364
rect 4162 10362 4186 10364
rect 4242 10362 4266 10364
rect 4322 10362 4346 10364
rect 4402 10362 4408 10364
rect 4162 10310 4164 10362
rect 4344 10310 4346 10362
rect 4100 10308 4106 10310
rect 4162 10308 4186 10310
rect 4242 10308 4266 10310
rect 4322 10308 4346 10310
rect 4402 10308 4408 10310
rect 4100 10299 4408 10308
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3804 8974 3832 9318
rect 3988 9042 4016 9386
rect 4100 9276 4408 9285
rect 4100 9274 4106 9276
rect 4162 9274 4186 9276
rect 4242 9274 4266 9276
rect 4322 9274 4346 9276
rect 4402 9274 4408 9276
rect 4162 9222 4164 9274
rect 4344 9222 4346 9274
rect 4100 9220 4106 9222
rect 4162 9220 4186 9222
rect 4242 9220 4266 9222
rect 4322 9220 4346 9222
rect 4402 9220 4408 9222
rect 4100 9211 4408 9220
rect 4448 9042 4476 9658
rect 4540 9518 4568 10526
rect 4724 10198 4752 11494
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4632 9654 4660 9998
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4816 9450 4844 11630
rect 4908 11252 4936 11766
rect 4896 11246 4948 11252
rect 4896 11188 4948 11194
rect 4988 11144 5040 11150
rect 4986 11112 4988 11121
rect 5040 11112 5042 11121
rect 4986 11047 5042 11056
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 4804 9444 4856 9450
rect 4804 9386 4856 9392
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4632 9178 4660 9318
rect 4908 9178 4936 9522
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 3988 8548 4016 8978
rect 4068 8560 4120 8566
rect 3988 8520 4068 8548
rect 4068 8502 4120 8508
rect 4448 8498 4476 8978
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3620 6254 3648 6938
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3620 5778 3648 6190
rect 3712 5846 3740 8298
rect 3804 6866 3832 8298
rect 4100 8188 4408 8197
rect 4100 8186 4106 8188
rect 4162 8186 4186 8188
rect 4242 8186 4266 8188
rect 4322 8186 4346 8188
rect 4402 8186 4408 8188
rect 4162 8134 4164 8186
rect 4344 8134 4346 8186
rect 4100 8132 4106 8134
rect 4162 8132 4186 8134
rect 4242 8132 4266 8134
rect 4322 8132 4346 8134
rect 4402 8132 4408 8134
rect 4100 8123 4408 8132
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4080 7410 4108 7822
rect 4448 7546 4476 8434
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4540 7750 4568 8366
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4724 7954 4752 8230
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4632 7342 4660 7822
rect 4724 7342 4752 7890
rect 4816 7546 4844 8366
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4908 7886 4936 8230
rect 5000 8022 5028 10542
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5092 9926 5120 10066
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5092 8838 5120 9522
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5184 8430 5212 12406
rect 5736 12374 5764 12582
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 5632 12232 5684 12238
rect 5828 12186 5856 13670
rect 6472 13394 6500 14486
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6564 14006 6592 14214
rect 6552 14000 6604 14006
rect 6552 13942 6604 13948
rect 6932 13938 6960 14214
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 5951 13084 6259 13093
rect 5951 13082 5957 13084
rect 6013 13082 6037 13084
rect 6093 13082 6117 13084
rect 6173 13082 6197 13084
rect 6253 13082 6259 13084
rect 6013 13030 6015 13082
rect 6195 13030 6197 13082
rect 5951 13028 5957 13030
rect 6013 13028 6037 13030
rect 6093 13028 6117 13030
rect 6173 13028 6197 13030
rect 6253 13028 6259 13030
rect 5951 13019 6259 13028
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5920 12306 5948 12582
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 5632 12174 5684 12180
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5276 11257 5304 11290
rect 5262 11248 5318 11257
rect 5262 11183 5318 11192
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5276 10266 5304 10678
rect 5368 10606 5396 10950
rect 5460 10742 5488 11562
rect 5552 11218 5580 12038
rect 5644 11898 5672 12174
rect 5736 12158 5856 12186
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5736 11830 5764 12158
rect 5951 11996 6259 12005
rect 5951 11994 5957 11996
rect 6013 11994 6037 11996
rect 6093 11994 6117 11996
rect 6173 11994 6197 11996
rect 6253 11994 6259 11996
rect 6013 11942 6015 11994
rect 6195 11942 6197 11994
rect 5951 11940 5957 11942
rect 6013 11940 6037 11942
rect 6093 11940 6117 11942
rect 6173 11940 6197 11942
rect 6253 11940 6259 11942
rect 5951 11931 6259 11940
rect 6288 11898 6316 12242
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 5724 11824 5776 11830
rect 5724 11766 5776 11772
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 11286 6408 11494
rect 6368 11280 6420 11286
rect 6368 11222 6420 11228
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5736 10810 5764 11086
rect 5816 11008 5868 11014
rect 5816 10950 5868 10956
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5828 10742 5856 10950
rect 5951 10908 6259 10917
rect 5951 10906 5957 10908
rect 6013 10906 6037 10908
rect 6093 10906 6117 10908
rect 6173 10906 6197 10908
rect 6253 10906 6259 10908
rect 6013 10854 6015 10906
rect 6195 10854 6197 10906
rect 5951 10852 5957 10854
rect 6013 10852 6037 10854
rect 6093 10852 6117 10854
rect 6173 10852 6197 10854
rect 6253 10852 6259 10854
rect 5951 10843 6259 10852
rect 5448 10736 5500 10742
rect 5448 10678 5500 10684
rect 5816 10736 5868 10742
rect 6472 10690 6500 13126
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7208 11694 7236 12038
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 6564 10810 6592 11630
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 5816 10678 5868 10684
rect 5828 10606 5856 10678
rect 6380 10674 6500 10690
rect 6368 10668 6500 10674
rect 6420 10662 6500 10668
rect 6368 10610 6420 10616
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 10266 5396 10406
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5460 10130 5488 10474
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5276 9518 5304 9862
rect 5644 9518 5672 9862
rect 5951 9820 6259 9829
rect 5951 9818 5957 9820
rect 6013 9818 6037 9820
rect 6093 9818 6117 9820
rect 6173 9818 6197 9820
rect 6253 9818 6259 9820
rect 6013 9766 6015 9818
rect 6195 9766 6197 9818
rect 5951 9764 5957 9766
rect 6013 9764 6037 9766
rect 6093 9764 6117 9766
rect 6173 9764 6197 9766
rect 6253 9764 6259 9766
rect 5951 9755 6259 9764
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5276 8634 5304 9454
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5552 9110 5580 9318
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 3896 6866 3924 7142
rect 4100 7100 4408 7109
rect 4100 7098 4106 7100
rect 4162 7098 4186 7100
rect 4242 7098 4266 7100
rect 4322 7098 4346 7100
rect 4402 7098 4408 7100
rect 4162 7046 4164 7098
rect 4344 7046 4346 7098
rect 4100 7044 4106 7046
rect 4162 7044 4186 7046
rect 4242 7044 4266 7046
rect 4322 7044 4346 7046
rect 4402 7044 4408 7046
rect 4100 7035 4408 7044
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3804 6202 3832 6802
rect 4540 6798 4568 7142
rect 4724 6934 4752 7278
rect 4908 7206 4936 7822
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 5368 7002 5396 7210
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4436 6656 4488 6662
rect 4436 6598 4488 6604
rect 4172 6458 4200 6598
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4448 6254 4476 6598
rect 4540 6458 4568 6734
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4540 6254 4568 6394
rect 4724 6254 4752 6870
rect 5552 6390 5580 9046
rect 5644 8566 5672 9454
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6288 9110 6316 9318
rect 6276 9104 6328 9110
rect 6380 9081 6408 10610
rect 6932 10606 6960 10950
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6656 10266 6684 10542
rect 6828 10532 6880 10538
rect 6828 10474 6880 10480
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6840 9994 6868 10474
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6460 9512 6512 9518
rect 6840 9500 6868 9930
rect 7104 9512 7156 9518
rect 6840 9472 7104 9500
rect 6460 9454 6512 9460
rect 7104 9454 7156 9460
rect 6276 9046 6328 9052
rect 6366 9072 6422 9081
rect 6366 9007 6422 9016
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5632 8560 5684 8566
rect 5632 8502 5684 8508
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5644 8022 5672 8230
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5736 6662 5764 8842
rect 5828 7818 5856 8910
rect 5951 8732 6259 8741
rect 5951 8730 5957 8732
rect 6013 8730 6037 8732
rect 6093 8730 6117 8732
rect 6173 8730 6197 8732
rect 6253 8730 6259 8732
rect 6013 8678 6015 8730
rect 6195 8678 6197 8730
rect 5951 8676 5957 8678
rect 6013 8676 6037 8678
rect 6093 8676 6117 8678
rect 6173 8676 6197 8678
rect 6253 8676 6259 8678
rect 5951 8667 6259 8676
rect 6380 8498 6408 9007
rect 6472 8634 6500 9454
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6564 8430 6592 9318
rect 7208 9178 7236 9386
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7300 9110 7328 12378
rect 7392 12102 7420 14554
rect 7576 14482 7604 14758
rect 7802 14716 8110 14725
rect 7802 14714 7808 14716
rect 7864 14714 7888 14716
rect 7944 14714 7968 14716
rect 8024 14714 8048 14716
rect 8104 14714 8110 14716
rect 7864 14662 7866 14714
rect 8046 14662 8048 14714
rect 7802 14660 7808 14662
rect 7864 14660 7888 14662
rect 7944 14660 7968 14662
rect 8024 14660 8048 14662
rect 8104 14660 8110 14662
rect 7802 14651 8110 14660
rect 8404 14618 8432 14894
rect 8484 14884 8536 14890
rect 8484 14826 8536 14832
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 7576 13734 7604 14418
rect 8312 14074 8340 14418
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 7564 13728 7616 13734
rect 7564 13670 7616 13676
rect 7802 13628 8110 13637
rect 7802 13626 7808 13628
rect 7864 13626 7888 13628
rect 7944 13626 7968 13628
rect 8024 13626 8048 13628
rect 8104 13626 8110 13628
rect 7864 13574 7866 13626
rect 8046 13574 8048 13626
rect 7802 13572 7808 13574
rect 7864 13572 7888 13574
rect 7944 13572 7968 13574
rect 8024 13572 8048 13574
rect 8104 13572 8110 13574
rect 7802 13563 8110 13572
rect 8496 13326 8524 14826
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8588 13274 8616 14010
rect 8956 13938 8984 14758
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8680 13394 8708 13806
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7668 12782 7696 13126
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7576 12306 7604 12582
rect 7802 12540 8110 12549
rect 7802 12538 7808 12540
rect 7864 12538 7888 12540
rect 7944 12538 7968 12540
rect 8024 12538 8048 12540
rect 8104 12538 8110 12540
rect 7864 12486 7866 12538
rect 8046 12486 8048 12538
rect 7802 12484 7808 12486
rect 7864 12484 7888 12486
rect 7944 12484 7968 12486
rect 8024 12484 8048 12486
rect 8104 12484 8110 12486
rect 7802 12475 8110 12484
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7392 11694 7420 12038
rect 7484 11898 7512 12242
rect 8496 12238 8524 13262
rect 8588 13246 8708 13274
rect 8680 13190 8708 13246
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7668 11694 7696 12106
rect 8128 11694 8156 12106
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11694 8248 12038
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 7802 11452 8110 11461
rect 7802 11450 7808 11452
rect 7864 11450 7888 11452
rect 7944 11450 7968 11452
rect 8024 11450 8048 11452
rect 8104 11450 8110 11452
rect 7864 11398 7866 11450
rect 8046 11398 8048 11450
rect 7802 11396 7808 11398
rect 7864 11396 7888 11398
rect 7944 11396 7968 11398
rect 8024 11396 8048 11398
rect 8104 11396 8110 11398
rect 7802 11387 8110 11396
rect 8312 11218 8340 11562
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8312 10810 8340 11154
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 7484 9518 7512 10542
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7802 10364 8110 10373
rect 7802 10362 7808 10364
rect 7864 10362 7888 10364
rect 7944 10362 7968 10364
rect 8024 10362 8048 10364
rect 8104 10362 8110 10364
rect 7864 10310 7866 10362
rect 8046 10310 8048 10362
rect 7802 10308 7808 10310
rect 7864 10308 7888 10310
rect 7944 10308 7968 10310
rect 8024 10308 8048 10310
rect 8104 10308 8110 10310
rect 7802 10299 8110 10308
rect 8220 9722 8248 10406
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 7944 9518 7972 9658
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7564 9512 7616 9518
rect 7932 9512 7984 9518
rect 7564 9454 7616 9460
rect 7668 9460 7932 9466
rect 7668 9454 7984 9460
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7392 7954 7420 8366
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 5816 7812 5868 7818
rect 5816 7754 5868 7760
rect 5828 7342 5856 7754
rect 5951 7644 6259 7653
rect 5951 7642 5957 7644
rect 6013 7642 6037 7644
rect 6093 7642 6117 7644
rect 6173 7642 6197 7644
rect 6253 7642 6259 7644
rect 6013 7590 6015 7642
rect 6195 7590 6197 7642
rect 5951 7588 5957 7590
rect 6013 7588 6037 7590
rect 6093 7588 6117 7590
rect 6173 7588 6197 7590
rect 6253 7588 6259 7590
rect 5951 7579 6259 7588
rect 6368 7472 6420 7478
rect 6368 7414 6420 7420
rect 7484 7426 7512 9454
rect 7576 9382 7604 9454
rect 7668 9450 7972 9454
rect 7656 9444 7972 9450
rect 7708 9438 7972 9444
rect 7656 9386 7708 9392
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7576 8838 7604 9318
rect 7802 9276 8110 9285
rect 7802 9274 7808 9276
rect 7864 9274 7888 9276
rect 7944 9274 7968 9276
rect 8024 9274 8048 9276
rect 8104 9274 8110 9276
rect 7864 9222 7866 9274
rect 8046 9222 8048 9274
rect 7802 9220 7808 9222
rect 7864 9220 7888 9222
rect 7944 9220 7968 9222
rect 8024 9220 8048 9222
rect 8104 9220 8110 9222
rect 7802 9211 8110 9220
rect 8404 9178 8432 10542
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 7802 8188 8110 8197
rect 7802 8186 7808 8188
rect 7864 8186 7888 8188
rect 7944 8186 7968 8188
rect 8024 8186 8048 8188
rect 8104 8186 8110 8188
rect 7864 8134 7866 8186
rect 8046 8134 8048 8186
rect 7802 8132 7808 8134
rect 7864 8132 7888 8134
rect 7944 8132 7968 8134
rect 8024 8132 8048 8134
rect 8104 8132 8110 8134
rect 7802 8123 8110 8132
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7668 7546 7696 7890
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 6380 6866 6408 7414
rect 7484 7398 7696 7426
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5828 6338 5856 6802
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 5951 6556 6259 6565
rect 5951 6554 5957 6556
rect 6013 6554 6037 6556
rect 6093 6554 6117 6556
rect 6173 6554 6197 6556
rect 6253 6554 6259 6556
rect 6013 6502 6015 6554
rect 6195 6502 6197 6554
rect 5951 6500 5957 6502
rect 6013 6500 6037 6502
rect 6093 6500 6117 6502
rect 6173 6500 6197 6502
rect 6253 6500 6259 6502
rect 5951 6491 6259 6500
rect 5828 6310 6040 6338
rect 6012 6254 6040 6310
rect 6288 6254 6316 6598
rect 6380 6390 6408 6802
rect 6656 6390 6684 6802
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6748 6458 6776 6666
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6368 6384 6420 6390
rect 6368 6326 6420 6332
rect 6644 6384 6696 6390
rect 6644 6326 6696 6332
rect 4436 6248 4488 6254
rect 3804 6174 4016 6202
rect 4436 6190 4488 6196
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3896 5914 3924 6054
rect 3988 5914 4016 6174
rect 4100 6012 4408 6021
rect 4100 6010 4106 6012
rect 4162 6010 4186 6012
rect 4242 6010 4266 6012
rect 4322 6010 4346 6012
rect 4402 6010 4408 6012
rect 4162 5958 4164 6010
rect 4344 5958 4346 6010
rect 4100 5956 4106 5958
rect 4162 5956 4186 5958
rect 4242 5956 4266 5958
rect 4322 5956 4346 5958
rect 4402 5956 4408 5958
rect 4100 5947 4408 5956
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3700 5840 3752 5846
rect 3700 5782 3752 5788
rect 4724 5778 4752 6190
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 5778 5764 6054
rect 6012 5914 6040 6190
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3712 5098 3740 5510
rect 4724 5370 4752 5714
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 6012 5534 6040 5714
rect 6104 5710 6132 6190
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6564 5794 6592 5850
rect 6380 5778 6592 5794
rect 6656 5778 6684 6054
rect 6368 5772 6592 5778
rect 6420 5766 6592 5772
rect 6644 5772 6696 5778
rect 6368 5714 6420 5720
rect 6644 5714 6696 5720
rect 6748 5710 6776 6122
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6840 5914 6868 6054
rect 7392 5914 7420 6190
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7484 5778 7512 7210
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 7002 7604 7142
rect 7668 7002 7696 7398
rect 8220 7342 8248 8230
rect 7748 7336 7800 7342
rect 8208 7336 8260 7342
rect 7838 7304 7894 7313
rect 7800 7284 7838 7290
rect 7748 7278 7838 7284
rect 7760 7262 7838 7278
rect 8208 7278 8260 7284
rect 7838 7239 7894 7248
rect 7802 7100 8110 7109
rect 7802 7098 7808 7100
rect 7864 7098 7888 7100
rect 7944 7098 7968 7100
rect 8024 7098 8048 7100
rect 8104 7098 8110 7100
rect 7864 7046 7866 7098
rect 8046 7046 8048 7098
rect 7802 7044 7808 7046
rect 7864 7044 7888 7046
rect 7944 7044 7968 7046
rect 8024 7044 8048 7046
rect 8104 7044 8110 7046
rect 7802 7035 8110 7044
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 7852 6118 7880 6258
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7802 6012 8110 6021
rect 7802 6010 7808 6012
rect 7864 6010 7888 6012
rect 7944 6010 7968 6012
rect 8024 6010 8048 6012
rect 8104 6010 8110 6012
rect 7864 5958 7866 6010
rect 8046 5958 8048 6010
rect 7802 5956 7808 5958
rect 7864 5956 7888 5958
rect 7944 5956 7968 5958
rect 8024 5956 8048 5958
rect 8104 5956 8110 5958
rect 7802 5947 8110 5956
rect 8404 5846 8432 9114
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8496 6866 8524 8230
rect 8588 7954 8616 13126
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8772 12102 8800 12582
rect 8864 12306 8892 13330
rect 9048 13258 9076 14758
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 8852 12300 8904 12306
rect 8852 12242 8904 12248
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 9048 11898 9076 12582
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8680 11354 8708 11630
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8772 8430 8800 9590
rect 8864 8430 8892 10610
rect 8956 8430 8984 11154
rect 9048 11150 9076 11834
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 9140 10266 9168 11494
rect 9324 11098 9352 12854
rect 9416 12170 9444 14554
rect 9508 13938 9536 14758
rect 10152 14618 10180 14894
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 9653 14172 9961 14181
rect 9653 14170 9659 14172
rect 9715 14170 9739 14172
rect 9795 14170 9819 14172
rect 9875 14170 9899 14172
rect 9955 14170 9961 14172
rect 9715 14118 9717 14170
rect 9897 14118 9899 14170
rect 9653 14116 9659 14118
rect 9715 14116 9739 14118
rect 9795 14116 9819 14118
rect 9875 14116 9899 14118
rect 9955 14116 9961 14118
rect 9653 14107 9961 14116
rect 10244 14074 10272 14418
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9968 13394 9996 13806
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9508 12306 9536 13126
rect 9653 13084 9961 13093
rect 9653 13082 9659 13084
rect 9715 13082 9739 13084
rect 9795 13082 9819 13084
rect 9875 13082 9899 13084
rect 9955 13082 9961 13084
rect 9715 13030 9717 13082
rect 9897 13030 9899 13082
rect 9653 13028 9659 13030
rect 9715 13028 9739 13030
rect 9795 13028 9819 13030
rect 9875 13028 9899 13030
rect 9955 13028 9961 13030
rect 9653 13019 9961 13028
rect 10060 12714 10088 13126
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10152 12442 10180 13262
rect 10336 12850 10364 14418
rect 10428 13870 10456 14758
rect 11348 13938 11376 14758
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9416 11762 9444 12106
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9508 11778 9536 12038
rect 9653 11996 9961 12005
rect 9653 11994 9659 11996
rect 9715 11994 9739 11996
rect 9795 11994 9819 11996
rect 9875 11994 9899 11996
rect 9955 11994 9961 11996
rect 9715 11942 9717 11994
rect 9897 11942 9899 11994
rect 9653 11940 9659 11942
rect 9715 11940 9739 11942
rect 9795 11940 9819 11942
rect 9875 11940 9899 11942
rect 9955 11940 9961 11942
rect 9653 11931 9961 11940
rect 9508 11762 9628 11778
rect 9404 11756 9456 11762
rect 9508 11756 9640 11762
rect 9508 11750 9588 11756
rect 9404 11698 9456 11704
rect 9588 11698 9640 11704
rect 9416 11218 9444 11698
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9588 11620 9640 11626
rect 9508 11580 9588 11608
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9324 11070 9444 11098
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9324 10266 9352 10950
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8496 6254 8524 6802
rect 8864 6730 8892 8366
rect 9048 8294 9076 9658
rect 9140 9586 9168 9862
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9232 9178 9260 9318
rect 9324 9178 9352 9862
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9310 9072 9366 9081
rect 9310 9007 9366 9016
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9140 8430 9168 8774
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 8864 6361 8892 6666
rect 8850 6352 8906 6361
rect 8850 6287 8906 6296
rect 9048 6254 9076 7890
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 9048 5778 9076 6054
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6748 5574 6776 5646
rect 6736 5568 6788 5574
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 5276 5166 5304 5510
rect 6012 5506 6316 5534
rect 6736 5510 6788 5516
rect 7748 5568 7800 5574
rect 9140 5534 9168 6054
rect 9232 5914 9260 8434
rect 9324 7750 9352 9007
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9416 7342 9444 11070
rect 9508 9518 9536 11580
rect 9588 11562 9640 11568
rect 9692 11286 9720 11630
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9968 11218 9996 11494
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9653 10908 9961 10917
rect 9653 10906 9659 10908
rect 9715 10906 9739 10908
rect 9795 10906 9819 10908
rect 9875 10906 9899 10908
rect 9955 10906 9961 10908
rect 9715 10854 9717 10906
rect 9897 10854 9899 10906
rect 9653 10852 9659 10854
rect 9715 10852 9739 10854
rect 9795 10852 9819 10854
rect 9875 10852 9899 10854
rect 9955 10852 9961 10854
rect 9653 10843 9961 10852
rect 10060 10742 10088 11154
rect 10048 10736 10100 10742
rect 10048 10678 10100 10684
rect 10244 10690 10272 12242
rect 10336 10810 10364 12786
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10244 10662 10364 10690
rect 9653 9820 9961 9829
rect 9653 9818 9659 9820
rect 9715 9818 9739 9820
rect 9795 9818 9819 9820
rect 9875 9818 9899 9820
rect 9955 9818 9961 9820
rect 9715 9766 9717 9818
rect 9897 9766 9899 9818
rect 9653 9764 9659 9766
rect 9715 9764 9739 9766
rect 9795 9764 9819 9766
rect 9875 9764 9899 9766
rect 9955 9764 9961 9766
rect 9653 9755 9961 9764
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9508 8362 9536 9454
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 9586 9072 9642 9081
rect 9642 9042 9720 9058
rect 9642 9036 9732 9042
rect 9642 9030 9680 9036
rect 9586 9007 9642 9016
rect 9680 8978 9732 8984
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9968 8906 9996 8978
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9653 8732 9961 8741
rect 9653 8730 9659 8732
rect 9715 8730 9739 8732
rect 9795 8730 9819 8732
rect 9875 8730 9899 8732
rect 9955 8730 9961 8732
rect 9715 8678 9717 8730
rect 9897 8678 9899 8730
rect 9653 8676 9659 8678
rect 9715 8676 9739 8678
rect 9795 8676 9819 8678
rect 9875 8676 9899 8678
rect 9955 8676 9961 8678
rect 9653 8667 9961 8676
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9508 8090 9536 8298
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9653 7644 9961 7653
rect 9653 7642 9659 7644
rect 9715 7642 9739 7644
rect 9795 7642 9819 7644
rect 9875 7642 9899 7644
rect 9955 7642 9961 7644
rect 9715 7590 9717 7642
rect 9897 7590 9899 7642
rect 9653 7588 9659 7590
rect 9715 7588 9739 7590
rect 9795 7588 9819 7590
rect 9875 7588 9899 7590
rect 9955 7588 9961 7590
rect 9653 7579 9961 7588
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9508 7002 9536 7142
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9653 6556 9961 6565
rect 9653 6554 9659 6556
rect 9715 6554 9739 6556
rect 9795 6554 9819 6556
rect 9875 6554 9899 6556
rect 9955 6554 9961 6556
rect 9715 6502 9717 6554
rect 9897 6502 9899 6554
rect 9653 6500 9659 6502
rect 9715 6500 9739 6502
rect 9795 6500 9819 6502
rect 9875 6500 9899 6502
rect 9955 6500 9961 6502
rect 9653 6491 9961 6500
rect 10060 6458 10088 9114
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 10152 8430 10180 8774
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 10244 8090 10272 9046
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 7478 10272 7686
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9772 6384 9824 6390
rect 9692 6332 9772 6338
rect 9692 6326 9824 6332
rect 10046 6352 10102 6361
rect 9692 6310 9812 6326
rect 9692 6254 9720 6310
rect 10046 6287 10102 6296
rect 10060 6254 10088 6287
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 9784 5914 9812 6190
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9232 5794 9260 5850
rect 9232 5766 9536 5794
rect 7800 5516 7972 5534
rect 7748 5510 7972 5516
rect 5951 5468 6259 5477
rect 5951 5466 5957 5468
rect 6013 5466 6037 5468
rect 6093 5466 6117 5468
rect 6173 5466 6197 5468
rect 6253 5466 6259 5468
rect 6013 5414 6015 5466
rect 6195 5414 6197 5466
rect 5951 5412 5957 5414
rect 6013 5412 6037 5414
rect 6093 5412 6117 5414
rect 6173 5412 6197 5414
rect 6253 5412 6259 5414
rect 5951 5403 6259 5412
rect 6288 5370 6316 5506
rect 6748 5370 6776 5510
rect 7760 5506 7972 5510
rect 9140 5506 9352 5534
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 7944 5166 7972 5506
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 9324 5098 9352 5506
rect 9508 5166 9536 5766
rect 9653 5468 9961 5477
rect 9653 5466 9659 5468
rect 9715 5466 9739 5468
rect 9795 5466 9819 5468
rect 9875 5466 9899 5468
rect 9955 5466 9961 5468
rect 9715 5414 9717 5466
rect 9897 5414 9899 5466
rect 9653 5412 9659 5414
rect 9715 5412 9739 5414
rect 9795 5412 9819 5414
rect 9875 5412 9899 5414
rect 9955 5412 9961 5414
rect 9653 5403 9961 5412
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 3700 5092 3752 5098
rect 3700 5034 3752 5040
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 4100 4924 4408 4933
rect 4100 4922 4106 4924
rect 4162 4922 4186 4924
rect 4242 4922 4266 4924
rect 4322 4922 4346 4924
rect 4402 4922 4408 4924
rect 4162 4870 4164 4922
rect 4344 4870 4346 4922
rect 4100 4868 4106 4870
rect 4162 4868 4186 4870
rect 4242 4868 4266 4870
rect 4322 4868 4346 4870
rect 4402 4868 4408 4870
rect 4100 4859 4408 4868
rect 7802 4924 8110 4933
rect 7802 4922 7808 4924
rect 7864 4922 7888 4924
rect 7944 4922 7968 4924
rect 8024 4922 8048 4924
rect 8104 4922 8110 4924
rect 7864 4870 7866 4922
rect 8046 4870 8048 4922
rect 7802 4868 7808 4870
rect 7864 4868 7888 4870
rect 7944 4868 7968 4870
rect 8024 4868 8048 4870
rect 8104 4868 8110 4870
rect 7802 4859 8110 4868
rect 2249 4380 2557 4389
rect 2249 4378 2255 4380
rect 2311 4378 2335 4380
rect 2391 4378 2415 4380
rect 2471 4378 2495 4380
rect 2551 4378 2557 4380
rect 2311 4326 2313 4378
rect 2493 4326 2495 4378
rect 2249 4324 2255 4326
rect 2311 4324 2335 4326
rect 2391 4324 2415 4326
rect 2471 4324 2495 4326
rect 2551 4324 2557 4326
rect 2249 4315 2557 4324
rect 5951 4380 6259 4389
rect 5951 4378 5957 4380
rect 6013 4378 6037 4380
rect 6093 4378 6117 4380
rect 6173 4378 6197 4380
rect 6253 4378 6259 4380
rect 6013 4326 6015 4378
rect 6195 4326 6197 4378
rect 5951 4324 5957 4326
rect 6013 4324 6037 4326
rect 6093 4324 6117 4326
rect 6173 4324 6197 4326
rect 6253 4324 6259 4326
rect 5951 4315 6259 4324
rect 9508 4146 9536 5102
rect 9653 4380 9961 4389
rect 9653 4378 9659 4380
rect 9715 4378 9739 4380
rect 9795 4378 9819 4380
rect 9875 4378 9899 4380
rect 9955 4378 9961 4380
rect 9715 4326 9717 4378
rect 9897 4326 9899 4378
rect 9653 4324 9659 4326
rect 9715 4324 9739 4326
rect 9795 4324 9819 4326
rect 9875 4324 9899 4326
rect 9955 4324 9961 4326
rect 9653 4315 9961 4324
rect 10152 4162 10180 7414
rect 10336 7290 10364 10662
rect 10428 8090 10456 13806
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10520 7342 10548 13670
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10612 12306 10640 12582
rect 11256 12442 11284 13262
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10612 11830 10640 12242
rect 11440 12102 11468 15098
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11504 14716 11812 14725
rect 11504 14714 11510 14716
rect 11566 14714 11590 14716
rect 11646 14714 11670 14716
rect 11726 14714 11750 14716
rect 11806 14714 11812 14716
rect 11566 14662 11568 14714
rect 11748 14662 11750 14714
rect 11504 14660 11510 14662
rect 11566 14660 11590 14662
rect 11646 14660 11670 14662
rect 11726 14660 11750 14662
rect 11806 14660 11812 14662
rect 11504 14651 11812 14660
rect 11992 14618 12020 14758
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11504 13628 11812 13637
rect 11504 13626 11510 13628
rect 11566 13626 11590 13628
rect 11646 13626 11670 13628
rect 11726 13626 11750 13628
rect 11806 13626 11812 13628
rect 11566 13574 11568 13626
rect 11748 13574 11750 13626
rect 11504 13572 11510 13574
rect 11566 13572 11590 13574
rect 11646 13572 11670 13574
rect 11726 13572 11750 13574
rect 11806 13572 11812 13574
rect 11504 13563 11812 13572
rect 11900 13394 11928 13806
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11900 12714 11928 13126
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11992 12594 12020 14554
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 12084 14074 12112 14418
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12176 13870 12204 15302
rect 12452 14958 12480 15600
rect 13355 15260 13663 15269
rect 13355 15258 13361 15260
rect 13417 15258 13441 15260
rect 13497 15258 13521 15260
rect 13577 15258 13601 15260
rect 13657 15258 13663 15260
rect 13417 15206 13419 15258
rect 13599 15206 13601 15258
rect 13355 15204 13361 15206
rect 13417 15204 13441 15206
rect 13497 15204 13521 15206
rect 13577 15204 13601 15206
rect 13657 15204 13663 15206
rect 13355 15195 13663 15204
rect 12808 15088 12860 15094
rect 12808 15030 12860 15036
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12268 14006 12296 14758
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 12176 12866 12204 13806
rect 11900 12566 12020 12594
rect 12084 12838 12204 12866
rect 11504 12540 11812 12549
rect 11504 12538 11510 12540
rect 11566 12538 11590 12540
rect 11646 12538 11670 12540
rect 11726 12538 11750 12540
rect 11806 12538 11812 12540
rect 11566 12486 11568 12538
rect 11748 12486 11750 12538
rect 11504 12484 11510 12486
rect 11566 12484 11590 12486
rect 11646 12484 11670 12486
rect 11726 12484 11750 12486
rect 11806 12484 11812 12486
rect 11504 12475 11812 12484
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11900 11898 11928 12566
rect 12084 11898 12112 12838
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 12176 12306 12204 12718
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10612 11014 10640 11766
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10704 11286 10732 11562
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10704 10130 10732 11222
rect 11164 11218 11192 11494
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10888 10606 10916 11086
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11072 10674 11100 10950
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 11348 10538 11376 11494
rect 11440 10606 11468 11494
rect 11504 11452 11812 11461
rect 11504 11450 11510 11452
rect 11566 11450 11590 11452
rect 11646 11450 11670 11452
rect 11726 11450 11750 11452
rect 11806 11450 11812 11452
rect 11566 11398 11568 11450
rect 11748 11398 11750 11450
rect 11504 11396 11510 11398
rect 11566 11396 11590 11398
rect 11646 11396 11670 11398
rect 11726 11396 11750 11398
rect 11806 11396 11812 11398
rect 11504 11387 11812 11396
rect 11900 11150 11928 11834
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11992 11218 12020 11494
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11504 10364 11812 10373
rect 11504 10362 11510 10364
rect 11566 10362 11590 10364
rect 11646 10362 11670 10364
rect 11726 10362 11750 10364
rect 11806 10362 11812 10364
rect 11566 10310 11568 10362
rect 11748 10310 11750 10362
rect 11504 10308 11510 10310
rect 11566 10308 11590 10310
rect 11646 10308 11670 10310
rect 11726 10308 11750 10310
rect 11806 10308 11812 10310
rect 11504 10299 11812 10308
rect 11992 10130 12020 11154
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10612 9042 10640 9318
rect 10704 9178 10732 10066
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10612 7954 10640 8978
rect 10704 8906 10732 9114
rect 10796 9042 10824 9386
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10888 9042 10916 9318
rect 11440 9178 11468 9386
rect 11532 9382 11560 9998
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11504 9276 11812 9285
rect 11504 9274 11510 9276
rect 11566 9274 11590 9276
rect 11646 9274 11670 9276
rect 11726 9274 11750 9276
rect 11806 9274 11812 9276
rect 11566 9222 11568 9274
rect 11748 9222 11750 9274
rect 11504 9220 11510 9222
rect 11566 9220 11590 9222
rect 11646 9220 11670 9222
rect 11726 9220 11750 9222
rect 11806 9220 11812 9222
rect 11504 9211 11812 9220
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11992 9042 12020 9862
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11256 8634 11284 8842
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11504 8188 11812 8197
rect 11504 8186 11510 8188
rect 11566 8186 11590 8188
rect 11646 8186 11670 8188
rect 11726 8186 11750 8188
rect 11806 8186 11812 8188
rect 11566 8134 11568 8186
rect 11748 8134 11750 8186
rect 11504 8132 11510 8134
rect 11566 8132 11590 8134
rect 11646 8132 11670 8134
rect 11726 8132 11750 8134
rect 11806 8132 11812 8134
rect 11504 8123 11812 8132
rect 11992 7954 12020 8230
rect 12084 8022 12112 11834
rect 12268 9450 12296 13942
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12360 10713 12388 13262
rect 12452 11150 12480 14214
rect 12728 13530 12756 14758
rect 12820 14482 12848 15030
rect 13740 14958 13768 15600
rect 15028 14958 15056 15600
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 13188 14618 13216 14894
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 12820 13938 12848 14418
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12636 12918 12664 13330
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12636 11218 12664 12854
rect 12728 11354 12756 13466
rect 12912 12764 12940 14418
rect 13004 13274 13032 14418
rect 13096 14074 13124 14418
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13280 13870 13308 14758
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13355 14172 13663 14181
rect 13355 14170 13361 14172
rect 13417 14170 13441 14172
rect 13497 14170 13521 14172
rect 13577 14170 13601 14172
rect 13657 14170 13663 14172
rect 13417 14118 13419 14170
rect 13599 14118 13601 14170
rect 13355 14116 13361 14118
rect 13417 14116 13441 14118
rect 13497 14116 13521 14118
rect 13577 14116 13601 14118
rect 13657 14116 13663 14118
rect 13355 14107 13663 14116
rect 13740 14074 13768 14350
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13832 13954 13860 14758
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 13740 13926 13860 13954
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13004 13246 13124 13274
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 13004 12986 13032 13126
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 12992 12776 13044 12782
rect 12912 12744 12992 12764
rect 13044 12744 13046 12753
rect 12912 12736 12990 12744
rect 13096 12714 13124 13246
rect 12990 12679 13046 12688
rect 13084 12708 13136 12714
rect 13084 12650 13136 12656
rect 13096 12442 13124 12650
rect 13280 12458 13308 13670
rect 13372 13326 13400 13670
rect 13740 13462 13768 13926
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 13530 13860 13806
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13728 13456 13780 13462
rect 13780 13404 13860 13410
rect 13728 13398 13860 13404
rect 13740 13382 13860 13398
rect 14016 13394 14044 14214
rect 14200 13394 14228 14758
rect 15206 14716 15514 14725
rect 15206 14714 15212 14716
rect 15268 14714 15292 14716
rect 15348 14714 15372 14716
rect 15428 14714 15452 14716
rect 15508 14714 15514 14716
rect 15268 14662 15270 14714
rect 15450 14662 15452 14714
rect 15206 14660 15212 14662
rect 15268 14660 15292 14662
rect 15348 14660 15372 14662
rect 15428 14660 15452 14662
rect 15508 14660 15514 14662
rect 15206 14651 15514 14660
rect 15014 14512 15070 14521
rect 15014 14447 15016 14456
rect 15068 14447 15070 14456
rect 15016 14418 15068 14424
rect 15028 13938 15056 14418
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 15206 13628 15514 13637
rect 15206 13626 15212 13628
rect 15268 13626 15292 13628
rect 15348 13626 15372 13628
rect 15428 13626 15452 13628
rect 15508 13626 15514 13628
rect 15268 13574 15270 13626
rect 15450 13574 15452 13626
rect 15206 13572 15212 13574
rect 15268 13572 15292 13574
rect 15348 13572 15372 13574
rect 15428 13572 15452 13574
rect 15508 13572 15514 13574
rect 15206 13563 15514 13572
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13355 13084 13663 13093
rect 13355 13082 13361 13084
rect 13417 13082 13441 13084
rect 13497 13082 13521 13084
rect 13577 13082 13601 13084
rect 13657 13082 13663 13084
rect 13417 13030 13419 13082
rect 13599 13030 13601 13082
rect 13355 13028 13361 13030
rect 13417 13028 13441 13030
rect 13497 13028 13521 13030
rect 13577 13028 13601 13030
rect 13657 13028 13663 13030
rect 13355 13019 13663 13028
rect 13740 12986 13768 13262
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13464 12617 13492 12650
rect 13544 12640 13596 12646
rect 13450 12608 13506 12617
rect 13740 12628 13768 12718
rect 13596 12600 13768 12628
rect 13544 12582 13596 12588
rect 13450 12543 13506 12552
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13188 12430 13308 12458
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12346 10704 12402 10713
rect 12346 10639 12402 10648
rect 12452 10282 12480 11086
rect 12360 10254 12480 10282
rect 12256 9444 12308 9450
rect 12256 9386 12308 9392
rect 12360 8566 12388 10254
rect 12636 10130 12664 11154
rect 12912 10810 12940 11154
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12452 9654 12480 10066
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12438 9072 12494 9081
rect 12636 9042 12664 10066
rect 13004 9602 13032 11154
rect 13188 11054 13216 12430
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13280 11218 13308 12242
rect 13355 11996 13663 12005
rect 13355 11994 13361 11996
rect 13417 11994 13441 11996
rect 13497 11994 13521 11996
rect 13577 11994 13601 11996
rect 13657 11994 13663 11996
rect 13417 11942 13419 11994
rect 13599 11942 13601 11994
rect 13355 11940 13361 11942
rect 13417 11940 13441 11942
rect 13497 11940 13521 11942
rect 13577 11940 13601 11942
rect 13657 11940 13663 11942
rect 13355 11931 13663 11940
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13648 11054 13676 11086
rect 13832 11054 13860 13382
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 13924 12306 13952 13126
rect 14200 12792 14228 13126
rect 14188 12786 14240 12792
rect 14476 12782 14504 13330
rect 14188 12728 14240 12734
rect 14280 12776 14332 12782
rect 14464 12776 14516 12782
rect 14280 12718 14332 12724
rect 14462 12744 14464 12753
rect 14516 12744 14518 12753
rect 14004 12640 14056 12646
rect 14002 12608 14004 12617
rect 14056 12608 14058 12617
rect 14002 12543 14058 12552
rect 14292 12442 14320 12718
rect 14462 12679 14518 12688
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 13188 11026 13308 11054
rect 13648 11026 13768 11054
rect 13832 11026 13952 11054
rect 12912 9574 13032 9602
rect 12912 9178 12940 9574
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 12900 9172 12952 9178
rect 12820 9132 12900 9160
rect 12438 9007 12440 9016
rect 12492 9007 12494 9016
rect 12624 9036 12676 9042
rect 12440 8978 12492 8984
rect 12624 8978 12676 8984
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 10244 7262 10364 7290
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10612 7274 10640 7890
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10600 7268 10652 7274
rect 10244 6390 10272 7262
rect 10600 7210 10652 7216
rect 10980 6458 11008 7482
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 11072 7002 11100 7210
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 10244 6186 10272 6326
rect 11256 6254 11284 7142
rect 11348 6474 11376 7890
rect 11888 7880 11940 7886
rect 12360 7834 12388 8502
rect 12636 8430 12664 8978
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12636 8022 12664 8366
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 11888 7822 11940 7828
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11440 6934 11468 7278
rect 11504 7100 11812 7109
rect 11504 7098 11510 7100
rect 11566 7098 11590 7100
rect 11646 7098 11670 7100
rect 11726 7098 11750 7100
rect 11806 7098 11812 7100
rect 11566 7046 11568 7098
rect 11748 7046 11750 7098
rect 11504 7044 11510 7046
rect 11566 7044 11590 7046
rect 11646 7044 11670 7046
rect 11726 7044 11750 7046
rect 11806 7044 11812 7046
rect 11504 7035 11812 7044
rect 11428 6928 11480 6934
rect 11900 6914 11928 7822
rect 12268 7806 12388 7834
rect 12268 7546 12296 7806
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12162 7304 12218 7313
rect 12162 7239 12218 7248
rect 11900 6886 12112 6914
rect 11428 6870 11480 6876
rect 11348 6446 11468 6474
rect 11440 6254 11468 6446
rect 12084 6390 12112 6886
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 10336 5710 10364 6054
rect 11164 5710 11192 6054
rect 11348 5914 11376 6054
rect 11504 6012 11812 6021
rect 11504 6010 11510 6012
rect 11566 6010 11590 6012
rect 11646 6010 11670 6012
rect 11726 6010 11750 6012
rect 11806 6010 11812 6012
rect 11566 5958 11568 6010
rect 11748 5958 11750 6010
rect 11504 5956 11510 5958
rect 11566 5956 11590 5958
rect 11646 5956 11670 5958
rect 11726 5956 11750 5958
rect 11806 5956 11812 5958
rect 11504 5947 11812 5956
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 12084 5778 12112 6326
rect 12176 5914 12204 7239
rect 12268 7206 12296 7482
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12360 6254 12388 7686
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12452 7002 12480 7278
rect 12544 7274 12572 7890
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12532 7268 12584 7274
rect 12532 7210 12584 7216
rect 12544 7002 12572 7210
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12452 6610 12480 6938
rect 12636 6730 12664 7686
rect 12728 7206 12756 7822
rect 12820 7818 12848 9132
rect 12900 9114 12952 9120
rect 13004 8974 13032 9454
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 13096 9178 13124 9318
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 12912 8634 12940 8910
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 13004 6866 13032 8910
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 13188 8022 13216 8366
rect 13176 8016 13228 8022
rect 13176 7958 13228 7964
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 13096 7546 13124 7890
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 13280 7313 13308 11026
rect 13355 10908 13663 10917
rect 13355 10906 13361 10908
rect 13417 10906 13441 10908
rect 13497 10906 13521 10908
rect 13577 10906 13601 10908
rect 13657 10906 13663 10908
rect 13417 10854 13419 10906
rect 13599 10854 13601 10906
rect 13355 10852 13361 10854
rect 13417 10852 13441 10854
rect 13497 10852 13521 10854
rect 13577 10852 13601 10854
rect 13657 10852 13663 10854
rect 13355 10843 13663 10852
rect 13740 10810 13768 11026
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13924 10606 13952 11026
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 14016 10606 14044 10950
rect 14108 10742 14136 12174
rect 14292 11218 14320 12378
rect 14476 12238 14504 12582
rect 15028 12374 15056 12650
rect 15206 12540 15514 12549
rect 15206 12538 15212 12540
rect 15268 12538 15292 12540
rect 15348 12538 15372 12540
rect 15428 12538 15452 12540
rect 15508 12538 15514 12540
rect 15268 12486 15270 12538
rect 15450 12486 15452 12538
rect 15206 12484 15212 12486
rect 15268 12484 15292 12486
rect 15348 12484 15372 12486
rect 15428 12484 15452 12486
rect 15508 12484 15514 12486
rect 15206 12475 15514 12484
rect 15016 12368 15068 12374
rect 15014 12336 15016 12345
rect 15068 12336 15070 12345
rect 15014 12271 15070 12280
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 15206 11452 15514 11461
rect 15206 11450 15212 11452
rect 15268 11450 15292 11452
rect 15348 11450 15372 11452
rect 15428 11450 15452 11452
rect 15508 11450 15514 11452
rect 15268 11398 15270 11450
rect 15450 11398 15452 11450
rect 15206 11396 15212 11398
rect 15268 11396 15292 11398
rect 15348 11396 15372 11398
rect 15428 11396 15452 11398
rect 15508 11396 15514 11398
rect 15206 11387 15514 11396
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 14292 10810 14320 11154
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14186 10704 14242 10713
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 13740 10470 13768 10542
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13355 9820 13663 9829
rect 13355 9818 13361 9820
rect 13417 9818 13441 9820
rect 13497 9818 13521 9820
rect 13577 9818 13601 9820
rect 13657 9818 13663 9820
rect 13417 9766 13419 9818
rect 13599 9766 13601 9818
rect 13355 9764 13361 9766
rect 13417 9764 13441 9766
rect 13497 9764 13521 9766
rect 13577 9764 13601 9766
rect 13657 9764 13663 9766
rect 13355 9755 13663 9764
rect 13355 8732 13663 8741
rect 13355 8730 13361 8732
rect 13417 8730 13441 8732
rect 13497 8730 13521 8732
rect 13577 8730 13601 8732
rect 13657 8730 13663 8732
rect 13417 8678 13419 8730
rect 13599 8678 13601 8730
rect 13355 8676 13361 8678
rect 13417 8676 13441 8678
rect 13497 8676 13521 8678
rect 13577 8676 13601 8678
rect 13657 8676 13663 8678
rect 13355 8667 13663 8676
rect 13924 8294 13952 10542
rect 14108 9586 14136 10678
rect 14186 10639 14242 10648
rect 14200 10606 14228 10639
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14096 8832 14148 8838
rect 14200 8786 14228 10542
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 14292 9450 14320 10406
rect 14568 9518 14596 10746
rect 14936 10713 14964 10950
rect 14922 10704 14978 10713
rect 14922 10639 14978 10648
rect 14936 10538 14964 10639
rect 14924 10532 14976 10538
rect 14924 10474 14976 10480
rect 15206 10364 15514 10373
rect 15206 10362 15212 10364
rect 15268 10362 15292 10364
rect 15348 10362 15372 10364
rect 15428 10362 15452 10364
rect 15508 10362 15514 10364
rect 15268 10310 15270 10362
rect 15450 10310 15452 10362
rect 15206 10308 15212 10310
rect 15268 10308 15292 10310
rect 15348 10308 15372 10310
rect 15428 10308 15452 10310
rect 15508 10308 15514 10310
rect 15206 10299 15514 10308
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14148 8780 14228 8786
rect 14096 8774 14228 8780
rect 14108 8758 14228 8774
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13355 7644 13663 7653
rect 13355 7642 13361 7644
rect 13417 7642 13441 7644
rect 13497 7642 13521 7644
rect 13577 7642 13601 7644
rect 13657 7642 13663 7644
rect 13417 7590 13419 7642
rect 13599 7590 13601 7642
rect 13355 7588 13361 7590
rect 13417 7588 13441 7590
rect 13497 7588 13521 7590
rect 13577 7588 13601 7590
rect 13657 7588 13663 7590
rect 13355 7579 13663 7588
rect 13924 7342 13952 8230
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14016 7342 14044 7686
rect 14200 7342 14228 8758
rect 14292 8430 14320 9386
rect 14568 9178 14596 9454
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 15028 8838 15056 9386
rect 15206 9276 15514 9285
rect 15206 9274 15212 9276
rect 15268 9274 15292 9276
rect 15348 9274 15372 9276
rect 15428 9274 15452 9276
rect 15508 9274 15514 9276
rect 15268 9222 15270 9274
rect 15450 9222 15452 9274
rect 15206 9220 15212 9222
rect 15268 9220 15292 9222
rect 15348 9220 15372 9222
rect 15428 9220 15452 9222
rect 15508 9220 15514 9222
rect 15206 9211 15514 9220
rect 15016 8832 15068 8838
rect 15014 8800 15016 8809
rect 15068 8800 15070 8809
rect 15014 8735 15070 8744
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 13912 7336 13964 7342
rect 13266 7304 13322 7313
rect 13912 7278 13964 7284
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 13266 7239 13322 7248
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13648 6866 13676 7142
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12716 6656 12768 6662
rect 12452 6604 12716 6610
rect 12452 6598 12768 6604
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12452 6582 12756 6598
rect 12452 6390 12480 6582
rect 12440 6384 12492 6390
rect 12440 6326 12492 6332
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 12544 5778 12572 6054
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 10336 5370 10364 5646
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 11624 5166 11652 5510
rect 12728 5370 12756 6582
rect 12820 6118 12848 6598
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 11612 5160 11664 5166
rect 11612 5102 11664 5108
rect 11504 4924 11812 4933
rect 11504 4922 11510 4924
rect 11566 4922 11590 4924
rect 11646 4922 11670 4924
rect 11726 4922 11750 4924
rect 11806 4922 11812 4924
rect 11566 4870 11568 4922
rect 11748 4870 11750 4922
rect 11504 4868 11510 4870
rect 11566 4868 11590 4870
rect 11646 4868 11670 4870
rect 11726 4868 11750 4870
rect 11806 4868 11812 4870
rect 11504 4859 11812 4868
rect 12820 4282 12848 6054
rect 13004 5710 13032 6802
rect 13355 6556 13663 6565
rect 13355 6554 13361 6556
rect 13417 6554 13441 6556
rect 13497 6554 13521 6556
rect 13577 6554 13601 6556
rect 13657 6554 13663 6556
rect 13417 6502 13419 6554
rect 13599 6502 13601 6554
rect 13355 6500 13361 6502
rect 13417 6500 13441 6502
rect 13497 6500 13521 6502
rect 13577 6500 13601 6502
rect 13657 6500 13663 6502
rect 13355 6491 13663 6500
rect 14292 6458 14320 8366
rect 15206 8188 15514 8197
rect 15206 8186 15212 8188
rect 15268 8186 15292 8188
rect 15348 8186 15372 8188
rect 15428 8186 15452 8188
rect 15508 8186 15514 8188
rect 15268 8134 15270 8186
rect 15450 8134 15452 8186
rect 15206 8132 15212 8134
rect 15268 8132 15292 8134
rect 15348 8132 15372 8134
rect 15428 8132 15452 8134
rect 15508 8132 15514 8134
rect 15206 8123 15514 8132
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 14464 6928 14516 6934
rect 15028 6905 15056 7278
rect 15206 7100 15514 7109
rect 15206 7098 15212 7100
rect 15268 7098 15292 7100
rect 15348 7098 15372 7100
rect 15428 7098 15452 7100
rect 15508 7098 15514 7100
rect 15268 7046 15270 7098
rect 15450 7046 15452 7098
rect 15206 7044 15212 7046
rect 15268 7044 15292 7046
rect 15348 7044 15372 7046
rect 15428 7044 15452 7046
rect 15508 7044 15514 7046
rect 15206 7035 15514 7044
rect 14464 6870 14516 6876
rect 15014 6896 15070 6905
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14476 6254 14504 6870
rect 15014 6831 15016 6840
rect 15068 6831 15070 6840
rect 15016 6802 15068 6808
rect 15028 6390 15056 6802
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 13004 5234 13032 5646
rect 14476 5574 14504 6190
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14464 5568 14516 5574
rect 14462 5536 14464 5545
rect 14516 5536 14518 5545
rect 13355 5468 13663 5477
rect 14462 5471 14518 5480
rect 13355 5466 13361 5468
rect 13417 5466 13441 5468
rect 13497 5466 13521 5468
rect 13577 5466 13601 5468
rect 13657 5466 13663 5468
rect 13417 5414 13419 5466
rect 13599 5414 13601 5466
rect 13355 5412 13361 5414
rect 13417 5412 13441 5414
rect 13497 5412 13521 5414
rect 13577 5412 13601 5414
rect 13657 5412 13663 5414
rect 13355 5403 13663 5412
rect 14568 5370 14596 6054
rect 15206 6012 15514 6021
rect 15206 6010 15212 6012
rect 15268 6010 15292 6012
rect 15348 6010 15372 6012
rect 15428 6010 15452 6012
rect 15508 6010 15514 6012
rect 15268 5958 15270 6010
rect 15450 5958 15452 6010
rect 15206 5956 15212 5958
rect 15268 5956 15292 5958
rect 15348 5956 15372 5958
rect 15428 5956 15452 5958
rect 15508 5956 15514 5958
rect 15206 5947 15514 5956
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13355 4380 13663 4389
rect 13355 4378 13361 4380
rect 13417 4378 13441 4380
rect 13497 4378 13521 4380
rect 13577 4378 13601 4380
rect 13657 4378 13663 4380
rect 13417 4326 13419 4378
rect 13599 4326 13601 4378
rect 13355 4324 13361 4326
rect 13417 4324 13441 4326
rect 13497 4324 13521 4326
rect 13577 4324 13601 4326
rect 13657 4324 13663 4326
rect 13355 4315 13663 4324
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 9968 4146 10180 4162
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9956 4140 10180 4146
rect 10008 4134 10180 4140
rect 9956 4082 10008 4088
rect 4100 3836 4408 3845
rect 4100 3834 4106 3836
rect 4162 3834 4186 3836
rect 4242 3834 4266 3836
rect 4322 3834 4346 3836
rect 4402 3834 4408 3836
rect 4162 3782 4164 3834
rect 4344 3782 4346 3834
rect 4100 3780 4106 3782
rect 4162 3780 4186 3782
rect 4242 3780 4266 3782
rect 4322 3780 4346 3782
rect 4402 3780 4408 3782
rect 4100 3771 4408 3780
rect 7802 3836 8110 3845
rect 7802 3834 7808 3836
rect 7864 3834 7888 3836
rect 7944 3834 7968 3836
rect 8024 3834 8048 3836
rect 8104 3834 8110 3836
rect 7864 3782 7866 3834
rect 8046 3782 8048 3834
rect 7802 3780 7808 3782
rect 7864 3780 7888 3782
rect 7944 3780 7968 3782
rect 8024 3780 8048 3782
rect 8104 3780 8110 3782
rect 7802 3771 8110 3780
rect 11504 3836 11812 3845
rect 11504 3834 11510 3836
rect 11566 3834 11590 3836
rect 11646 3834 11670 3836
rect 11726 3834 11750 3836
rect 11806 3834 11812 3836
rect 11566 3782 11568 3834
rect 11748 3782 11750 3834
rect 11504 3780 11510 3782
rect 11566 3780 11590 3782
rect 11646 3780 11670 3782
rect 11726 3780 11750 3782
rect 11806 3780 11812 3782
rect 11504 3771 11812 3780
rect 2249 3292 2557 3301
rect 2249 3290 2255 3292
rect 2311 3290 2335 3292
rect 2391 3290 2415 3292
rect 2471 3290 2495 3292
rect 2551 3290 2557 3292
rect 2311 3238 2313 3290
rect 2493 3238 2495 3290
rect 2249 3236 2255 3238
rect 2311 3236 2335 3238
rect 2391 3236 2415 3238
rect 2471 3236 2495 3238
rect 2551 3236 2557 3238
rect 2249 3227 2557 3236
rect 5951 3292 6259 3301
rect 5951 3290 5957 3292
rect 6013 3290 6037 3292
rect 6093 3290 6117 3292
rect 6173 3290 6197 3292
rect 6253 3290 6259 3292
rect 6013 3238 6015 3290
rect 6195 3238 6197 3290
rect 5951 3236 5957 3238
rect 6013 3236 6037 3238
rect 6093 3236 6117 3238
rect 6173 3236 6197 3238
rect 6253 3236 6259 3238
rect 5951 3227 6259 3236
rect 9653 3292 9961 3301
rect 9653 3290 9659 3292
rect 9715 3290 9739 3292
rect 9795 3290 9819 3292
rect 9875 3290 9899 3292
rect 9955 3290 9961 3292
rect 9715 3238 9717 3290
rect 9897 3238 9899 3290
rect 9653 3236 9659 3238
rect 9715 3236 9739 3238
rect 9795 3236 9819 3238
rect 9875 3236 9899 3238
rect 9955 3236 9961 3238
rect 9653 3227 9961 3236
rect 4100 2748 4408 2757
rect 4100 2746 4106 2748
rect 4162 2746 4186 2748
rect 4242 2746 4266 2748
rect 4322 2746 4346 2748
rect 4402 2746 4408 2748
rect 4162 2694 4164 2746
rect 4344 2694 4346 2746
rect 4100 2692 4106 2694
rect 4162 2692 4186 2694
rect 4242 2692 4266 2694
rect 4322 2692 4346 2694
rect 4402 2692 4408 2694
rect 4100 2683 4408 2692
rect 7802 2748 8110 2757
rect 7802 2746 7808 2748
rect 7864 2746 7888 2748
rect 7944 2746 7968 2748
rect 8024 2746 8048 2748
rect 8104 2746 8110 2748
rect 7864 2694 7866 2746
rect 8046 2694 8048 2746
rect 7802 2692 7808 2694
rect 7864 2692 7888 2694
rect 7944 2692 7968 2694
rect 8024 2692 8048 2694
rect 8104 2692 8110 2694
rect 7802 2683 8110 2692
rect 11504 2748 11812 2757
rect 11504 2746 11510 2748
rect 11566 2746 11590 2748
rect 11646 2746 11670 2748
rect 11726 2746 11750 2748
rect 11806 2746 11812 2748
rect 11566 2694 11568 2746
rect 11748 2694 11750 2746
rect 11504 2692 11510 2694
rect 11566 2692 11590 2694
rect 11646 2692 11670 2694
rect 11726 2692 11750 2694
rect 11806 2692 11812 2694
rect 11504 2683 11812 2692
rect 2249 2204 2557 2213
rect 2249 2202 2255 2204
rect 2311 2202 2335 2204
rect 2391 2202 2415 2204
rect 2471 2202 2495 2204
rect 2551 2202 2557 2204
rect 2311 2150 2313 2202
rect 2493 2150 2495 2202
rect 2249 2148 2255 2150
rect 2311 2148 2335 2150
rect 2391 2148 2415 2150
rect 2471 2148 2495 2150
rect 2551 2148 2557 2150
rect 2249 2139 2557 2148
rect 5951 2204 6259 2213
rect 5951 2202 5957 2204
rect 6013 2202 6037 2204
rect 6093 2202 6117 2204
rect 6173 2202 6197 2204
rect 6253 2202 6259 2204
rect 6013 2150 6015 2202
rect 6195 2150 6197 2202
rect 5951 2148 5957 2150
rect 6013 2148 6037 2150
rect 6093 2148 6117 2150
rect 6173 2148 6197 2150
rect 6253 2148 6259 2150
rect 5951 2139 6259 2148
rect 9653 2204 9961 2213
rect 9653 2202 9659 2204
rect 9715 2202 9739 2204
rect 9795 2202 9819 2204
rect 9875 2202 9899 2204
rect 9955 2202 9961 2204
rect 9715 2150 9717 2202
rect 9897 2150 9899 2202
rect 9653 2148 9659 2150
rect 9715 2148 9739 2150
rect 9795 2148 9819 2150
rect 9875 2148 9899 2150
rect 9955 2148 9961 2150
rect 9653 2139 9961 2148
rect 4100 1660 4408 1669
rect 4100 1658 4106 1660
rect 4162 1658 4186 1660
rect 4242 1658 4266 1660
rect 4322 1658 4346 1660
rect 4402 1658 4408 1660
rect 4162 1606 4164 1658
rect 4344 1606 4346 1658
rect 4100 1604 4106 1606
rect 4162 1604 4186 1606
rect 4242 1604 4266 1606
rect 4322 1604 4346 1606
rect 4402 1604 4408 1606
rect 4100 1595 4408 1604
rect 7802 1660 8110 1669
rect 7802 1658 7808 1660
rect 7864 1658 7888 1660
rect 7944 1658 7968 1660
rect 8024 1658 8048 1660
rect 8104 1658 8110 1660
rect 7864 1606 7866 1658
rect 8046 1606 8048 1658
rect 7802 1604 7808 1606
rect 7864 1604 7888 1606
rect 7944 1604 7968 1606
rect 8024 1604 8048 1606
rect 8104 1604 8110 1606
rect 7802 1595 8110 1604
rect 11504 1660 11812 1669
rect 11504 1658 11510 1660
rect 11566 1658 11590 1660
rect 11646 1658 11670 1660
rect 11726 1658 11750 1660
rect 11806 1658 11812 1660
rect 11566 1606 11568 1658
rect 11748 1606 11750 1658
rect 11504 1604 11510 1606
rect 11566 1604 11590 1606
rect 11646 1604 11670 1606
rect 11726 1604 11750 1606
rect 11806 1604 11812 1606
rect 11504 1595 11812 1604
rect 12360 1329 12388 4218
rect 13355 3292 13663 3301
rect 13355 3290 13361 3292
rect 13417 3290 13441 3292
rect 13497 3290 13521 3292
rect 13577 3290 13601 3292
rect 13657 3290 13663 3292
rect 13417 3238 13419 3290
rect 13599 3238 13601 3290
rect 13355 3236 13361 3238
rect 13417 3236 13441 3238
rect 13497 3236 13521 3238
rect 13577 3236 13601 3238
rect 13657 3236 13663 3238
rect 13355 3227 13663 3236
rect 14568 3097 14596 5306
rect 15206 4924 15514 4933
rect 15206 4922 15212 4924
rect 15268 4922 15292 4924
rect 15348 4922 15372 4924
rect 15428 4922 15452 4924
rect 15508 4922 15514 4924
rect 15268 4870 15270 4922
rect 15450 4870 15452 4922
rect 15206 4868 15212 4870
rect 15268 4868 15292 4870
rect 15348 4868 15372 4870
rect 15428 4868 15452 4870
rect 15508 4868 15514 4870
rect 15206 4859 15514 4868
rect 15206 3836 15514 3845
rect 15206 3834 15212 3836
rect 15268 3834 15292 3836
rect 15348 3834 15372 3836
rect 15428 3834 15452 3836
rect 15508 3834 15514 3836
rect 15268 3782 15270 3834
rect 15450 3782 15452 3834
rect 15206 3780 15212 3782
rect 15268 3780 15292 3782
rect 15348 3780 15372 3782
rect 15428 3780 15452 3782
rect 15508 3780 15514 3782
rect 15206 3771 15514 3780
rect 14554 3088 14610 3097
rect 14554 3023 14610 3032
rect 15206 2748 15514 2757
rect 15206 2746 15212 2748
rect 15268 2746 15292 2748
rect 15348 2746 15372 2748
rect 15428 2746 15452 2748
rect 15508 2746 15514 2748
rect 15268 2694 15270 2746
rect 15450 2694 15452 2746
rect 15206 2692 15212 2694
rect 15268 2692 15292 2694
rect 15348 2692 15372 2694
rect 15428 2692 15452 2694
rect 15508 2692 15514 2694
rect 15206 2683 15514 2692
rect 13355 2204 13663 2213
rect 13355 2202 13361 2204
rect 13417 2202 13441 2204
rect 13497 2202 13521 2204
rect 13577 2202 13601 2204
rect 13657 2202 13663 2204
rect 13417 2150 13419 2202
rect 13599 2150 13601 2202
rect 13355 2148 13361 2150
rect 13417 2148 13441 2150
rect 13497 2148 13521 2150
rect 13577 2148 13601 2150
rect 13657 2148 13663 2150
rect 13355 2139 13663 2148
rect 15206 1660 15514 1669
rect 15206 1658 15212 1660
rect 15268 1658 15292 1660
rect 15348 1658 15372 1660
rect 15428 1658 15452 1660
rect 15508 1658 15514 1660
rect 15268 1606 15270 1658
rect 15450 1606 15452 1658
rect 15206 1604 15212 1606
rect 15268 1604 15292 1606
rect 15348 1604 15372 1606
rect 15428 1604 15452 1606
rect 15508 1604 15514 1606
rect 15206 1595 15514 1604
rect 12346 1320 12402 1329
rect 12346 1255 12402 1264
rect 2249 1116 2557 1125
rect 2249 1114 2255 1116
rect 2311 1114 2335 1116
rect 2391 1114 2415 1116
rect 2471 1114 2495 1116
rect 2551 1114 2557 1116
rect 2311 1062 2313 1114
rect 2493 1062 2495 1114
rect 2249 1060 2255 1062
rect 2311 1060 2335 1062
rect 2391 1060 2415 1062
rect 2471 1060 2495 1062
rect 2551 1060 2557 1062
rect 2249 1051 2557 1060
rect 5951 1116 6259 1125
rect 5951 1114 5957 1116
rect 6013 1114 6037 1116
rect 6093 1114 6117 1116
rect 6173 1114 6197 1116
rect 6253 1114 6259 1116
rect 6013 1062 6015 1114
rect 6195 1062 6197 1114
rect 5951 1060 5957 1062
rect 6013 1060 6037 1062
rect 6093 1060 6117 1062
rect 6173 1060 6197 1062
rect 6253 1060 6259 1062
rect 5951 1051 6259 1060
rect 9653 1116 9961 1125
rect 9653 1114 9659 1116
rect 9715 1114 9739 1116
rect 9795 1114 9819 1116
rect 9875 1114 9899 1116
rect 9955 1114 9961 1116
rect 9715 1062 9717 1114
rect 9897 1062 9899 1114
rect 9653 1060 9659 1062
rect 9715 1060 9739 1062
rect 9795 1060 9819 1062
rect 9875 1060 9899 1062
rect 9955 1060 9961 1062
rect 9653 1051 9961 1060
rect 13355 1116 13663 1125
rect 13355 1114 13361 1116
rect 13417 1114 13441 1116
rect 13497 1114 13521 1116
rect 13577 1114 13601 1116
rect 13657 1114 13663 1116
rect 13417 1062 13419 1114
rect 13599 1062 13601 1114
rect 13355 1060 13361 1062
rect 13417 1060 13441 1062
rect 13497 1060 13521 1062
rect 13577 1060 13601 1062
rect 13657 1060 13663 1062
rect 13355 1051 13663 1060
rect 4100 572 4408 581
rect 4100 570 4106 572
rect 4162 570 4186 572
rect 4242 570 4266 572
rect 4322 570 4346 572
rect 4402 570 4408 572
rect 4162 518 4164 570
rect 4344 518 4346 570
rect 4100 516 4106 518
rect 4162 516 4186 518
rect 4242 516 4266 518
rect 4322 516 4346 518
rect 4402 516 4408 518
rect 4100 507 4408 516
rect 7802 572 8110 581
rect 7802 570 7808 572
rect 7864 570 7888 572
rect 7944 570 7968 572
rect 8024 570 8048 572
rect 8104 570 8110 572
rect 7864 518 7866 570
rect 8046 518 8048 570
rect 7802 516 7808 518
rect 7864 516 7888 518
rect 7944 516 7968 518
rect 8024 516 8048 518
rect 8104 516 8110 518
rect 7802 507 8110 516
rect 11504 572 11812 581
rect 11504 570 11510 572
rect 11566 570 11590 572
rect 11646 570 11670 572
rect 11726 570 11750 572
rect 11806 570 11812 572
rect 11566 518 11568 570
rect 11748 518 11750 570
rect 11504 516 11510 518
rect 11566 516 11590 518
rect 11646 516 11670 518
rect 11726 516 11750 518
rect 11806 516 11812 518
rect 11504 507 11812 516
rect 15206 572 15514 581
rect 15206 570 15212 572
rect 15268 570 15292 572
rect 15348 570 15372 572
rect 15428 570 15452 572
rect 15508 570 15514 572
rect 15268 518 15270 570
rect 15450 518 15452 570
rect 15206 516 15212 518
rect 15268 516 15292 518
rect 15348 516 15372 518
rect 15428 516 15452 518
rect 15508 516 15514 518
rect 15206 507 15514 516
<< via2 >>
rect 2255 15258 2311 15260
rect 2335 15258 2391 15260
rect 2415 15258 2471 15260
rect 2495 15258 2551 15260
rect 2255 15206 2301 15258
rect 2301 15206 2311 15258
rect 2335 15206 2365 15258
rect 2365 15206 2377 15258
rect 2377 15206 2391 15258
rect 2415 15206 2429 15258
rect 2429 15206 2441 15258
rect 2441 15206 2471 15258
rect 2495 15206 2505 15258
rect 2505 15206 2551 15258
rect 2255 15204 2311 15206
rect 2335 15204 2391 15206
rect 2415 15204 2471 15206
rect 2495 15204 2551 15206
rect 5957 15258 6013 15260
rect 6037 15258 6093 15260
rect 6117 15258 6173 15260
rect 6197 15258 6253 15260
rect 5957 15206 6003 15258
rect 6003 15206 6013 15258
rect 6037 15206 6067 15258
rect 6067 15206 6079 15258
rect 6079 15206 6093 15258
rect 6117 15206 6131 15258
rect 6131 15206 6143 15258
rect 6143 15206 6173 15258
rect 6197 15206 6207 15258
rect 6207 15206 6253 15258
rect 5957 15204 6013 15206
rect 6037 15204 6093 15206
rect 6117 15204 6173 15206
rect 6197 15204 6253 15206
rect 2255 14170 2311 14172
rect 2335 14170 2391 14172
rect 2415 14170 2471 14172
rect 2495 14170 2551 14172
rect 2255 14118 2301 14170
rect 2301 14118 2311 14170
rect 2335 14118 2365 14170
rect 2365 14118 2377 14170
rect 2377 14118 2391 14170
rect 2415 14118 2429 14170
rect 2429 14118 2441 14170
rect 2441 14118 2471 14170
rect 2495 14118 2505 14170
rect 2505 14118 2551 14170
rect 2255 14116 2311 14118
rect 2335 14116 2391 14118
rect 2415 14116 2471 14118
rect 2495 14116 2551 14118
rect 4106 14714 4162 14716
rect 4186 14714 4242 14716
rect 4266 14714 4322 14716
rect 4346 14714 4402 14716
rect 4106 14662 4152 14714
rect 4152 14662 4162 14714
rect 4186 14662 4216 14714
rect 4216 14662 4228 14714
rect 4228 14662 4242 14714
rect 4266 14662 4280 14714
rect 4280 14662 4292 14714
rect 4292 14662 4322 14714
rect 4346 14662 4356 14714
rect 4356 14662 4402 14714
rect 4106 14660 4162 14662
rect 4186 14660 4242 14662
rect 4266 14660 4322 14662
rect 4346 14660 4402 14662
rect 2255 13082 2311 13084
rect 2335 13082 2391 13084
rect 2415 13082 2471 13084
rect 2495 13082 2551 13084
rect 2255 13030 2301 13082
rect 2301 13030 2311 13082
rect 2335 13030 2365 13082
rect 2365 13030 2377 13082
rect 2377 13030 2391 13082
rect 2415 13030 2429 13082
rect 2429 13030 2441 13082
rect 2441 13030 2471 13082
rect 2495 13030 2505 13082
rect 2505 13030 2551 13082
rect 2255 13028 2311 13030
rect 2335 13028 2391 13030
rect 2415 13028 2471 13030
rect 2495 13028 2551 13030
rect 2255 11994 2311 11996
rect 2335 11994 2391 11996
rect 2415 11994 2471 11996
rect 2495 11994 2551 11996
rect 2255 11942 2301 11994
rect 2301 11942 2311 11994
rect 2335 11942 2365 11994
rect 2365 11942 2377 11994
rect 2377 11942 2391 11994
rect 2415 11942 2429 11994
rect 2429 11942 2441 11994
rect 2441 11942 2471 11994
rect 2495 11942 2505 11994
rect 2505 11942 2551 11994
rect 2255 11940 2311 11942
rect 2335 11940 2391 11942
rect 2415 11940 2471 11942
rect 2495 11940 2551 11942
rect 2255 10906 2311 10908
rect 2335 10906 2391 10908
rect 2415 10906 2471 10908
rect 2495 10906 2551 10908
rect 2255 10854 2301 10906
rect 2301 10854 2311 10906
rect 2335 10854 2365 10906
rect 2365 10854 2377 10906
rect 2377 10854 2391 10906
rect 2415 10854 2429 10906
rect 2429 10854 2441 10906
rect 2441 10854 2471 10906
rect 2495 10854 2505 10906
rect 2505 10854 2551 10906
rect 2255 10852 2311 10854
rect 2335 10852 2391 10854
rect 2415 10852 2471 10854
rect 2495 10852 2551 10854
rect 2255 9818 2311 9820
rect 2335 9818 2391 9820
rect 2415 9818 2471 9820
rect 2495 9818 2551 9820
rect 2255 9766 2301 9818
rect 2301 9766 2311 9818
rect 2335 9766 2365 9818
rect 2365 9766 2377 9818
rect 2377 9766 2391 9818
rect 2415 9766 2429 9818
rect 2429 9766 2441 9818
rect 2441 9766 2471 9818
rect 2495 9766 2505 9818
rect 2505 9766 2551 9818
rect 2255 9764 2311 9766
rect 2335 9764 2391 9766
rect 2415 9764 2471 9766
rect 2495 9764 2551 9766
rect 2255 8730 2311 8732
rect 2335 8730 2391 8732
rect 2415 8730 2471 8732
rect 2495 8730 2551 8732
rect 2255 8678 2301 8730
rect 2301 8678 2311 8730
rect 2335 8678 2365 8730
rect 2365 8678 2377 8730
rect 2377 8678 2391 8730
rect 2415 8678 2429 8730
rect 2429 8678 2441 8730
rect 2441 8678 2471 8730
rect 2495 8678 2505 8730
rect 2505 8678 2551 8730
rect 2255 8676 2311 8678
rect 2335 8676 2391 8678
rect 2415 8676 2471 8678
rect 2495 8676 2551 8678
rect 4106 13626 4162 13628
rect 4186 13626 4242 13628
rect 4266 13626 4322 13628
rect 4346 13626 4402 13628
rect 4106 13574 4152 13626
rect 4152 13574 4162 13626
rect 4186 13574 4216 13626
rect 4216 13574 4228 13626
rect 4228 13574 4242 13626
rect 4266 13574 4280 13626
rect 4280 13574 4292 13626
rect 4292 13574 4322 13626
rect 4346 13574 4356 13626
rect 4356 13574 4402 13626
rect 4106 13572 4162 13574
rect 4186 13572 4242 13574
rect 4266 13572 4322 13574
rect 4346 13572 4402 13574
rect 4106 12538 4162 12540
rect 4186 12538 4242 12540
rect 4266 12538 4322 12540
rect 4346 12538 4402 12540
rect 4106 12486 4152 12538
rect 4152 12486 4162 12538
rect 4186 12486 4216 12538
rect 4216 12486 4228 12538
rect 4228 12486 4242 12538
rect 4266 12486 4280 12538
rect 4280 12486 4292 12538
rect 4292 12486 4322 12538
rect 4346 12486 4356 12538
rect 4356 12486 4402 12538
rect 4106 12484 4162 12486
rect 4186 12484 4242 12486
rect 4266 12484 4322 12486
rect 4346 12484 4402 12486
rect 3514 11212 3570 11248
rect 3514 11192 3516 11212
rect 3516 11192 3568 11212
rect 3568 11192 3570 11212
rect 2255 7642 2311 7644
rect 2335 7642 2391 7644
rect 2415 7642 2471 7644
rect 2495 7642 2551 7644
rect 2255 7590 2301 7642
rect 2301 7590 2311 7642
rect 2335 7590 2365 7642
rect 2365 7590 2377 7642
rect 2377 7590 2391 7642
rect 2415 7590 2429 7642
rect 2429 7590 2441 7642
rect 2441 7590 2471 7642
rect 2495 7590 2505 7642
rect 2505 7590 2551 7642
rect 2255 7588 2311 7590
rect 2335 7588 2391 7590
rect 2415 7588 2471 7590
rect 2495 7588 2551 7590
rect 5957 14170 6013 14172
rect 6037 14170 6093 14172
rect 6117 14170 6173 14172
rect 6197 14170 6253 14172
rect 5957 14118 6003 14170
rect 6003 14118 6013 14170
rect 6037 14118 6067 14170
rect 6067 14118 6079 14170
rect 6079 14118 6093 14170
rect 6117 14118 6131 14170
rect 6131 14118 6143 14170
rect 6143 14118 6173 14170
rect 6197 14118 6207 14170
rect 6207 14118 6253 14170
rect 5957 14116 6013 14118
rect 6037 14116 6093 14118
rect 6117 14116 6173 14118
rect 6197 14116 6253 14118
rect 9659 15258 9715 15260
rect 9739 15258 9795 15260
rect 9819 15258 9875 15260
rect 9899 15258 9955 15260
rect 9659 15206 9705 15258
rect 9705 15206 9715 15258
rect 9739 15206 9769 15258
rect 9769 15206 9781 15258
rect 9781 15206 9795 15258
rect 9819 15206 9833 15258
rect 9833 15206 9845 15258
rect 9845 15206 9875 15258
rect 9899 15206 9909 15258
rect 9909 15206 9955 15258
rect 9659 15204 9715 15206
rect 9739 15204 9795 15206
rect 9819 15204 9875 15206
rect 9899 15204 9955 15206
rect 4106 11450 4162 11452
rect 4186 11450 4242 11452
rect 4266 11450 4322 11452
rect 4346 11450 4402 11452
rect 4106 11398 4152 11450
rect 4152 11398 4162 11450
rect 4186 11398 4216 11450
rect 4216 11398 4228 11450
rect 4228 11398 4242 11450
rect 4266 11398 4280 11450
rect 4280 11398 4292 11450
rect 4292 11398 4322 11450
rect 4346 11398 4356 11450
rect 4356 11398 4402 11450
rect 4106 11396 4162 11398
rect 4186 11396 4242 11398
rect 4266 11396 4322 11398
rect 4346 11396 4402 11398
rect 4066 11212 4122 11248
rect 4066 11192 4068 11212
rect 4068 11192 4120 11212
rect 4120 11192 4122 11212
rect 2255 6554 2311 6556
rect 2335 6554 2391 6556
rect 2415 6554 2471 6556
rect 2495 6554 2551 6556
rect 2255 6502 2301 6554
rect 2301 6502 2311 6554
rect 2335 6502 2365 6554
rect 2365 6502 2377 6554
rect 2377 6502 2391 6554
rect 2415 6502 2429 6554
rect 2429 6502 2441 6554
rect 2441 6502 2471 6554
rect 2495 6502 2505 6554
rect 2505 6502 2551 6554
rect 2255 6500 2311 6502
rect 2335 6500 2391 6502
rect 2415 6500 2471 6502
rect 2495 6500 2551 6502
rect 2255 5466 2311 5468
rect 2335 5466 2391 5468
rect 2415 5466 2471 5468
rect 2495 5466 2551 5468
rect 2255 5414 2301 5466
rect 2301 5414 2311 5466
rect 2335 5414 2365 5466
rect 2365 5414 2377 5466
rect 2377 5414 2391 5466
rect 2415 5414 2429 5466
rect 2429 5414 2441 5466
rect 2441 5414 2471 5466
rect 2495 5414 2505 5466
rect 2505 5414 2551 5466
rect 2255 5412 2311 5414
rect 2335 5412 2391 5414
rect 2415 5412 2471 5414
rect 2495 5412 2551 5414
rect 4618 11192 4674 11248
rect 4526 11092 4528 11112
rect 4528 11092 4580 11112
rect 4580 11092 4582 11112
rect 4526 11056 4582 11092
rect 4106 10362 4162 10364
rect 4186 10362 4242 10364
rect 4266 10362 4322 10364
rect 4346 10362 4402 10364
rect 4106 10310 4152 10362
rect 4152 10310 4162 10362
rect 4186 10310 4216 10362
rect 4216 10310 4228 10362
rect 4228 10310 4242 10362
rect 4266 10310 4280 10362
rect 4280 10310 4292 10362
rect 4292 10310 4322 10362
rect 4346 10310 4356 10362
rect 4356 10310 4402 10362
rect 4106 10308 4162 10310
rect 4186 10308 4242 10310
rect 4266 10308 4322 10310
rect 4346 10308 4402 10310
rect 4106 9274 4162 9276
rect 4186 9274 4242 9276
rect 4266 9274 4322 9276
rect 4346 9274 4402 9276
rect 4106 9222 4152 9274
rect 4152 9222 4162 9274
rect 4186 9222 4216 9274
rect 4216 9222 4228 9274
rect 4228 9222 4242 9274
rect 4266 9222 4280 9274
rect 4280 9222 4292 9274
rect 4292 9222 4322 9274
rect 4346 9222 4356 9274
rect 4356 9222 4402 9274
rect 4106 9220 4162 9222
rect 4186 9220 4242 9222
rect 4266 9220 4322 9222
rect 4346 9220 4402 9222
rect 4986 11092 4988 11112
rect 4988 11092 5040 11112
rect 5040 11092 5042 11112
rect 4986 11056 5042 11092
rect 4106 8186 4162 8188
rect 4186 8186 4242 8188
rect 4266 8186 4322 8188
rect 4346 8186 4402 8188
rect 4106 8134 4152 8186
rect 4152 8134 4162 8186
rect 4186 8134 4216 8186
rect 4216 8134 4228 8186
rect 4228 8134 4242 8186
rect 4266 8134 4280 8186
rect 4280 8134 4292 8186
rect 4292 8134 4322 8186
rect 4346 8134 4356 8186
rect 4356 8134 4402 8186
rect 4106 8132 4162 8134
rect 4186 8132 4242 8134
rect 4266 8132 4322 8134
rect 4346 8132 4402 8134
rect 5957 13082 6013 13084
rect 6037 13082 6093 13084
rect 6117 13082 6173 13084
rect 6197 13082 6253 13084
rect 5957 13030 6003 13082
rect 6003 13030 6013 13082
rect 6037 13030 6067 13082
rect 6067 13030 6079 13082
rect 6079 13030 6093 13082
rect 6117 13030 6131 13082
rect 6131 13030 6143 13082
rect 6143 13030 6173 13082
rect 6197 13030 6207 13082
rect 6207 13030 6253 13082
rect 5957 13028 6013 13030
rect 6037 13028 6093 13030
rect 6117 13028 6173 13030
rect 6197 13028 6253 13030
rect 5262 11192 5318 11248
rect 5957 11994 6013 11996
rect 6037 11994 6093 11996
rect 6117 11994 6173 11996
rect 6197 11994 6253 11996
rect 5957 11942 6003 11994
rect 6003 11942 6013 11994
rect 6037 11942 6067 11994
rect 6067 11942 6079 11994
rect 6079 11942 6093 11994
rect 6117 11942 6131 11994
rect 6131 11942 6143 11994
rect 6143 11942 6173 11994
rect 6197 11942 6207 11994
rect 6207 11942 6253 11994
rect 5957 11940 6013 11942
rect 6037 11940 6093 11942
rect 6117 11940 6173 11942
rect 6197 11940 6253 11942
rect 5957 10906 6013 10908
rect 6037 10906 6093 10908
rect 6117 10906 6173 10908
rect 6197 10906 6253 10908
rect 5957 10854 6003 10906
rect 6003 10854 6013 10906
rect 6037 10854 6067 10906
rect 6067 10854 6079 10906
rect 6079 10854 6093 10906
rect 6117 10854 6131 10906
rect 6131 10854 6143 10906
rect 6143 10854 6173 10906
rect 6197 10854 6207 10906
rect 6207 10854 6253 10906
rect 5957 10852 6013 10854
rect 6037 10852 6093 10854
rect 6117 10852 6173 10854
rect 6197 10852 6253 10854
rect 5957 9818 6013 9820
rect 6037 9818 6093 9820
rect 6117 9818 6173 9820
rect 6197 9818 6253 9820
rect 5957 9766 6003 9818
rect 6003 9766 6013 9818
rect 6037 9766 6067 9818
rect 6067 9766 6079 9818
rect 6079 9766 6093 9818
rect 6117 9766 6131 9818
rect 6131 9766 6143 9818
rect 6143 9766 6173 9818
rect 6197 9766 6207 9818
rect 6207 9766 6253 9818
rect 5957 9764 6013 9766
rect 6037 9764 6093 9766
rect 6117 9764 6173 9766
rect 6197 9764 6253 9766
rect 4106 7098 4162 7100
rect 4186 7098 4242 7100
rect 4266 7098 4322 7100
rect 4346 7098 4402 7100
rect 4106 7046 4152 7098
rect 4152 7046 4162 7098
rect 4186 7046 4216 7098
rect 4216 7046 4228 7098
rect 4228 7046 4242 7098
rect 4266 7046 4280 7098
rect 4280 7046 4292 7098
rect 4292 7046 4322 7098
rect 4346 7046 4356 7098
rect 4356 7046 4402 7098
rect 4106 7044 4162 7046
rect 4186 7044 4242 7046
rect 4266 7044 4322 7046
rect 4346 7044 4402 7046
rect 6366 9016 6422 9072
rect 5957 8730 6013 8732
rect 6037 8730 6093 8732
rect 6117 8730 6173 8732
rect 6197 8730 6253 8732
rect 5957 8678 6003 8730
rect 6003 8678 6013 8730
rect 6037 8678 6067 8730
rect 6067 8678 6079 8730
rect 6079 8678 6093 8730
rect 6117 8678 6131 8730
rect 6131 8678 6143 8730
rect 6143 8678 6173 8730
rect 6197 8678 6207 8730
rect 6207 8678 6253 8730
rect 5957 8676 6013 8678
rect 6037 8676 6093 8678
rect 6117 8676 6173 8678
rect 6197 8676 6253 8678
rect 7808 14714 7864 14716
rect 7888 14714 7944 14716
rect 7968 14714 8024 14716
rect 8048 14714 8104 14716
rect 7808 14662 7854 14714
rect 7854 14662 7864 14714
rect 7888 14662 7918 14714
rect 7918 14662 7930 14714
rect 7930 14662 7944 14714
rect 7968 14662 7982 14714
rect 7982 14662 7994 14714
rect 7994 14662 8024 14714
rect 8048 14662 8058 14714
rect 8058 14662 8104 14714
rect 7808 14660 7864 14662
rect 7888 14660 7944 14662
rect 7968 14660 8024 14662
rect 8048 14660 8104 14662
rect 7808 13626 7864 13628
rect 7888 13626 7944 13628
rect 7968 13626 8024 13628
rect 8048 13626 8104 13628
rect 7808 13574 7854 13626
rect 7854 13574 7864 13626
rect 7888 13574 7918 13626
rect 7918 13574 7930 13626
rect 7930 13574 7944 13626
rect 7968 13574 7982 13626
rect 7982 13574 7994 13626
rect 7994 13574 8024 13626
rect 8048 13574 8058 13626
rect 8058 13574 8104 13626
rect 7808 13572 7864 13574
rect 7888 13572 7944 13574
rect 7968 13572 8024 13574
rect 8048 13572 8104 13574
rect 7808 12538 7864 12540
rect 7888 12538 7944 12540
rect 7968 12538 8024 12540
rect 8048 12538 8104 12540
rect 7808 12486 7854 12538
rect 7854 12486 7864 12538
rect 7888 12486 7918 12538
rect 7918 12486 7930 12538
rect 7930 12486 7944 12538
rect 7968 12486 7982 12538
rect 7982 12486 7994 12538
rect 7994 12486 8024 12538
rect 8048 12486 8058 12538
rect 8058 12486 8104 12538
rect 7808 12484 7864 12486
rect 7888 12484 7944 12486
rect 7968 12484 8024 12486
rect 8048 12484 8104 12486
rect 7808 11450 7864 11452
rect 7888 11450 7944 11452
rect 7968 11450 8024 11452
rect 8048 11450 8104 11452
rect 7808 11398 7854 11450
rect 7854 11398 7864 11450
rect 7888 11398 7918 11450
rect 7918 11398 7930 11450
rect 7930 11398 7944 11450
rect 7968 11398 7982 11450
rect 7982 11398 7994 11450
rect 7994 11398 8024 11450
rect 8048 11398 8058 11450
rect 8058 11398 8104 11450
rect 7808 11396 7864 11398
rect 7888 11396 7944 11398
rect 7968 11396 8024 11398
rect 8048 11396 8104 11398
rect 7808 10362 7864 10364
rect 7888 10362 7944 10364
rect 7968 10362 8024 10364
rect 8048 10362 8104 10364
rect 7808 10310 7854 10362
rect 7854 10310 7864 10362
rect 7888 10310 7918 10362
rect 7918 10310 7930 10362
rect 7930 10310 7944 10362
rect 7968 10310 7982 10362
rect 7982 10310 7994 10362
rect 7994 10310 8024 10362
rect 8048 10310 8058 10362
rect 8058 10310 8104 10362
rect 7808 10308 7864 10310
rect 7888 10308 7944 10310
rect 7968 10308 8024 10310
rect 8048 10308 8104 10310
rect 5957 7642 6013 7644
rect 6037 7642 6093 7644
rect 6117 7642 6173 7644
rect 6197 7642 6253 7644
rect 5957 7590 6003 7642
rect 6003 7590 6013 7642
rect 6037 7590 6067 7642
rect 6067 7590 6079 7642
rect 6079 7590 6093 7642
rect 6117 7590 6131 7642
rect 6131 7590 6143 7642
rect 6143 7590 6173 7642
rect 6197 7590 6207 7642
rect 6207 7590 6253 7642
rect 5957 7588 6013 7590
rect 6037 7588 6093 7590
rect 6117 7588 6173 7590
rect 6197 7588 6253 7590
rect 7808 9274 7864 9276
rect 7888 9274 7944 9276
rect 7968 9274 8024 9276
rect 8048 9274 8104 9276
rect 7808 9222 7854 9274
rect 7854 9222 7864 9274
rect 7888 9222 7918 9274
rect 7918 9222 7930 9274
rect 7930 9222 7944 9274
rect 7968 9222 7982 9274
rect 7982 9222 7994 9274
rect 7994 9222 8024 9274
rect 8048 9222 8058 9274
rect 8058 9222 8104 9274
rect 7808 9220 7864 9222
rect 7888 9220 7944 9222
rect 7968 9220 8024 9222
rect 8048 9220 8104 9222
rect 7808 8186 7864 8188
rect 7888 8186 7944 8188
rect 7968 8186 8024 8188
rect 8048 8186 8104 8188
rect 7808 8134 7854 8186
rect 7854 8134 7864 8186
rect 7888 8134 7918 8186
rect 7918 8134 7930 8186
rect 7930 8134 7944 8186
rect 7968 8134 7982 8186
rect 7982 8134 7994 8186
rect 7994 8134 8024 8186
rect 8048 8134 8058 8186
rect 8058 8134 8104 8186
rect 7808 8132 7864 8134
rect 7888 8132 7944 8134
rect 7968 8132 8024 8134
rect 8048 8132 8104 8134
rect 5957 6554 6013 6556
rect 6037 6554 6093 6556
rect 6117 6554 6173 6556
rect 6197 6554 6253 6556
rect 5957 6502 6003 6554
rect 6003 6502 6013 6554
rect 6037 6502 6067 6554
rect 6067 6502 6079 6554
rect 6079 6502 6093 6554
rect 6117 6502 6131 6554
rect 6131 6502 6143 6554
rect 6143 6502 6173 6554
rect 6197 6502 6207 6554
rect 6207 6502 6253 6554
rect 5957 6500 6013 6502
rect 6037 6500 6093 6502
rect 6117 6500 6173 6502
rect 6197 6500 6253 6502
rect 4106 6010 4162 6012
rect 4186 6010 4242 6012
rect 4266 6010 4322 6012
rect 4346 6010 4402 6012
rect 4106 5958 4152 6010
rect 4152 5958 4162 6010
rect 4186 5958 4216 6010
rect 4216 5958 4228 6010
rect 4228 5958 4242 6010
rect 4266 5958 4280 6010
rect 4280 5958 4292 6010
rect 4292 5958 4322 6010
rect 4346 5958 4356 6010
rect 4356 5958 4402 6010
rect 4106 5956 4162 5958
rect 4186 5956 4242 5958
rect 4266 5956 4322 5958
rect 4346 5956 4402 5958
rect 7838 7248 7894 7304
rect 7808 7098 7864 7100
rect 7888 7098 7944 7100
rect 7968 7098 8024 7100
rect 8048 7098 8104 7100
rect 7808 7046 7854 7098
rect 7854 7046 7864 7098
rect 7888 7046 7918 7098
rect 7918 7046 7930 7098
rect 7930 7046 7944 7098
rect 7968 7046 7982 7098
rect 7982 7046 7994 7098
rect 7994 7046 8024 7098
rect 8048 7046 8058 7098
rect 8058 7046 8104 7098
rect 7808 7044 7864 7046
rect 7888 7044 7944 7046
rect 7968 7044 8024 7046
rect 8048 7044 8104 7046
rect 7808 6010 7864 6012
rect 7888 6010 7944 6012
rect 7968 6010 8024 6012
rect 8048 6010 8104 6012
rect 7808 5958 7854 6010
rect 7854 5958 7864 6010
rect 7888 5958 7918 6010
rect 7918 5958 7930 6010
rect 7930 5958 7944 6010
rect 7968 5958 7982 6010
rect 7982 5958 7994 6010
rect 7994 5958 8024 6010
rect 8048 5958 8058 6010
rect 8058 5958 8104 6010
rect 7808 5956 7864 5958
rect 7888 5956 7944 5958
rect 7968 5956 8024 5958
rect 8048 5956 8104 5958
rect 9659 14170 9715 14172
rect 9739 14170 9795 14172
rect 9819 14170 9875 14172
rect 9899 14170 9955 14172
rect 9659 14118 9705 14170
rect 9705 14118 9715 14170
rect 9739 14118 9769 14170
rect 9769 14118 9781 14170
rect 9781 14118 9795 14170
rect 9819 14118 9833 14170
rect 9833 14118 9845 14170
rect 9845 14118 9875 14170
rect 9899 14118 9909 14170
rect 9909 14118 9955 14170
rect 9659 14116 9715 14118
rect 9739 14116 9795 14118
rect 9819 14116 9875 14118
rect 9899 14116 9955 14118
rect 9659 13082 9715 13084
rect 9739 13082 9795 13084
rect 9819 13082 9875 13084
rect 9899 13082 9955 13084
rect 9659 13030 9705 13082
rect 9705 13030 9715 13082
rect 9739 13030 9769 13082
rect 9769 13030 9781 13082
rect 9781 13030 9795 13082
rect 9819 13030 9833 13082
rect 9833 13030 9845 13082
rect 9845 13030 9875 13082
rect 9899 13030 9909 13082
rect 9909 13030 9955 13082
rect 9659 13028 9715 13030
rect 9739 13028 9795 13030
rect 9819 13028 9875 13030
rect 9899 13028 9955 13030
rect 9659 11994 9715 11996
rect 9739 11994 9795 11996
rect 9819 11994 9875 11996
rect 9899 11994 9955 11996
rect 9659 11942 9705 11994
rect 9705 11942 9715 11994
rect 9739 11942 9769 11994
rect 9769 11942 9781 11994
rect 9781 11942 9795 11994
rect 9819 11942 9833 11994
rect 9833 11942 9845 11994
rect 9845 11942 9875 11994
rect 9899 11942 9909 11994
rect 9909 11942 9955 11994
rect 9659 11940 9715 11942
rect 9739 11940 9795 11942
rect 9819 11940 9875 11942
rect 9899 11940 9955 11942
rect 9310 9016 9366 9072
rect 8850 6296 8906 6352
rect 9659 10906 9715 10908
rect 9739 10906 9795 10908
rect 9819 10906 9875 10908
rect 9899 10906 9955 10908
rect 9659 10854 9705 10906
rect 9705 10854 9715 10906
rect 9739 10854 9769 10906
rect 9769 10854 9781 10906
rect 9781 10854 9795 10906
rect 9819 10854 9833 10906
rect 9833 10854 9845 10906
rect 9845 10854 9875 10906
rect 9899 10854 9909 10906
rect 9909 10854 9955 10906
rect 9659 10852 9715 10854
rect 9739 10852 9795 10854
rect 9819 10852 9875 10854
rect 9899 10852 9955 10854
rect 9659 9818 9715 9820
rect 9739 9818 9795 9820
rect 9819 9818 9875 9820
rect 9899 9818 9955 9820
rect 9659 9766 9705 9818
rect 9705 9766 9715 9818
rect 9739 9766 9769 9818
rect 9769 9766 9781 9818
rect 9781 9766 9795 9818
rect 9819 9766 9833 9818
rect 9833 9766 9845 9818
rect 9845 9766 9875 9818
rect 9899 9766 9909 9818
rect 9909 9766 9955 9818
rect 9659 9764 9715 9766
rect 9739 9764 9795 9766
rect 9819 9764 9875 9766
rect 9899 9764 9955 9766
rect 9586 9016 9642 9072
rect 9659 8730 9715 8732
rect 9739 8730 9795 8732
rect 9819 8730 9875 8732
rect 9899 8730 9955 8732
rect 9659 8678 9705 8730
rect 9705 8678 9715 8730
rect 9739 8678 9769 8730
rect 9769 8678 9781 8730
rect 9781 8678 9795 8730
rect 9819 8678 9833 8730
rect 9833 8678 9845 8730
rect 9845 8678 9875 8730
rect 9899 8678 9909 8730
rect 9909 8678 9955 8730
rect 9659 8676 9715 8678
rect 9739 8676 9795 8678
rect 9819 8676 9875 8678
rect 9899 8676 9955 8678
rect 9659 7642 9715 7644
rect 9739 7642 9795 7644
rect 9819 7642 9875 7644
rect 9899 7642 9955 7644
rect 9659 7590 9705 7642
rect 9705 7590 9715 7642
rect 9739 7590 9769 7642
rect 9769 7590 9781 7642
rect 9781 7590 9795 7642
rect 9819 7590 9833 7642
rect 9833 7590 9845 7642
rect 9845 7590 9875 7642
rect 9899 7590 9909 7642
rect 9909 7590 9955 7642
rect 9659 7588 9715 7590
rect 9739 7588 9795 7590
rect 9819 7588 9875 7590
rect 9899 7588 9955 7590
rect 9659 6554 9715 6556
rect 9739 6554 9795 6556
rect 9819 6554 9875 6556
rect 9899 6554 9955 6556
rect 9659 6502 9705 6554
rect 9705 6502 9715 6554
rect 9739 6502 9769 6554
rect 9769 6502 9781 6554
rect 9781 6502 9795 6554
rect 9819 6502 9833 6554
rect 9833 6502 9845 6554
rect 9845 6502 9875 6554
rect 9899 6502 9909 6554
rect 9909 6502 9955 6554
rect 9659 6500 9715 6502
rect 9739 6500 9795 6502
rect 9819 6500 9875 6502
rect 9899 6500 9955 6502
rect 10046 6296 10102 6352
rect 5957 5466 6013 5468
rect 6037 5466 6093 5468
rect 6117 5466 6173 5468
rect 6197 5466 6253 5468
rect 5957 5414 6003 5466
rect 6003 5414 6013 5466
rect 6037 5414 6067 5466
rect 6067 5414 6079 5466
rect 6079 5414 6093 5466
rect 6117 5414 6131 5466
rect 6131 5414 6143 5466
rect 6143 5414 6173 5466
rect 6197 5414 6207 5466
rect 6207 5414 6253 5466
rect 5957 5412 6013 5414
rect 6037 5412 6093 5414
rect 6117 5412 6173 5414
rect 6197 5412 6253 5414
rect 9659 5466 9715 5468
rect 9739 5466 9795 5468
rect 9819 5466 9875 5468
rect 9899 5466 9955 5468
rect 9659 5414 9705 5466
rect 9705 5414 9715 5466
rect 9739 5414 9769 5466
rect 9769 5414 9781 5466
rect 9781 5414 9795 5466
rect 9819 5414 9833 5466
rect 9833 5414 9845 5466
rect 9845 5414 9875 5466
rect 9899 5414 9909 5466
rect 9909 5414 9955 5466
rect 9659 5412 9715 5414
rect 9739 5412 9795 5414
rect 9819 5412 9875 5414
rect 9899 5412 9955 5414
rect 4106 4922 4162 4924
rect 4186 4922 4242 4924
rect 4266 4922 4322 4924
rect 4346 4922 4402 4924
rect 4106 4870 4152 4922
rect 4152 4870 4162 4922
rect 4186 4870 4216 4922
rect 4216 4870 4228 4922
rect 4228 4870 4242 4922
rect 4266 4870 4280 4922
rect 4280 4870 4292 4922
rect 4292 4870 4322 4922
rect 4346 4870 4356 4922
rect 4356 4870 4402 4922
rect 4106 4868 4162 4870
rect 4186 4868 4242 4870
rect 4266 4868 4322 4870
rect 4346 4868 4402 4870
rect 7808 4922 7864 4924
rect 7888 4922 7944 4924
rect 7968 4922 8024 4924
rect 8048 4922 8104 4924
rect 7808 4870 7854 4922
rect 7854 4870 7864 4922
rect 7888 4870 7918 4922
rect 7918 4870 7930 4922
rect 7930 4870 7944 4922
rect 7968 4870 7982 4922
rect 7982 4870 7994 4922
rect 7994 4870 8024 4922
rect 8048 4870 8058 4922
rect 8058 4870 8104 4922
rect 7808 4868 7864 4870
rect 7888 4868 7944 4870
rect 7968 4868 8024 4870
rect 8048 4868 8104 4870
rect 2255 4378 2311 4380
rect 2335 4378 2391 4380
rect 2415 4378 2471 4380
rect 2495 4378 2551 4380
rect 2255 4326 2301 4378
rect 2301 4326 2311 4378
rect 2335 4326 2365 4378
rect 2365 4326 2377 4378
rect 2377 4326 2391 4378
rect 2415 4326 2429 4378
rect 2429 4326 2441 4378
rect 2441 4326 2471 4378
rect 2495 4326 2505 4378
rect 2505 4326 2551 4378
rect 2255 4324 2311 4326
rect 2335 4324 2391 4326
rect 2415 4324 2471 4326
rect 2495 4324 2551 4326
rect 5957 4378 6013 4380
rect 6037 4378 6093 4380
rect 6117 4378 6173 4380
rect 6197 4378 6253 4380
rect 5957 4326 6003 4378
rect 6003 4326 6013 4378
rect 6037 4326 6067 4378
rect 6067 4326 6079 4378
rect 6079 4326 6093 4378
rect 6117 4326 6131 4378
rect 6131 4326 6143 4378
rect 6143 4326 6173 4378
rect 6197 4326 6207 4378
rect 6207 4326 6253 4378
rect 5957 4324 6013 4326
rect 6037 4324 6093 4326
rect 6117 4324 6173 4326
rect 6197 4324 6253 4326
rect 9659 4378 9715 4380
rect 9739 4378 9795 4380
rect 9819 4378 9875 4380
rect 9899 4378 9955 4380
rect 9659 4326 9705 4378
rect 9705 4326 9715 4378
rect 9739 4326 9769 4378
rect 9769 4326 9781 4378
rect 9781 4326 9795 4378
rect 9819 4326 9833 4378
rect 9833 4326 9845 4378
rect 9845 4326 9875 4378
rect 9899 4326 9909 4378
rect 9909 4326 9955 4378
rect 9659 4324 9715 4326
rect 9739 4324 9795 4326
rect 9819 4324 9875 4326
rect 9899 4324 9955 4326
rect 11510 14714 11566 14716
rect 11590 14714 11646 14716
rect 11670 14714 11726 14716
rect 11750 14714 11806 14716
rect 11510 14662 11556 14714
rect 11556 14662 11566 14714
rect 11590 14662 11620 14714
rect 11620 14662 11632 14714
rect 11632 14662 11646 14714
rect 11670 14662 11684 14714
rect 11684 14662 11696 14714
rect 11696 14662 11726 14714
rect 11750 14662 11760 14714
rect 11760 14662 11806 14714
rect 11510 14660 11566 14662
rect 11590 14660 11646 14662
rect 11670 14660 11726 14662
rect 11750 14660 11806 14662
rect 11510 13626 11566 13628
rect 11590 13626 11646 13628
rect 11670 13626 11726 13628
rect 11750 13626 11806 13628
rect 11510 13574 11556 13626
rect 11556 13574 11566 13626
rect 11590 13574 11620 13626
rect 11620 13574 11632 13626
rect 11632 13574 11646 13626
rect 11670 13574 11684 13626
rect 11684 13574 11696 13626
rect 11696 13574 11726 13626
rect 11750 13574 11760 13626
rect 11760 13574 11806 13626
rect 11510 13572 11566 13574
rect 11590 13572 11646 13574
rect 11670 13572 11726 13574
rect 11750 13572 11806 13574
rect 13361 15258 13417 15260
rect 13441 15258 13497 15260
rect 13521 15258 13577 15260
rect 13601 15258 13657 15260
rect 13361 15206 13407 15258
rect 13407 15206 13417 15258
rect 13441 15206 13471 15258
rect 13471 15206 13483 15258
rect 13483 15206 13497 15258
rect 13521 15206 13535 15258
rect 13535 15206 13547 15258
rect 13547 15206 13577 15258
rect 13601 15206 13611 15258
rect 13611 15206 13657 15258
rect 13361 15204 13417 15206
rect 13441 15204 13497 15206
rect 13521 15204 13577 15206
rect 13601 15204 13657 15206
rect 11510 12538 11566 12540
rect 11590 12538 11646 12540
rect 11670 12538 11726 12540
rect 11750 12538 11806 12540
rect 11510 12486 11556 12538
rect 11556 12486 11566 12538
rect 11590 12486 11620 12538
rect 11620 12486 11632 12538
rect 11632 12486 11646 12538
rect 11670 12486 11684 12538
rect 11684 12486 11696 12538
rect 11696 12486 11726 12538
rect 11750 12486 11760 12538
rect 11760 12486 11806 12538
rect 11510 12484 11566 12486
rect 11590 12484 11646 12486
rect 11670 12484 11726 12486
rect 11750 12484 11806 12486
rect 11510 11450 11566 11452
rect 11590 11450 11646 11452
rect 11670 11450 11726 11452
rect 11750 11450 11806 11452
rect 11510 11398 11556 11450
rect 11556 11398 11566 11450
rect 11590 11398 11620 11450
rect 11620 11398 11632 11450
rect 11632 11398 11646 11450
rect 11670 11398 11684 11450
rect 11684 11398 11696 11450
rect 11696 11398 11726 11450
rect 11750 11398 11760 11450
rect 11760 11398 11806 11450
rect 11510 11396 11566 11398
rect 11590 11396 11646 11398
rect 11670 11396 11726 11398
rect 11750 11396 11806 11398
rect 11510 10362 11566 10364
rect 11590 10362 11646 10364
rect 11670 10362 11726 10364
rect 11750 10362 11806 10364
rect 11510 10310 11556 10362
rect 11556 10310 11566 10362
rect 11590 10310 11620 10362
rect 11620 10310 11632 10362
rect 11632 10310 11646 10362
rect 11670 10310 11684 10362
rect 11684 10310 11696 10362
rect 11696 10310 11726 10362
rect 11750 10310 11760 10362
rect 11760 10310 11806 10362
rect 11510 10308 11566 10310
rect 11590 10308 11646 10310
rect 11670 10308 11726 10310
rect 11750 10308 11806 10310
rect 11510 9274 11566 9276
rect 11590 9274 11646 9276
rect 11670 9274 11726 9276
rect 11750 9274 11806 9276
rect 11510 9222 11556 9274
rect 11556 9222 11566 9274
rect 11590 9222 11620 9274
rect 11620 9222 11632 9274
rect 11632 9222 11646 9274
rect 11670 9222 11684 9274
rect 11684 9222 11696 9274
rect 11696 9222 11726 9274
rect 11750 9222 11760 9274
rect 11760 9222 11806 9274
rect 11510 9220 11566 9222
rect 11590 9220 11646 9222
rect 11670 9220 11726 9222
rect 11750 9220 11806 9222
rect 11510 8186 11566 8188
rect 11590 8186 11646 8188
rect 11670 8186 11726 8188
rect 11750 8186 11806 8188
rect 11510 8134 11556 8186
rect 11556 8134 11566 8186
rect 11590 8134 11620 8186
rect 11620 8134 11632 8186
rect 11632 8134 11646 8186
rect 11670 8134 11684 8186
rect 11684 8134 11696 8186
rect 11696 8134 11726 8186
rect 11750 8134 11760 8186
rect 11760 8134 11806 8186
rect 11510 8132 11566 8134
rect 11590 8132 11646 8134
rect 11670 8132 11726 8134
rect 11750 8132 11806 8134
rect 13361 14170 13417 14172
rect 13441 14170 13497 14172
rect 13521 14170 13577 14172
rect 13601 14170 13657 14172
rect 13361 14118 13407 14170
rect 13407 14118 13417 14170
rect 13441 14118 13471 14170
rect 13471 14118 13483 14170
rect 13483 14118 13497 14170
rect 13521 14118 13535 14170
rect 13535 14118 13547 14170
rect 13547 14118 13577 14170
rect 13601 14118 13611 14170
rect 13611 14118 13657 14170
rect 13361 14116 13417 14118
rect 13441 14116 13497 14118
rect 13521 14116 13577 14118
rect 13601 14116 13657 14118
rect 12990 12724 12992 12744
rect 12992 12724 13044 12744
rect 13044 12724 13046 12744
rect 12990 12688 13046 12724
rect 15212 14714 15268 14716
rect 15292 14714 15348 14716
rect 15372 14714 15428 14716
rect 15452 14714 15508 14716
rect 15212 14662 15258 14714
rect 15258 14662 15268 14714
rect 15292 14662 15322 14714
rect 15322 14662 15334 14714
rect 15334 14662 15348 14714
rect 15372 14662 15386 14714
rect 15386 14662 15398 14714
rect 15398 14662 15428 14714
rect 15452 14662 15462 14714
rect 15462 14662 15508 14714
rect 15212 14660 15268 14662
rect 15292 14660 15348 14662
rect 15372 14660 15428 14662
rect 15452 14660 15508 14662
rect 15014 14476 15070 14512
rect 15014 14456 15016 14476
rect 15016 14456 15068 14476
rect 15068 14456 15070 14476
rect 15212 13626 15268 13628
rect 15292 13626 15348 13628
rect 15372 13626 15428 13628
rect 15452 13626 15508 13628
rect 15212 13574 15258 13626
rect 15258 13574 15268 13626
rect 15292 13574 15322 13626
rect 15322 13574 15334 13626
rect 15334 13574 15348 13626
rect 15372 13574 15386 13626
rect 15386 13574 15398 13626
rect 15398 13574 15428 13626
rect 15452 13574 15462 13626
rect 15462 13574 15508 13626
rect 15212 13572 15268 13574
rect 15292 13572 15348 13574
rect 15372 13572 15428 13574
rect 15452 13572 15508 13574
rect 13361 13082 13417 13084
rect 13441 13082 13497 13084
rect 13521 13082 13577 13084
rect 13601 13082 13657 13084
rect 13361 13030 13407 13082
rect 13407 13030 13417 13082
rect 13441 13030 13471 13082
rect 13471 13030 13483 13082
rect 13483 13030 13497 13082
rect 13521 13030 13535 13082
rect 13535 13030 13547 13082
rect 13547 13030 13577 13082
rect 13601 13030 13611 13082
rect 13611 13030 13657 13082
rect 13361 13028 13417 13030
rect 13441 13028 13497 13030
rect 13521 13028 13577 13030
rect 13601 13028 13657 13030
rect 13450 12552 13506 12608
rect 12346 10648 12402 10704
rect 12438 9036 12494 9072
rect 13361 11994 13417 11996
rect 13441 11994 13497 11996
rect 13521 11994 13577 11996
rect 13601 11994 13657 11996
rect 13361 11942 13407 11994
rect 13407 11942 13417 11994
rect 13441 11942 13471 11994
rect 13471 11942 13483 11994
rect 13483 11942 13497 11994
rect 13521 11942 13535 11994
rect 13535 11942 13547 11994
rect 13547 11942 13577 11994
rect 13601 11942 13611 11994
rect 13611 11942 13657 11994
rect 13361 11940 13417 11942
rect 13441 11940 13497 11942
rect 13521 11940 13577 11942
rect 13601 11940 13657 11942
rect 14462 12724 14464 12744
rect 14464 12724 14516 12744
rect 14516 12724 14518 12744
rect 14002 12588 14004 12608
rect 14004 12588 14056 12608
rect 14056 12588 14058 12608
rect 14002 12552 14058 12588
rect 14462 12688 14518 12724
rect 12438 9016 12440 9036
rect 12440 9016 12492 9036
rect 12492 9016 12494 9036
rect 11510 7098 11566 7100
rect 11590 7098 11646 7100
rect 11670 7098 11726 7100
rect 11750 7098 11806 7100
rect 11510 7046 11556 7098
rect 11556 7046 11566 7098
rect 11590 7046 11620 7098
rect 11620 7046 11632 7098
rect 11632 7046 11646 7098
rect 11670 7046 11684 7098
rect 11684 7046 11696 7098
rect 11696 7046 11726 7098
rect 11750 7046 11760 7098
rect 11760 7046 11806 7098
rect 11510 7044 11566 7046
rect 11590 7044 11646 7046
rect 11670 7044 11726 7046
rect 11750 7044 11806 7046
rect 12162 7248 12218 7304
rect 11510 6010 11566 6012
rect 11590 6010 11646 6012
rect 11670 6010 11726 6012
rect 11750 6010 11806 6012
rect 11510 5958 11556 6010
rect 11556 5958 11566 6010
rect 11590 5958 11620 6010
rect 11620 5958 11632 6010
rect 11632 5958 11646 6010
rect 11670 5958 11684 6010
rect 11684 5958 11696 6010
rect 11696 5958 11726 6010
rect 11750 5958 11760 6010
rect 11760 5958 11806 6010
rect 11510 5956 11566 5958
rect 11590 5956 11646 5958
rect 11670 5956 11726 5958
rect 11750 5956 11806 5958
rect 13361 10906 13417 10908
rect 13441 10906 13497 10908
rect 13521 10906 13577 10908
rect 13601 10906 13657 10908
rect 13361 10854 13407 10906
rect 13407 10854 13417 10906
rect 13441 10854 13471 10906
rect 13471 10854 13483 10906
rect 13483 10854 13497 10906
rect 13521 10854 13535 10906
rect 13535 10854 13547 10906
rect 13547 10854 13577 10906
rect 13601 10854 13611 10906
rect 13611 10854 13657 10906
rect 13361 10852 13417 10854
rect 13441 10852 13497 10854
rect 13521 10852 13577 10854
rect 13601 10852 13657 10854
rect 15212 12538 15268 12540
rect 15292 12538 15348 12540
rect 15372 12538 15428 12540
rect 15452 12538 15508 12540
rect 15212 12486 15258 12538
rect 15258 12486 15268 12538
rect 15292 12486 15322 12538
rect 15322 12486 15334 12538
rect 15334 12486 15348 12538
rect 15372 12486 15386 12538
rect 15386 12486 15398 12538
rect 15398 12486 15428 12538
rect 15452 12486 15462 12538
rect 15462 12486 15508 12538
rect 15212 12484 15268 12486
rect 15292 12484 15348 12486
rect 15372 12484 15428 12486
rect 15452 12484 15508 12486
rect 15014 12316 15016 12336
rect 15016 12316 15068 12336
rect 15068 12316 15070 12336
rect 15014 12280 15070 12316
rect 15212 11450 15268 11452
rect 15292 11450 15348 11452
rect 15372 11450 15428 11452
rect 15452 11450 15508 11452
rect 15212 11398 15258 11450
rect 15258 11398 15268 11450
rect 15292 11398 15322 11450
rect 15322 11398 15334 11450
rect 15334 11398 15348 11450
rect 15372 11398 15386 11450
rect 15386 11398 15398 11450
rect 15398 11398 15428 11450
rect 15452 11398 15462 11450
rect 15462 11398 15508 11450
rect 15212 11396 15268 11398
rect 15292 11396 15348 11398
rect 15372 11396 15428 11398
rect 15452 11396 15508 11398
rect 13361 9818 13417 9820
rect 13441 9818 13497 9820
rect 13521 9818 13577 9820
rect 13601 9818 13657 9820
rect 13361 9766 13407 9818
rect 13407 9766 13417 9818
rect 13441 9766 13471 9818
rect 13471 9766 13483 9818
rect 13483 9766 13497 9818
rect 13521 9766 13535 9818
rect 13535 9766 13547 9818
rect 13547 9766 13577 9818
rect 13601 9766 13611 9818
rect 13611 9766 13657 9818
rect 13361 9764 13417 9766
rect 13441 9764 13497 9766
rect 13521 9764 13577 9766
rect 13601 9764 13657 9766
rect 13361 8730 13417 8732
rect 13441 8730 13497 8732
rect 13521 8730 13577 8732
rect 13601 8730 13657 8732
rect 13361 8678 13407 8730
rect 13407 8678 13417 8730
rect 13441 8678 13471 8730
rect 13471 8678 13483 8730
rect 13483 8678 13497 8730
rect 13521 8678 13535 8730
rect 13535 8678 13547 8730
rect 13547 8678 13577 8730
rect 13601 8678 13611 8730
rect 13611 8678 13657 8730
rect 13361 8676 13417 8678
rect 13441 8676 13497 8678
rect 13521 8676 13577 8678
rect 13601 8676 13657 8678
rect 14186 10648 14242 10704
rect 14922 10648 14978 10704
rect 15212 10362 15268 10364
rect 15292 10362 15348 10364
rect 15372 10362 15428 10364
rect 15452 10362 15508 10364
rect 15212 10310 15258 10362
rect 15258 10310 15268 10362
rect 15292 10310 15322 10362
rect 15322 10310 15334 10362
rect 15334 10310 15348 10362
rect 15372 10310 15386 10362
rect 15386 10310 15398 10362
rect 15398 10310 15428 10362
rect 15452 10310 15462 10362
rect 15462 10310 15508 10362
rect 15212 10308 15268 10310
rect 15292 10308 15348 10310
rect 15372 10308 15428 10310
rect 15452 10308 15508 10310
rect 13361 7642 13417 7644
rect 13441 7642 13497 7644
rect 13521 7642 13577 7644
rect 13601 7642 13657 7644
rect 13361 7590 13407 7642
rect 13407 7590 13417 7642
rect 13441 7590 13471 7642
rect 13471 7590 13483 7642
rect 13483 7590 13497 7642
rect 13521 7590 13535 7642
rect 13535 7590 13547 7642
rect 13547 7590 13577 7642
rect 13601 7590 13611 7642
rect 13611 7590 13657 7642
rect 13361 7588 13417 7590
rect 13441 7588 13497 7590
rect 13521 7588 13577 7590
rect 13601 7588 13657 7590
rect 15212 9274 15268 9276
rect 15292 9274 15348 9276
rect 15372 9274 15428 9276
rect 15452 9274 15508 9276
rect 15212 9222 15258 9274
rect 15258 9222 15268 9274
rect 15292 9222 15322 9274
rect 15322 9222 15334 9274
rect 15334 9222 15348 9274
rect 15372 9222 15386 9274
rect 15386 9222 15398 9274
rect 15398 9222 15428 9274
rect 15452 9222 15462 9274
rect 15462 9222 15508 9274
rect 15212 9220 15268 9222
rect 15292 9220 15348 9222
rect 15372 9220 15428 9222
rect 15452 9220 15508 9222
rect 15014 8780 15016 8800
rect 15016 8780 15068 8800
rect 15068 8780 15070 8800
rect 15014 8744 15070 8780
rect 13266 7248 13322 7304
rect 11510 4922 11566 4924
rect 11590 4922 11646 4924
rect 11670 4922 11726 4924
rect 11750 4922 11806 4924
rect 11510 4870 11556 4922
rect 11556 4870 11566 4922
rect 11590 4870 11620 4922
rect 11620 4870 11632 4922
rect 11632 4870 11646 4922
rect 11670 4870 11684 4922
rect 11684 4870 11696 4922
rect 11696 4870 11726 4922
rect 11750 4870 11760 4922
rect 11760 4870 11806 4922
rect 11510 4868 11566 4870
rect 11590 4868 11646 4870
rect 11670 4868 11726 4870
rect 11750 4868 11806 4870
rect 13361 6554 13417 6556
rect 13441 6554 13497 6556
rect 13521 6554 13577 6556
rect 13601 6554 13657 6556
rect 13361 6502 13407 6554
rect 13407 6502 13417 6554
rect 13441 6502 13471 6554
rect 13471 6502 13483 6554
rect 13483 6502 13497 6554
rect 13521 6502 13535 6554
rect 13535 6502 13547 6554
rect 13547 6502 13577 6554
rect 13601 6502 13611 6554
rect 13611 6502 13657 6554
rect 13361 6500 13417 6502
rect 13441 6500 13497 6502
rect 13521 6500 13577 6502
rect 13601 6500 13657 6502
rect 15212 8186 15268 8188
rect 15292 8186 15348 8188
rect 15372 8186 15428 8188
rect 15452 8186 15508 8188
rect 15212 8134 15258 8186
rect 15258 8134 15268 8186
rect 15292 8134 15322 8186
rect 15322 8134 15334 8186
rect 15334 8134 15348 8186
rect 15372 8134 15386 8186
rect 15386 8134 15398 8186
rect 15398 8134 15428 8186
rect 15452 8134 15462 8186
rect 15462 8134 15508 8186
rect 15212 8132 15268 8134
rect 15292 8132 15348 8134
rect 15372 8132 15428 8134
rect 15452 8132 15508 8134
rect 15212 7098 15268 7100
rect 15292 7098 15348 7100
rect 15372 7098 15428 7100
rect 15452 7098 15508 7100
rect 15212 7046 15258 7098
rect 15258 7046 15268 7098
rect 15292 7046 15322 7098
rect 15322 7046 15334 7098
rect 15334 7046 15348 7098
rect 15372 7046 15386 7098
rect 15386 7046 15398 7098
rect 15398 7046 15428 7098
rect 15452 7046 15462 7098
rect 15462 7046 15508 7098
rect 15212 7044 15268 7046
rect 15292 7044 15348 7046
rect 15372 7044 15428 7046
rect 15452 7044 15508 7046
rect 15014 6860 15070 6896
rect 15014 6840 15016 6860
rect 15016 6840 15068 6860
rect 15068 6840 15070 6860
rect 14462 5516 14464 5536
rect 14464 5516 14516 5536
rect 14516 5516 14518 5536
rect 14462 5480 14518 5516
rect 13361 5466 13417 5468
rect 13441 5466 13497 5468
rect 13521 5466 13577 5468
rect 13601 5466 13657 5468
rect 13361 5414 13407 5466
rect 13407 5414 13417 5466
rect 13441 5414 13471 5466
rect 13471 5414 13483 5466
rect 13483 5414 13497 5466
rect 13521 5414 13535 5466
rect 13535 5414 13547 5466
rect 13547 5414 13577 5466
rect 13601 5414 13611 5466
rect 13611 5414 13657 5466
rect 13361 5412 13417 5414
rect 13441 5412 13497 5414
rect 13521 5412 13577 5414
rect 13601 5412 13657 5414
rect 15212 6010 15268 6012
rect 15292 6010 15348 6012
rect 15372 6010 15428 6012
rect 15452 6010 15508 6012
rect 15212 5958 15258 6010
rect 15258 5958 15268 6010
rect 15292 5958 15322 6010
rect 15322 5958 15334 6010
rect 15334 5958 15348 6010
rect 15372 5958 15386 6010
rect 15386 5958 15398 6010
rect 15398 5958 15428 6010
rect 15452 5958 15462 6010
rect 15462 5958 15508 6010
rect 15212 5956 15268 5958
rect 15292 5956 15348 5958
rect 15372 5956 15428 5958
rect 15452 5956 15508 5958
rect 13361 4378 13417 4380
rect 13441 4378 13497 4380
rect 13521 4378 13577 4380
rect 13601 4378 13657 4380
rect 13361 4326 13407 4378
rect 13407 4326 13417 4378
rect 13441 4326 13471 4378
rect 13471 4326 13483 4378
rect 13483 4326 13497 4378
rect 13521 4326 13535 4378
rect 13535 4326 13547 4378
rect 13547 4326 13577 4378
rect 13601 4326 13611 4378
rect 13611 4326 13657 4378
rect 13361 4324 13417 4326
rect 13441 4324 13497 4326
rect 13521 4324 13577 4326
rect 13601 4324 13657 4326
rect 4106 3834 4162 3836
rect 4186 3834 4242 3836
rect 4266 3834 4322 3836
rect 4346 3834 4402 3836
rect 4106 3782 4152 3834
rect 4152 3782 4162 3834
rect 4186 3782 4216 3834
rect 4216 3782 4228 3834
rect 4228 3782 4242 3834
rect 4266 3782 4280 3834
rect 4280 3782 4292 3834
rect 4292 3782 4322 3834
rect 4346 3782 4356 3834
rect 4356 3782 4402 3834
rect 4106 3780 4162 3782
rect 4186 3780 4242 3782
rect 4266 3780 4322 3782
rect 4346 3780 4402 3782
rect 7808 3834 7864 3836
rect 7888 3834 7944 3836
rect 7968 3834 8024 3836
rect 8048 3834 8104 3836
rect 7808 3782 7854 3834
rect 7854 3782 7864 3834
rect 7888 3782 7918 3834
rect 7918 3782 7930 3834
rect 7930 3782 7944 3834
rect 7968 3782 7982 3834
rect 7982 3782 7994 3834
rect 7994 3782 8024 3834
rect 8048 3782 8058 3834
rect 8058 3782 8104 3834
rect 7808 3780 7864 3782
rect 7888 3780 7944 3782
rect 7968 3780 8024 3782
rect 8048 3780 8104 3782
rect 11510 3834 11566 3836
rect 11590 3834 11646 3836
rect 11670 3834 11726 3836
rect 11750 3834 11806 3836
rect 11510 3782 11556 3834
rect 11556 3782 11566 3834
rect 11590 3782 11620 3834
rect 11620 3782 11632 3834
rect 11632 3782 11646 3834
rect 11670 3782 11684 3834
rect 11684 3782 11696 3834
rect 11696 3782 11726 3834
rect 11750 3782 11760 3834
rect 11760 3782 11806 3834
rect 11510 3780 11566 3782
rect 11590 3780 11646 3782
rect 11670 3780 11726 3782
rect 11750 3780 11806 3782
rect 2255 3290 2311 3292
rect 2335 3290 2391 3292
rect 2415 3290 2471 3292
rect 2495 3290 2551 3292
rect 2255 3238 2301 3290
rect 2301 3238 2311 3290
rect 2335 3238 2365 3290
rect 2365 3238 2377 3290
rect 2377 3238 2391 3290
rect 2415 3238 2429 3290
rect 2429 3238 2441 3290
rect 2441 3238 2471 3290
rect 2495 3238 2505 3290
rect 2505 3238 2551 3290
rect 2255 3236 2311 3238
rect 2335 3236 2391 3238
rect 2415 3236 2471 3238
rect 2495 3236 2551 3238
rect 5957 3290 6013 3292
rect 6037 3290 6093 3292
rect 6117 3290 6173 3292
rect 6197 3290 6253 3292
rect 5957 3238 6003 3290
rect 6003 3238 6013 3290
rect 6037 3238 6067 3290
rect 6067 3238 6079 3290
rect 6079 3238 6093 3290
rect 6117 3238 6131 3290
rect 6131 3238 6143 3290
rect 6143 3238 6173 3290
rect 6197 3238 6207 3290
rect 6207 3238 6253 3290
rect 5957 3236 6013 3238
rect 6037 3236 6093 3238
rect 6117 3236 6173 3238
rect 6197 3236 6253 3238
rect 9659 3290 9715 3292
rect 9739 3290 9795 3292
rect 9819 3290 9875 3292
rect 9899 3290 9955 3292
rect 9659 3238 9705 3290
rect 9705 3238 9715 3290
rect 9739 3238 9769 3290
rect 9769 3238 9781 3290
rect 9781 3238 9795 3290
rect 9819 3238 9833 3290
rect 9833 3238 9845 3290
rect 9845 3238 9875 3290
rect 9899 3238 9909 3290
rect 9909 3238 9955 3290
rect 9659 3236 9715 3238
rect 9739 3236 9795 3238
rect 9819 3236 9875 3238
rect 9899 3236 9955 3238
rect 4106 2746 4162 2748
rect 4186 2746 4242 2748
rect 4266 2746 4322 2748
rect 4346 2746 4402 2748
rect 4106 2694 4152 2746
rect 4152 2694 4162 2746
rect 4186 2694 4216 2746
rect 4216 2694 4228 2746
rect 4228 2694 4242 2746
rect 4266 2694 4280 2746
rect 4280 2694 4292 2746
rect 4292 2694 4322 2746
rect 4346 2694 4356 2746
rect 4356 2694 4402 2746
rect 4106 2692 4162 2694
rect 4186 2692 4242 2694
rect 4266 2692 4322 2694
rect 4346 2692 4402 2694
rect 7808 2746 7864 2748
rect 7888 2746 7944 2748
rect 7968 2746 8024 2748
rect 8048 2746 8104 2748
rect 7808 2694 7854 2746
rect 7854 2694 7864 2746
rect 7888 2694 7918 2746
rect 7918 2694 7930 2746
rect 7930 2694 7944 2746
rect 7968 2694 7982 2746
rect 7982 2694 7994 2746
rect 7994 2694 8024 2746
rect 8048 2694 8058 2746
rect 8058 2694 8104 2746
rect 7808 2692 7864 2694
rect 7888 2692 7944 2694
rect 7968 2692 8024 2694
rect 8048 2692 8104 2694
rect 11510 2746 11566 2748
rect 11590 2746 11646 2748
rect 11670 2746 11726 2748
rect 11750 2746 11806 2748
rect 11510 2694 11556 2746
rect 11556 2694 11566 2746
rect 11590 2694 11620 2746
rect 11620 2694 11632 2746
rect 11632 2694 11646 2746
rect 11670 2694 11684 2746
rect 11684 2694 11696 2746
rect 11696 2694 11726 2746
rect 11750 2694 11760 2746
rect 11760 2694 11806 2746
rect 11510 2692 11566 2694
rect 11590 2692 11646 2694
rect 11670 2692 11726 2694
rect 11750 2692 11806 2694
rect 2255 2202 2311 2204
rect 2335 2202 2391 2204
rect 2415 2202 2471 2204
rect 2495 2202 2551 2204
rect 2255 2150 2301 2202
rect 2301 2150 2311 2202
rect 2335 2150 2365 2202
rect 2365 2150 2377 2202
rect 2377 2150 2391 2202
rect 2415 2150 2429 2202
rect 2429 2150 2441 2202
rect 2441 2150 2471 2202
rect 2495 2150 2505 2202
rect 2505 2150 2551 2202
rect 2255 2148 2311 2150
rect 2335 2148 2391 2150
rect 2415 2148 2471 2150
rect 2495 2148 2551 2150
rect 5957 2202 6013 2204
rect 6037 2202 6093 2204
rect 6117 2202 6173 2204
rect 6197 2202 6253 2204
rect 5957 2150 6003 2202
rect 6003 2150 6013 2202
rect 6037 2150 6067 2202
rect 6067 2150 6079 2202
rect 6079 2150 6093 2202
rect 6117 2150 6131 2202
rect 6131 2150 6143 2202
rect 6143 2150 6173 2202
rect 6197 2150 6207 2202
rect 6207 2150 6253 2202
rect 5957 2148 6013 2150
rect 6037 2148 6093 2150
rect 6117 2148 6173 2150
rect 6197 2148 6253 2150
rect 9659 2202 9715 2204
rect 9739 2202 9795 2204
rect 9819 2202 9875 2204
rect 9899 2202 9955 2204
rect 9659 2150 9705 2202
rect 9705 2150 9715 2202
rect 9739 2150 9769 2202
rect 9769 2150 9781 2202
rect 9781 2150 9795 2202
rect 9819 2150 9833 2202
rect 9833 2150 9845 2202
rect 9845 2150 9875 2202
rect 9899 2150 9909 2202
rect 9909 2150 9955 2202
rect 9659 2148 9715 2150
rect 9739 2148 9795 2150
rect 9819 2148 9875 2150
rect 9899 2148 9955 2150
rect 4106 1658 4162 1660
rect 4186 1658 4242 1660
rect 4266 1658 4322 1660
rect 4346 1658 4402 1660
rect 4106 1606 4152 1658
rect 4152 1606 4162 1658
rect 4186 1606 4216 1658
rect 4216 1606 4228 1658
rect 4228 1606 4242 1658
rect 4266 1606 4280 1658
rect 4280 1606 4292 1658
rect 4292 1606 4322 1658
rect 4346 1606 4356 1658
rect 4356 1606 4402 1658
rect 4106 1604 4162 1606
rect 4186 1604 4242 1606
rect 4266 1604 4322 1606
rect 4346 1604 4402 1606
rect 7808 1658 7864 1660
rect 7888 1658 7944 1660
rect 7968 1658 8024 1660
rect 8048 1658 8104 1660
rect 7808 1606 7854 1658
rect 7854 1606 7864 1658
rect 7888 1606 7918 1658
rect 7918 1606 7930 1658
rect 7930 1606 7944 1658
rect 7968 1606 7982 1658
rect 7982 1606 7994 1658
rect 7994 1606 8024 1658
rect 8048 1606 8058 1658
rect 8058 1606 8104 1658
rect 7808 1604 7864 1606
rect 7888 1604 7944 1606
rect 7968 1604 8024 1606
rect 8048 1604 8104 1606
rect 11510 1658 11566 1660
rect 11590 1658 11646 1660
rect 11670 1658 11726 1660
rect 11750 1658 11806 1660
rect 11510 1606 11556 1658
rect 11556 1606 11566 1658
rect 11590 1606 11620 1658
rect 11620 1606 11632 1658
rect 11632 1606 11646 1658
rect 11670 1606 11684 1658
rect 11684 1606 11696 1658
rect 11696 1606 11726 1658
rect 11750 1606 11760 1658
rect 11760 1606 11806 1658
rect 11510 1604 11566 1606
rect 11590 1604 11646 1606
rect 11670 1604 11726 1606
rect 11750 1604 11806 1606
rect 13361 3290 13417 3292
rect 13441 3290 13497 3292
rect 13521 3290 13577 3292
rect 13601 3290 13657 3292
rect 13361 3238 13407 3290
rect 13407 3238 13417 3290
rect 13441 3238 13471 3290
rect 13471 3238 13483 3290
rect 13483 3238 13497 3290
rect 13521 3238 13535 3290
rect 13535 3238 13547 3290
rect 13547 3238 13577 3290
rect 13601 3238 13611 3290
rect 13611 3238 13657 3290
rect 13361 3236 13417 3238
rect 13441 3236 13497 3238
rect 13521 3236 13577 3238
rect 13601 3236 13657 3238
rect 15212 4922 15268 4924
rect 15292 4922 15348 4924
rect 15372 4922 15428 4924
rect 15452 4922 15508 4924
rect 15212 4870 15258 4922
rect 15258 4870 15268 4922
rect 15292 4870 15322 4922
rect 15322 4870 15334 4922
rect 15334 4870 15348 4922
rect 15372 4870 15386 4922
rect 15386 4870 15398 4922
rect 15398 4870 15428 4922
rect 15452 4870 15462 4922
rect 15462 4870 15508 4922
rect 15212 4868 15268 4870
rect 15292 4868 15348 4870
rect 15372 4868 15428 4870
rect 15452 4868 15508 4870
rect 15212 3834 15268 3836
rect 15292 3834 15348 3836
rect 15372 3834 15428 3836
rect 15452 3834 15508 3836
rect 15212 3782 15258 3834
rect 15258 3782 15268 3834
rect 15292 3782 15322 3834
rect 15322 3782 15334 3834
rect 15334 3782 15348 3834
rect 15372 3782 15386 3834
rect 15386 3782 15398 3834
rect 15398 3782 15428 3834
rect 15452 3782 15462 3834
rect 15462 3782 15508 3834
rect 15212 3780 15268 3782
rect 15292 3780 15348 3782
rect 15372 3780 15428 3782
rect 15452 3780 15508 3782
rect 14554 3032 14610 3088
rect 15212 2746 15268 2748
rect 15292 2746 15348 2748
rect 15372 2746 15428 2748
rect 15452 2746 15508 2748
rect 15212 2694 15258 2746
rect 15258 2694 15268 2746
rect 15292 2694 15322 2746
rect 15322 2694 15334 2746
rect 15334 2694 15348 2746
rect 15372 2694 15386 2746
rect 15386 2694 15398 2746
rect 15398 2694 15428 2746
rect 15452 2694 15462 2746
rect 15462 2694 15508 2746
rect 15212 2692 15268 2694
rect 15292 2692 15348 2694
rect 15372 2692 15428 2694
rect 15452 2692 15508 2694
rect 13361 2202 13417 2204
rect 13441 2202 13497 2204
rect 13521 2202 13577 2204
rect 13601 2202 13657 2204
rect 13361 2150 13407 2202
rect 13407 2150 13417 2202
rect 13441 2150 13471 2202
rect 13471 2150 13483 2202
rect 13483 2150 13497 2202
rect 13521 2150 13535 2202
rect 13535 2150 13547 2202
rect 13547 2150 13577 2202
rect 13601 2150 13611 2202
rect 13611 2150 13657 2202
rect 13361 2148 13417 2150
rect 13441 2148 13497 2150
rect 13521 2148 13577 2150
rect 13601 2148 13657 2150
rect 15212 1658 15268 1660
rect 15292 1658 15348 1660
rect 15372 1658 15428 1660
rect 15452 1658 15508 1660
rect 15212 1606 15258 1658
rect 15258 1606 15268 1658
rect 15292 1606 15322 1658
rect 15322 1606 15334 1658
rect 15334 1606 15348 1658
rect 15372 1606 15386 1658
rect 15386 1606 15398 1658
rect 15398 1606 15428 1658
rect 15452 1606 15462 1658
rect 15462 1606 15508 1658
rect 15212 1604 15268 1606
rect 15292 1604 15348 1606
rect 15372 1604 15428 1606
rect 15452 1604 15508 1606
rect 12346 1264 12402 1320
rect 2255 1114 2311 1116
rect 2335 1114 2391 1116
rect 2415 1114 2471 1116
rect 2495 1114 2551 1116
rect 2255 1062 2301 1114
rect 2301 1062 2311 1114
rect 2335 1062 2365 1114
rect 2365 1062 2377 1114
rect 2377 1062 2391 1114
rect 2415 1062 2429 1114
rect 2429 1062 2441 1114
rect 2441 1062 2471 1114
rect 2495 1062 2505 1114
rect 2505 1062 2551 1114
rect 2255 1060 2311 1062
rect 2335 1060 2391 1062
rect 2415 1060 2471 1062
rect 2495 1060 2551 1062
rect 5957 1114 6013 1116
rect 6037 1114 6093 1116
rect 6117 1114 6173 1116
rect 6197 1114 6253 1116
rect 5957 1062 6003 1114
rect 6003 1062 6013 1114
rect 6037 1062 6067 1114
rect 6067 1062 6079 1114
rect 6079 1062 6093 1114
rect 6117 1062 6131 1114
rect 6131 1062 6143 1114
rect 6143 1062 6173 1114
rect 6197 1062 6207 1114
rect 6207 1062 6253 1114
rect 5957 1060 6013 1062
rect 6037 1060 6093 1062
rect 6117 1060 6173 1062
rect 6197 1060 6253 1062
rect 9659 1114 9715 1116
rect 9739 1114 9795 1116
rect 9819 1114 9875 1116
rect 9899 1114 9955 1116
rect 9659 1062 9705 1114
rect 9705 1062 9715 1114
rect 9739 1062 9769 1114
rect 9769 1062 9781 1114
rect 9781 1062 9795 1114
rect 9819 1062 9833 1114
rect 9833 1062 9845 1114
rect 9845 1062 9875 1114
rect 9899 1062 9909 1114
rect 9909 1062 9955 1114
rect 9659 1060 9715 1062
rect 9739 1060 9795 1062
rect 9819 1060 9875 1062
rect 9899 1060 9955 1062
rect 13361 1114 13417 1116
rect 13441 1114 13497 1116
rect 13521 1114 13577 1116
rect 13601 1114 13657 1116
rect 13361 1062 13407 1114
rect 13407 1062 13417 1114
rect 13441 1062 13471 1114
rect 13471 1062 13483 1114
rect 13483 1062 13497 1114
rect 13521 1062 13535 1114
rect 13535 1062 13547 1114
rect 13547 1062 13577 1114
rect 13601 1062 13611 1114
rect 13611 1062 13657 1114
rect 13361 1060 13417 1062
rect 13441 1060 13497 1062
rect 13521 1060 13577 1062
rect 13601 1060 13657 1062
rect 4106 570 4162 572
rect 4186 570 4242 572
rect 4266 570 4322 572
rect 4346 570 4402 572
rect 4106 518 4152 570
rect 4152 518 4162 570
rect 4186 518 4216 570
rect 4216 518 4228 570
rect 4228 518 4242 570
rect 4266 518 4280 570
rect 4280 518 4292 570
rect 4292 518 4322 570
rect 4346 518 4356 570
rect 4356 518 4402 570
rect 4106 516 4162 518
rect 4186 516 4242 518
rect 4266 516 4322 518
rect 4346 516 4402 518
rect 7808 570 7864 572
rect 7888 570 7944 572
rect 7968 570 8024 572
rect 8048 570 8104 572
rect 7808 518 7854 570
rect 7854 518 7864 570
rect 7888 518 7918 570
rect 7918 518 7930 570
rect 7930 518 7944 570
rect 7968 518 7982 570
rect 7982 518 7994 570
rect 7994 518 8024 570
rect 8048 518 8058 570
rect 8058 518 8104 570
rect 7808 516 7864 518
rect 7888 516 7944 518
rect 7968 516 8024 518
rect 8048 516 8104 518
rect 11510 570 11566 572
rect 11590 570 11646 572
rect 11670 570 11726 572
rect 11750 570 11806 572
rect 11510 518 11556 570
rect 11556 518 11566 570
rect 11590 518 11620 570
rect 11620 518 11632 570
rect 11632 518 11646 570
rect 11670 518 11684 570
rect 11684 518 11696 570
rect 11696 518 11726 570
rect 11750 518 11760 570
rect 11760 518 11806 570
rect 11510 516 11566 518
rect 11590 516 11646 518
rect 11670 516 11726 518
rect 11750 516 11806 518
rect 15212 570 15268 572
rect 15292 570 15348 572
rect 15372 570 15428 572
rect 15452 570 15508 572
rect 15212 518 15258 570
rect 15258 518 15268 570
rect 15292 518 15322 570
rect 15322 518 15334 570
rect 15334 518 15348 570
rect 15372 518 15386 570
rect 15386 518 15398 570
rect 15398 518 15428 570
rect 15452 518 15462 570
rect 15462 518 15508 570
rect 15212 516 15268 518
rect 15292 516 15348 518
rect 15372 516 15428 518
rect 15452 516 15508 518
<< metal3 >>
rect 2245 15264 2561 15265
rect 2245 15200 2251 15264
rect 2315 15200 2331 15264
rect 2395 15200 2411 15264
rect 2475 15200 2491 15264
rect 2555 15200 2561 15264
rect 2245 15199 2561 15200
rect 5947 15264 6263 15265
rect 5947 15200 5953 15264
rect 6017 15200 6033 15264
rect 6097 15200 6113 15264
rect 6177 15200 6193 15264
rect 6257 15200 6263 15264
rect 5947 15199 6263 15200
rect 9649 15264 9965 15265
rect 9649 15200 9655 15264
rect 9719 15200 9735 15264
rect 9799 15200 9815 15264
rect 9879 15200 9895 15264
rect 9959 15200 9965 15264
rect 9649 15199 9965 15200
rect 13351 15264 13667 15265
rect 13351 15200 13357 15264
rect 13421 15200 13437 15264
rect 13501 15200 13517 15264
rect 13581 15200 13597 15264
rect 13661 15200 13667 15264
rect 13351 15199 13667 15200
rect 4096 14720 4412 14721
rect 4096 14656 4102 14720
rect 4166 14656 4182 14720
rect 4246 14656 4262 14720
rect 4326 14656 4342 14720
rect 4406 14656 4412 14720
rect 4096 14655 4412 14656
rect 7798 14720 8114 14721
rect 7798 14656 7804 14720
rect 7868 14656 7884 14720
rect 7948 14656 7964 14720
rect 8028 14656 8044 14720
rect 8108 14656 8114 14720
rect 7798 14655 8114 14656
rect 11500 14720 11816 14721
rect 11500 14656 11506 14720
rect 11570 14656 11586 14720
rect 11650 14656 11666 14720
rect 11730 14656 11746 14720
rect 11810 14656 11816 14720
rect 11500 14655 11816 14656
rect 15202 14720 15518 14721
rect 15202 14656 15208 14720
rect 15272 14656 15288 14720
rect 15352 14656 15368 14720
rect 15432 14656 15448 14720
rect 15512 14656 15518 14720
rect 15202 14655 15518 14656
rect 15009 14514 15075 14517
rect 15600 14514 16000 14544
rect 15009 14512 16000 14514
rect 15009 14456 15014 14512
rect 15070 14456 16000 14512
rect 15009 14454 16000 14456
rect 15009 14451 15075 14454
rect 15600 14424 16000 14454
rect 2245 14176 2561 14177
rect 2245 14112 2251 14176
rect 2315 14112 2331 14176
rect 2395 14112 2411 14176
rect 2475 14112 2491 14176
rect 2555 14112 2561 14176
rect 2245 14111 2561 14112
rect 5947 14176 6263 14177
rect 5947 14112 5953 14176
rect 6017 14112 6033 14176
rect 6097 14112 6113 14176
rect 6177 14112 6193 14176
rect 6257 14112 6263 14176
rect 5947 14111 6263 14112
rect 9649 14176 9965 14177
rect 9649 14112 9655 14176
rect 9719 14112 9735 14176
rect 9799 14112 9815 14176
rect 9879 14112 9895 14176
rect 9959 14112 9965 14176
rect 9649 14111 9965 14112
rect 13351 14176 13667 14177
rect 13351 14112 13357 14176
rect 13421 14112 13437 14176
rect 13501 14112 13517 14176
rect 13581 14112 13597 14176
rect 13661 14112 13667 14176
rect 13351 14111 13667 14112
rect 4096 13632 4412 13633
rect 4096 13568 4102 13632
rect 4166 13568 4182 13632
rect 4246 13568 4262 13632
rect 4326 13568 4342 13632
rect 4406 13568 4412 13632
rect 4096 13567 4412 13568
rect 7798 13632 8114 13633
rect 7798 13568 7804 13632
rect 7868 13568 7884 13632
rect 7948 13568 7964 13632
rect 8028 13568 8044 13632
rect 8108 13568 8114 13632
rect 7798 13567 8114 13568
rect 11500 13632 11816 13633
rect 11500 13568 11506 13632
rect 11570 13568 11586 13632
rect 11650 13568 11666 13632
rect 11730 13568 11746 13632
rect 11810 13568 11816 13632
rect 11500 13567 11816 13568
rect 15202 13632 15518 13633
rect 15202 13568 15208 13632
rect 15272 13568 15288 13632
rect 15352 13568 15368 13632
rect 15432 13568 15448 13632
rect 15512 13568 15518 13632
rect 15202 13567 15518 13568
rect 2245 13088 2561 13089
rect 2245 13024 2251 13088
rect 2315 13024 2331 13088
rect 2395 13024 2411 13088
rect 2475 13024 2491 13088
rect 2555 13024 2561 13088
rect 2245 13023 2561 13024
rect 5947 13088 6263 13089
rect 5947 13024 5953 13088
rect 6017 13024 6033 13088
rect 6097 13024 6113 13088
rect 6177 13024 6193 13088
rect 6257 13024 6263 13088
rect 5947 13023 6263 13024
rect 9649 13088 9965 13089
rect 9649 13024 9655 13088
rect 9719 13024 9735 13088
rect 9799 13024 9815 13088
rect 9879 13024 9895 13088
rect 9959 13024 9965 13088
rect 9649 13023 9965 13024
rect 13351 13088 13667 13089
rect 13351 13024 13357 13088
rect 13421 13024 13437 13088
rect 13501 13024 13517 13088
rect 13581 13024 13597 13088
rect 13661 13024 13667 13088
rect 13351 13023 13667 13024
rect 12985 12746 13051 12749
rect 14457 12746 14523 12749
rect 12985 12744 14523 12746
rect 12985 12688 12990 12744
rect 13046 12688 14462 12744
rect 14518 12688 14523 12744
rect 12985 12686 14523 12688
rect 12985 12683 13051 12686
rect 14457 12683 14523 12686
rect 13445 12610 13511 12613
rect 13997 12610 14063 12613
rect 13445 12608 14063 12610
rect 13445 12552 13450 12608
rect 13506 12552 14002 12608
rect 14058 12552 14063 12608
rect 13445 12550 14063 12552
rect 13445 12547 13511 12550
rect 13997 12547 14063 12550
rect 4096 12544 4412 12545
rect 4096 12480 4102 12544
rect 4166 12480 4182 12544
rect 4246 12480 4262 12544
rect 4326 12480 4342 12544
rect 4406 12480 4412 12544
rect 4096 12479 4412 12480
rect 7798 12544 8114 12545
rect 7798 12480 7804 12544
rect 7868 12480 7884 12544
rect 7948 12480 7964 12544
rect 8028 12480 8044 12544
rect 8108 12480 8114 12544
rect 7798 12479 8114 12480
rect 11500 12544 11816 12545
rect 11500 12480 11506 12544
rect 11570 12480 11586 12544
rect 11650 12480 11666 12544
rect 11730 12480 11746 12544
rect 11810 12480 11816 12544
rect 11500 12479 11816 12480
rect 15202 12544 15518 12545
rect 15202 12480 15208 12544
rect 15272 12480 15288 12544
rect 15352 12480 15368 12544
rect 15432 12480 15448 12544
rect 15512 12480 15518 12544
rect 15600 12520 16000 12640
rect 15202 12479 15518 12480
rect 15009 12338 15075 12341
rect 15702 12338 15762 12520
rect 15009 12336 15762 12338
rect 15009 12280 15014 12336
rect 15070 12280 15762 12336
rect 15009 12278 15762 12280
rect 15009 12275 15075 12278
rect 2245 12000 2561 12001
rect 2245 11936 2251 12000
rect 2315 11936 2331 12000
rect 2395 11936 2411 12000
rect 2475 11936 2491 12000
rect 2555 11936 2561 12000
rect 2245 11935 2561 11936
rect 5947 12000 6263 12001
rect 5947 11936 5953 12000
rect 6017 11936 6033 12000
rect 6097 11936 6113 12000
rect 6177 11936 6193 12000
rect 6257 11936 6263 12000
rect 5947 11935 6263 11936
rect 9649 12000 9965 12001
rect 9649 11936 9655 12000
rect 9719 11936 9735 12000
rect 9799 11936 9815 12000
rect 9879 11936 9895 12000
rect 9959 11936 9965 12000
rect 9649 11935 9965 11936
rect 13351 12000 13667 12001
rect 13351 11936 13357 12000
rect 13421 11936 13437 12000
rect 13501 11936 13517 12000
rect 13581 11936 13597 12000
rect 13661 11936 13667 12000
rect 13351 11935 13667 11936
rect 4096 11456 4412 11457
rect 4096 11392 4102 11456
rect 4166 11392 4182 11456
rect 4246 11392 4262 11456
rect 4326 11392 4342 11456
rect 4406 11392 4412 11456
rect 4096 11391 4412 11392
rect 7798 11456 8114 11457
rect 7798 11392 7804 11456
rect 7868 11392 7884 11456
rect 7948 11392 7964 11456
rect 8028 11392 8044 11456
rect 8108 11392 8114 11456
rect 7798 11391 8114 11392
rect 11500 11456 11816 11457
rect 11500 11392 11506 11456
rect 11570 11392 11586 11456
rect 11650 11392 11666 11456
rect 11730 11392 11746 11456
rect 11810 11392 11816 11456
rect 11500 11391 11816 11392
rect 15202 11456 15518 11457
rect 15202 11392 15208 11456
rect 15272 11392 15288 11456
rect 15352 11392 15368 11456
rect 15432 11392 15448 11456
rect 15512 11392 15518 11456
rect 15202 11391 15518 11392
rect 3509 11250 3575 11253
rect 4061 11250 4127 11253
rect 4613 11250 4679 11253
rect 5257 11250 5323 11253
rect 3509 11248 5323 11250
rect 3509 11192 3514 11248
rect 3570 11192 4066 11248
rect 4122 11192 4618 11248
rect 4674 11192 5262 11248
rect 5318 11192 5323 11248
rect 3509 11190 5323 11192
rect 3509 11187 3575 11190
rect 4061 11187 4127 11190
rect 4613 11187 4679 11190
rect 5257 11187 5323 11190
rect 4521 11114 4587 11117
rect 4981 11114 5047 11117
rect 4521 11112 5047 11114
rect 4521 11056 4526 11112
rect 4582 11056 4986 11112
rect 5042 11056 5047 11112
rect 4521 11054 5047 11056
rect 4521 11051 4587 11054
rect 4981 11051 5047 11054
rect 2245 10912 2561 10913
rect 2245 10848 2251 10912
rect 2315 10848 2331 10912
rect 2395 10848 2411 10912
rect 2475 10848 2491 10912
rect 2555 10848 2561 10912
rect 2245 10847 2561 10848
rect 5947 10912 6263 10913
rect 5947 10848 5953 10912
rect 6017 10848 6033 10912
rect 6097 10848 6113 10912
rect 6177 10848 6193 10912
rect 6257 10848 6263 10912
rect 5947 10847 6263 10848
rect 9649 10912 9965 10913
rect 9649 10848 9655 10912
rect 9719 10848 9735 10912
rect 9799 10848 9815 10912
rect 9879 10848 9895 10912
rect 9959 10848 9965 10912
rect 9649 10847 9965 10848
rect 13351 10912 13667 10913
rect 13351 10848 13357 10912
rect 13421 10848 13437 10912
rect 13501 10848 13517 10912
rect 13581 10848 13597 10912
rect 13661 10848 13667 10912
rect 13351 10847 13667 10848
rect 12341 10706 12407 10709
rect 14181 10706 14247 10709
rect 12341 10704 14247 10706
rect 12341 10648 12346 10704
rect 12402 10648 14186 10704
rect 14242 10648 14247 10704
rect 12341 10646 14247 10648
rect 12341 10643 12407 10646
rect 14181 10643 14247 10646
rect 14917 10706 14983 10709
rect 15600 10706 16000 10736
rect 14917 10704 16000 10706
rect 14917 10648 14922 10704
rect 14978 10648 16000 10704
rect 14917 10646 16000 10648
rect 14917 10643 14983 10646
rect 15600 10616 16000 10646
rect 4096 10368 4412 10369
rect 4096 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4342 10368
rect 4406 10304 4412 10368
rect 4096 10303 4412 10304
rect 7798 10368 8114 10369
rect 7798 10304 7804 10368
rect 7868 10304 7884 10368
rect 7948 10304 7964 10368
rect 8028 10304 8044 10368
rect 8108 10304 8114 10368
rect 7798 10303 8114 10304
rect 11500 10368 11816 10369
rect 11500 10304 11506 10368
rect 11570 10304 11586 10368
rect 11650 10304 11666 10368
rect 11730 10304 11746 10368
rect 11810 10304 11816 10368
rect 11500 10303 11816 10304
rect 15202 10368 15518 10369
rect 15202 10304 15208 10368
rect 15272 10304 15288 10368
rect 15352 10304 15368 10368
rect 15432 10304 15448 10368
rect 15512 10304 15518 10368
rect 15202 10303 15518 10304
rect 2245 9824 2561 9825
rect 2245 9760 2251 9824
rect 2315 9760 2331 9824
rect 2395 9760 2411 9824
rect 2475 9760 2491 9824
rect 2555 9760 2561 9824
rect 2245 9759 2561 9760
rect 5947 9824 6263 9825
rect 5947 9760 5953 9824
rect 6017 9760 6033 9824
rect 6097 9760 6113 9824
rect 6177 9760 6193 9824
rect 6257 9760 6263 9824
rect 5947 9759 6263 9760
rect 9649 9824 9965 9825
rect 9649 9760 9655 9824
rect 9719 9760 9735 9824
rect 9799 9760 9815 9824
rect 9879 9760 9895 9824
rect 9959 9760 9965 9824
rect 9649 9759 9965 9760
rect 13351 9824 13667 9825
rect 13351 9760 13357 9824
rect 13421 9760 13437 9824
rect 13501 9760 13517 9824
rect 13581 9760 13597 9824
rect 13661 9760 13667 9824
rect 13351 9759 13667 9760
rect 4096 9280 4412 9281
rect 4096 9216 4102 9280
rect 4166 9216 4182 9280
rect 4246 9216 4262 9280
rect 4326 9216 4342 9280
rect 4406 9216 4412 9280
rect 4096 9215 4412 9216
rect 7798 9280 8114 9281
rect 7798 9216 7804 9280
rect 7868 9216 7884 9280
rect 7948 9216 7964 9280
rect 8028 9216 8044 9280
rect 8108 9216 8114 9280
rect 7798 9215 8114 9216
rect 11500 9280 11816 9281
rect 11500 9216 11506 9280
rect 11570 9216 11586 9280
rect 11650 9216 11666 9280
rect 11730 9216 11746 9280
rect 11810 9216 11816 9280
rect 11500 9215 11816 9216
rect 15202 9280 15518 9281
rect 15202 9216 15208 9280
rect 15272 9216 15288 9280
rect 15352 9216 15368 9280
rect 15432 9216 15448 9280
rect 15512 9216 15518 9280
rect 15202 9215 15518 9216
rect 6361 9074 6427 9077
rect 9305 9074 9371 9077
rect 9581 9074 9647 9077
rect 12433 9074 12499 9077
rect 6361 9072 12499 9074
rect 6361 9016 6366 9072
rect 6422 9016 9310 9072
rect 9366 9016 9586 9072
rect 9642 9016 12438 9072
rect 12494 9016 12499 9072
rect 6361 9014 12499 9016
rect 6361 9011 6427 9014
rect 9305 9011 9371 9014
rect 9581 9011 9647 9014
rect 12433 9011 12499 9014
rect 15009 8802 15075 8805
rect 15600 8802 16000 8832
rect 15009 8800 16000 8802
rect 15009 8744 15014 8800
rect 15070 8744 16000 8800
rect 15009 8742 16000 8744
rect 15009 8739 15075 8742
rect 2245 8736 2561 8737
rect 2245 8672 2251 8736
rect 2315 8672 2331 8736
rect 2395 8672 2411 8736
rect 2475 8672 2491 8736
rect 2555 8672 2561 8736
rect 2245 8671 2561 8672
rect 5947 8736 6263 8737
rect 5947 8672 5953 8736
rect 6017 8672 6033 8736
rect 6097 8672 6113 8736
rect 6177 8672 6193 8736
rect 6257 8672 6263 8736
rect 5947 8671 6263 8672
rect 9649 8736 9965 8737
rect 9649 8672 9655 8736
rect 9719 8672 9735 8736
rect 9799 8672 9815 8736
rect 9879 8672 9895 8736
rect 9959 8672 9965 8736
rect 9649 8671 9965 8672
rect 13351 8736 13667 8737
rect 13351 8672 13357 8736
rect 13421 8672 13437 8736
rect 13501 8672 13517 8736
rect 13581 8672 13597 8736
rect 13661 8672 13667 8736
rect 15600 8712 16000 8742
rect 13351 8671 13667 8672
rect 4096 8192 4412 8193
rect 4096 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4342 8192
rect 4406 8128 4412 8192
rect 4096 8127 4412 8128
rect 7798 8192 8114 8193
rect 7798 8128 7804 8192
rect 7868 8128 7884 8192
rect 7948 8128 7964 8192
rect 8028 8128 8044 8192
rect 8108 8128 8114 8192
rect 7798 8127 8114 8128
rect 11500 8192 11816 8193
rect 11500 8128 11506 8192
rect 11570 8128 11586 8192
rect 11650 8128 11666 8192
rect 11730 8128 11746 8192
rect 11810 8128 11816 8192
rect 11500 8127 11816 8128
rect 15202 8192 15518 8193
rect 15202 8128 15208 8192
rect 15272 8128 15288 8192
rect 15352 8128 15368 8192
rect 15432 8128 15448 8192
rect 15512 8128 15518 8192
rect 15202 8127 15518 8128
rect 2245 7648 2561 7649
rect 2245 7584 2251 7648
rect 2315 7584 2331 7648
rect 2395 7584 2411 7648
rect 2475 7584 2491 7648
rect 2555 7584 2561 7648
rect 2245 7583 2561 7584
rect 5947 7648 6263 7649
rect 5947 7584 5953 7648
rect 6017 7584 6033 7648
rect 6097 7584 6113 7648
rect 6177 7584 6193 7648
rect 6257 7584 6263 7648
rect 5947 7583 6263 7584
rect 9649 7648 9965 7649
rect 9649 7584 9655 7648
rect 9719 7584 9735 7648
rect 9799 7584 9815 7648
rect 9879 7584 9895 7648
rect 9959 7584 9965 7648
rect 9649 7583 9965 7584
rect 13351 7648 13667 7649
rect 13351 7584 13357 7648
rect 13421 7584 13437 7648
rect 13501 7584 13517 7648
rect 13581 7584 13597 7648
rect 13661 7584 13667 7648
rect 13351 7583 13667 7584
rect 7833 7306 7899 7309
rect 12157 7306 12223 7309
rect 13261 7306 13327 7309
rect 7833 7304 13327 7306
rect 7833 7248 7838 7304
rect 7894 7248 12162 7304
rect 12218 7248 13266 7304
rect 13322 7248 13327 7304
rect 7833 7246 13327 7248
rect 7833 7243 7899 7246
rect 12157 7243 12223 7246
rect 13261 7243 13327 7246
rect 4096 7104 4412 7105
rect 4096 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4342 7104
rect 4406 7040 4412 7104
rect 4096 7039 4412 7040
rect 7798 7104 8114 7105
rect 7798 7040 7804 7104
rect 7868 7040 7884 7104
rect 7948 7040 7964 7104
rect 8028 7040 8044 7104
rect 8108 7040 8114 7104
rect 7798 7039 8114 7040
rect 11500 7104 11816 7105
rect 11500 7040 11506 7104
rect 11570 7040 11586 7104
rect 11650 7040 11666 7104
rect 11730 7040 11746 7104
rect 11810 7040 11816 7104
rect 11500 7039 11816 7040
rect 15202 7104 15518 7105
rect 15202 7040 15208 7104
rect 15272 7040 15288 7104
rect 15352 7040 15368 7104
rect 15432 7040 15448 7104
rect 15512 7040 15518 7104
rect 15202 7039 15518 7040
rect 15009 6898 15075 6901
rect 15600 6898 16000 6928
rect 15009 6896 16000 6898
rect 15009 6840 15014 6896
rect 15070 6840 16000 6896
rect 15009 6838 16000 6840
rect 15009 6835 15075 6838
rect 15600 6808 16000 6838
rect 2245 6560 2561 6561
rect 2245 6496 2251 6560
rect 2315 6496 2331 6560
rect 2395 6496 2411 6560
rect 2475 6496 2491 6560
rect 2555 6496 2561 6560
rect 2245 6495 2561 6496
rect 5947 6560 6263 6561
rect 5947 6496 5953 6560
rect 6017 6496 6033 6560
rect 6097 6496 6113 6560
rect 6177 6496 6193 6560
rect 6257 6496 6263 6560
rect 5947 6495 6263 6496
rect 9649 6560 9965 6561
rect 9649 6496 9655 6560
rect 9719 6496 9735 6560
rect 9799 6496 9815 6560
rect 9879 6496 9895 6560
rect 9959 6496 9965 6560
rect 9649 6495 9965 6496
rect 13351 6560 13667 6561
rect 13351 6496 13357 6560
rect 13421 6496 13437 6560
rect 13501 6496 13517 6560
rect 13581 6496 13597 6560
rect 13661 6496 13667 6560
rect 13351 6495 13667 6496
rect 8845 6354 8911 6357
rect 10041 6354 10107 6357
rect 8845 6352 10107 6354
rect 8845 6296 8850 6352
rect 8906 6296 10046 6352
rect 10102 6296 10107 6352
rect 8845 6294 10107 6296
rect 8845 6291 8911 6294
rect 10041 6291 10107 6294
rect 4096 6016 4412 6017
rect 4096 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4342 6016
rect 4406 5952 4412 6016
rect 4096 5951 4412 5952
rect 7798 6016 8114 6017
rect 7798 5952 7804 6016
rect 7868 5952 7884 6016
rect 7948 5952 7964 6016
rect 8028 5952 8044 6016
rect 8108 5952 8114 6016
rect 7798 5951 8114 5952
rect 11500 6016 11816 6017
rect 11500 5952 11506 6016
rect 11570 5952 11586 6016
rect 11650 5952 11666 6016
rect 11730 5952 11746 6016
rect 11810 5952 11816 6016
rect 11500 5951 11816 5952
rect 15202 6016 15518 6017
rect 15202 5952 15208 6016
rect 15272 5952 15288 6016
rect 15352 5952 15368 6016
rect 15432 5952 15448 6016
rect 15512 5952 15518 6016
rect 15202 5951 15518 5952
rect 14457 5538 14523 5541
rect 14457 5536 15762 5538
rect 14457 5480 14462 5536
rect 14518 5480 15762 5536
rect 14457 5478 15762 5480
rect 14457 5475 14523 5478
rect 2245 5472 2561 5473
rect 2245 5408 2251 5472
rect 2315 5408 2331 5472
rect 2395 5408 2411 5472
rect 2475 5408 2491 5472
rect 2555 5408 2561 5472
rect 2245 5407 2561 5408
rect 5947 5472 6263 5473
rect 5947 5408 5953 5472
rect 6017 5408 6033 5472
rect 6097 5408 6113 5472
rect 6177 5408 6193 5472
rect 6257 5408 6263 5472
rect 5947 5407 6263 5408
rect 9649 5472 9965 5473
rect 9649 5408 9655 5472
rect 9719 5408 9735 5472
rect 9799 5408 9815 5472
rect 9879 5408 9895 5472
rect 9959 5408 9965 5472
rect 9649 5407 9965 5408
rect 13351 5472 13667 5473
rect 13351 5408 13357 5472
rect 13421 5408 13437 5472
rect 13501 5408 13517 5472
rect 13581 5408 13597 5472
rect 13661 5408 13667 5472
rect 13351 5407 13667 5408
rect 15702 5024 15762 5478
rect 4096 4928 4412 4929
rect 4096 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4342 4928
rect 4406 4864 4412 4928
rect 4096 4863 4412 4864
rect 7798 4928 8114 4929
rect 7798 4864 7804 4928
rect 7868 4864 7884 4928
rect 7948 4864 7964 4928
rect 8028 4864 8044 4928
rect 8108 4864 8114 4928
rect 7798 4863 8114 4864
rect 11500 4928 11816 4929
rect 11500 4864 11506 4928
rect 11570 4864 11586 4928
rect 11650 4864 11666 4928
rect 11730 4864 11746 4928
rect 11810 4864 11816 4928
rect 11500 4863 11816 4864
rect 15202 4928 15518 4929
rect 15202 4864 15208 4928
rect 15272 4864 15288 4928
rect 15352 4864 15368 4928
rect 15432 4864 15448 4928
rect 15512 4864 15518 4928
rect 15600 4904 16000 5024
rect 15202 4863 15518 4864
rect 2245 4384 2561 4385
rect 2245 4320 2251 4384
rect 2315 4320 2331 4384
rect 2395 4320 2411 4384
rect 2475 4320 2491 4384
rect 2555 4320 2561 4384
rect 2245 4319 2561 4320
rect 5947 4384 6263 4385
rect 5947 4320 5953 4384
rect 6017 4320 6033 4384
rect 6097 4320 6113 4384
rect 6177 4320 6193 4384
rect 6257 4320 6263 4384
rect 5947 4319 6263 4320
rect 9649 4384 9965 4385
rect 9649 4320 9655 4384
rect 9719 4320 9735 4384
rect 9799 4320 9815 4384
rect 9879 4320 9895 4384
rect 9959 4320 9965 4384
rect 9649 4319 9965 4320
rect 13351 4384 13667 4385
rect 13351 4320 13357 4384
rect 13421 4320 13437 4384
rect 13501 4320 13517 4384
rect 13581 4320 13597 4384
rect 13661 4320 13667 4384
rect 13351 4319 13667 4320
rect 4096 3840 4412 3841
rect 4096 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4342 3840
rect 4406 3776 4412 3840
rect 4096 3775 4412 3776
rect 7798 3840 8114 3841
rect 7798 3776 7804 3840
rect 7868 3776 7884 3840
rect 7948 3776 7964 3840
rect 8028 3776 8044 3840
rect 8108 3776 8114 3840
rect 7798 3775 8114 3776
rect 11500 3840 11816 3841
rect 11500 3776 11506 3840
rect 11570 3776 11586 3840
rect 11650 3776 11666 3840
rect 11730 3776 11746 3840
rect 11810 3776 11816 3840
rect 11500 3775 11816 3776
rect 15202 3840 15518 3841
rect 15202 3776 15208 3840
rect 15272 3776 15288 3840
rect 15352 3776 15368 3840
rect 15432 3776 15448 3840
rect 15512 3776 15518 3840
rect 15202 3775 15518 3776
rect 2245 3296 2561 3297
rect 2245 3232 2251 3296
rect 2315 3232 2331 3296
rect 2395 3232 2411 3296
rect 2475 3232 2491 3296
rect 2555 3232 2561 3296
rect 2245 3231 2561 3232
rect 5947 3296 6263 3297
rect 5947 3232 5953 3296
rect 6017 3232 6033 3296
rect 6097 3232 6113 3296
rect 6177 3232 6193 3296
rect 6257 3232 6263 3296
rect 5947 3231 6263 3232
rect 9649 3296 9965 3297
rect 9649 3232 9655 3296
rect 9719 3232 9735 3296
rect 9799 3232 9815 3296
rect 9879 3232 9895 3296
rect 9959 3232 9965 3296
rect 9649 3231 9965 3232
rect 13351 3296 13667 3297
rect 13351 3232 13357 3296
rect 13421 3232 13437 3296
rect 13501 3232 13517 3296
rect 13581 3232 13597 3296
rect 13661 3232 13667 3296
rect 13351 3231 13667 3232
rect 14549 3090 14615 3093
rect 15600 3090 16000 3120
rect 14549 3088 16000 3090
rect 14549 3032 14554 3088
rect 14610 3032 16000 3088
rect 14549 3030 16000 3032
rect 14549 3027 14615 3030
rect 15600 3000 16000 3030
rect 4096 2752 4412 2753
rect 4096 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4342 2752
rect 4406 2688 4412 2752
rect 4096 2687 4412 2688
rect 7798 2752 8114 2753
rect 7798 2688 7804 2752
rect 7868 2688 7884 2752
rect 7948 2688 7964 2752
rect 8028 2688 8044 2752
rect 8108 2688 8114 2752
rect 7798 2687 8114 2688
rect 11500 2752 11816 2753
rect 11500 2688 11506 2752
rect 11570 2688 11586 2752
rect 11650 2688 11666 2752
rect 11730 2688 11746 2752
rect 11810 2688 11816 2752
rect 11500 2687 11816 2688
rect 15202 2752 15518 2753
rect 15202 2688 15208 2752
rect 15272 2688 15288 2752
rect 15352 2688 15368 2752
rect 15432 2688 15448 2752
rect 15512 2688 15518 2752
rect 15202 2687 15518 2688
rect 2245 2208 2561 2209
rect 2245 2144 2251 2208
rect 2315 2144 2331 2208
rect 2395 2144 2411 2208
rect 2475 2144 2491 2208
rect 2555 2144 2561 2208
rect 2245 2143 2561 2144
rect 5947 2208 6263 2209
rect 5947 2144 5953 2208
rect 6017 2144 6033 2208
rect 6097 2144 6113 2208
rect 6177 2144 6193 2208
rect 6257 2144 6263 2208
rect 5947 2143 6263 2144
rect 9649 2208 9965 2209
rect 9649 2144 9655 2208
rect 9719 2144 9735 2208
rect 9799 2144 9815 2208
rect 9879 2144 9895 2208
rect 9959 2144 9965 2208
rect 9649 2143 9965 2144
rect 13351 2208 13667 2209
rect 13351 2144 13357 2208
rect 13421 2144 13437 2208
rect 13501 2144 13517 2208
rect 13581 2144 13597 2208
rect 13661 2144 13667 2208
rect 13351 2143 13667 2144
rect 4096 1664 4412 1665
rect 4096 1600 4102 1664
rect 4166 1600 4182 1664
rect 4246 1600 4262 1664
rect 4326 1600 4342 1664
rect 4406 1600 4412 1664
rect 4096 1599 4412 1600
rect 7798 1664 8114 1665
rect 7798 1600 7804 1664
rect 7868 1600 7884 1664
rect 7948 1600 7964 1664
rect 8028 1600 8044 1664
rect 8108 1600 8114 1664
rect 7798 1599 8114 1600
rect 11500 1664 11816 1665
rect 11500 1600 11506 1664
rect 11570 1600 11586 1664
rect 11650 1600 11666 1664
rect 11730 1600 11746 1664
rect 11810 1600 11816 1664
rect 11500 1599 11816 1600
rect 15202 1664 15518 1665
rect 15202 1600 15208 1664
rect 15272 1600 15288 1664
rect 15352 1600 15368 1664
rect 15432 1600 15448 1664
rect 15512 1600 15518 1664
rect 15202 1599 15518 1600
rect 12341 1322 12407 1325
rect 12341 1320 13922 1322
rect 12341 1264 12346 1320
rect 12402 1264 13922 1320
rect 12341 1262 13922 1264
rect 12341 1259 12407 1262
rect 13862 1186 13922 1262
rect 15600 1186 16000 1216
rect 13862 1126 16000 1186
rect 2245 1120 2561 1121
rect 2245 1056 2251 1120
rect 2315 1056 2331 1120
rect 2395 1056 2411 1120
rect 2475 1056 2491 1120
rect 2555 1056 2561 1120
rect 2245 1055 2561 1056
rect 5947 1120 6263 1121
rect 5947 1056 5953 1120
rect 6017 1056 6033 1120
rect 6097 1056 6113 1120
rect 6177 1056 6193 1120
rect 6257 1056 6263 1120
rect 5947 1055 6263 1056
rect 9649 1120 9965 1121
rect 9649 1056 9655 1120
rect 9719 1056 9735 1120
rect 9799 1056 9815 1120
rect 9879 1056 9895 1120
rect 9959 1056 9965 1120
rect 9649 1055 9965 1056
rect 13351 1120 13667 1121
rect 13351 1056 13357 1120
rect 13421 1056 13437 1120
rect 13501 1056 13517 1120
rect 13581 1056 13597 1120
rect 13661 1056 13667 1120
rect 15600 1096 16000 1126
rect 13351 1055 13667 1056
rect 4096 576 4412 577
rect 4096 512 4102 576
rect 4166 512 4182 576
rect 4246 512 4262 576
rect 4326 512 4342 576
rect 4406 512 4412 576
rect 4096 511 4412 512
rect 7798 576 8114 577
rect 7798 512 7804 576
rect 7868 512 7884 576
rect 7948 512 7964 576
rect 8028 512 8044 576
rect 8108 512 8114 576
rect 7798 511 8114 512
rect 11500 576 11816 577
rect 11500 512 11506 576
rect 11570 512 11586 576
rect 11650 512 11666 576
rect 11730 512 11746 576
rect 11810 512 11816 576
rect 11500 511 11816 512
rect 15202 576 15518 577
rect 15202 512 15208 576
rect 15272 512 15288 576
rect 15352 512 15368 576
rect 15432 512 15448 576
rect 15512 512 15518 576
rect 15202 511 15518 512
<< via3 >>
rect 2251 15260 2315 15264
rect 2251 15204 2255 15260
rect 2255 15204 2311 15260
rect 2311 15204 2315 15260
rect 2251 15200 2315 15204
rect 2331 15260 2395 15264
rect 2331 15204 2335 15260
rect 2335 15204 2391 15260
rect 2391 15204 2395 15260
rect 2331 15200 2395 15204
rect 2411 15260 2475 15264
rect 2411 15204 2415 15260
rect 2415 15204 2471 15260
rect 2471 15204 2475 15260
rect 2411 15200 2475 15204
rect 2491 15260 2555 15264
rect 2491 15204 2495 15260
rect 2495 15204 2551 15260
rect 2551 15204 2555 15260
rect 2491 15200 2555 15204
rect 5953 15260 6017 15264
rect 5953 15204 5957 15260
rect 5957 15204 6013 15260
rect 6013 15204 6017 15260
rect 5953 15200 6017 15204
rect 6033 15260 6097 15264
rect 6033 15204 6037 15260
rect 6037 15204 6093 15260
rect 6093 15204 6097 15260
rect 6033 15200 6097 15204
rect 6113 15260 6177 15264
rect 6113 15204 6117 15260
rect 6117 15204 6173 15260
rect 6173 15204 6177 15260
rect 6113 15200 6177 15204
rect 6193 15260 6257 15264
rect 6193 15204 6197 15260
rect 6197 15204 6253 15260
rect 6253 15204 6257 15260
rect 6193 15200 6257 15204
rect 9655 15260 9719 15264
rect 9655 15204 9659 15260
rect 9659 15204 9715 15260
rect 9715 15204 9719 15260
rect 9655 15200 9719 15204
rect 9735 15260 9799 15264
rect 9735 15204 9739 15260
rect 9739 15204 9795 15260
rect 9795 15204 9799 15260
rect 9735 15200 9799 15204
rect 9815 15260 9879 15264
rect 9815 15204 9819 15260
rect 9819 15204 9875 15260
rect 9875 15204 9879 15260
rect 9815 15200 9879 15204
rect 9895 15260 9959 15264
rect 9895 15204 9899 15260
rect 9899 15204 9955 15260
rect 9955 15204 9959 15260
rect 9895 15200 9959 15204
rect 13357 15260 13421 15264
rect 13357 15204 13361 15260
rect 13361 15204 13417 15260
rect 13417 15204 13421 15260
rect 13357 15200 13421 15204
rect 13437 15260 13501 15264
rect 13437 15204 13441 15260
rect 13441 15204 13497 15260
rect 13497 15204 13501 15260
rect 13437 15200 13501 15204
rect 13517 15260 13581 15264
rect 13517 15204 13521 15260
rect 13521 15204 13577 15260
rect 13577 15204 13581 15260
rect 13517 15200 13581 15204
rect 13597 15260 13661 15264
rect 13597 15204 13601 15260
rect 13601 15204 13657 15260
rect 13657 15204 13661 15260
rect 13597 15200 13661 15204
rect 4102 14716 4166 14720
rect 4102 14660 4106 14716
rect 4106 14660 4162 14716
rect 4162 14660 4166 14716
rect 4102 14656 4166 14660
rect 4182 14716 4246 14720
rect 4182 14660 4186 14716
rect 4186 14660 4242 14716
rect 4242 14660 4246 14716
rect 4182 14656 4246 14660
rect 4262 14716 4326 14720
rect 4262 14660 4266 14716
rect 4266 14660 4322 14716
rect 4322 14660 4326 14716
rect 4262 14656 4326 14660
rect 4342 14716 4406 14720
rect 4342 14660 4346 14716
rect 4346 14660 4402 14716
rect 4402 14660 4406 14716
rect 4342 14656 4406 14660
rect 7804 14716 7868 14720
rect 7804 14660 7808 14716
rect 7808 14660 7864 14716
rect 7864 14660 7868 14716
rect 7804 14656 7868 14660
rect 7884 14716 7948 14720
rect 7884 14660 7888 14716
rect 7888 14660 7944 14716
rect 7944 14660 7948 14716
rect 7884 14656 7948 14660
rect 7964 14716 8028 14720
rect 7964 14660 7968 14716
rect 7968 14660 8024 14716
rect 8024 14660 8028 14716
rect 7964 14656 8028 14660
rect 8044 14716 8108 14720
rect 8044 14660 8048 14716
rect 8048 14660 8104 14716
rect 8104 14660 8108 14716
rect 8044 14656 8108 14660
rect 11506 14716 11570 14720
rect 11506 14660 11510 14716
rect 11510 14660 11566 14716
rect 11566 14660 11570 14716
rect 11506 14656 11570 14660
rect 11586 14716 11650 14720
rect 11586 14660 11590 14716
rect 11590 14660 11646 14716
rect 11646 14660 11650 14716
rect 11586 14656 11650 14660
rect 11666 14716 11730 14720
rect 11666 14660 11670 14716
rect 11670 14660 11726 14716
rect 11726 14660 11730 14716
rect 11666 14656 11730 14660
rect 11746 14716 11810 14720
rect 11746 14660 11750 14716
rect 11750 14660 11806 14716
rect 11806 14660 11810 14716
rect 11746 14656 11810 14660
rect 15208 14716 15272 14720
rect 15208 14660 15212 14716
rect 15212 14660 15268 14716
rect 15268 14660 15272 14716
rect 15208 14656 15272 14660
rect 15288 14716 15352 14720
rect 15288 14660 15292 14716
rect 15292 14660 15348 14716
rect 15348 14660 15352 14716
rect 15288 14656 15352 14660
rect 15368 14716 15432 14720
rect 15368 14660 15372 14716
rect 15372 14660 15428 14716
rect 15428 14660 15432 14716
rect 15368 14656 15432 14660
rect 15448 14716 15512 14720
rect 15448 14660 15452 14716
rect 15452 14660 15508 14716
rect 15508 14660 15512 14716
rect 15448 14656 15512 14660
rect 2251 14172 2315 14176
rect 2251 14116 2255 14172
rect 2255 14116 2311 14172
rect 2311 14116 2315 14172
rect 2251 14112 2315 14116
rect 2331 14172 2395 14176
rect 2331 14116 2335 14172
rect 2335 14116 2391 14172
rect 2391 14116 2395 14172
rect 2331 14112 2395 14116
rect 2411 14172 2475 14176
rect 2411 14116 2415 14172
rect 2415 14116 2471 14172
rect 2471 14116 2475 14172
rect 2411 14112 2475 14116
rect 2491 14172 2555 14176
rect 2491 14116 2495 14172
rect 2495 14116 2551 14172
rect 2551 14116 2555 14172
rect 2491 14112 2555 14116
rect 5953 14172 6017 14176
rect 5953 14116 5957 14172
rect 5957 14116 6013 14172
rect 6013 14116 6017 14172
rect 5953 14112 6017 14116
rect 6033 14172 6097 14176
rect 6033 14116 6037 14172
rect 6037 14116 6093 14172
rect 6093 14116 6097 14172
rect 6033 14112 6097 14116
rect 6113 14172 6177 14176
rect 6113 14116 6117 14172
rect 6117 14116 6173 14172
rect 6173 14116 6177 14172
rect 6113 14112 6177 14116
rect 6193 14172 6257 14176
rect 6193 14116 6197 14172
rect 6197 14116 6253 14172
rect 6253 14116 6257 14172
rect 6193 14112 6257 14116
rect 9655 14172 9719 14176
rect 9655 14116 9659 14172
rect 9659 14116 9715 14172
rect 9715 14116 9719 14172
rect 9655 14112 9719 14116
rect 9735 14172 9799 14176
rect 9735 14116 9739 14172
rect 9739 14116 9795 14172
rect 9795 14116 9799 14172
rect 9735 14112 9799 14116
rect 9815 14172 9879 14176
rect 9815 14116 9819 14172
rect 9819 14116 9875 14172
rect 9875 14116 9879 14172
rect 9815 14112 9879 14116
rect 9895 14172 9959 14176
rect 9895 14116 9899 14172
rect 9899 14116 9955 14172
rect 9955 14116 9959 14172
rect 9895 14112 9959 14116
rect 13357 14172 13421 14176
rect 13357 14116 13361 14172
rect 13361 14116 13417 14172
rect 13417 14116 13421 14172
rect 13357 14112 13421 14116
rect 13437 14172 13501 14176
rect 13437 14116 13441 14172
rect 13441 14116 13497 14172
rect 13497 14116 13501 14172
rect 13437 14112 13501 14116
rect 13517 14172 13581 14176
rect 13517 14116 13521 14172
rect 13521 14116 13577 14172
rect 13577 14116 13581 14172
rect 13517 14112 13581 14116
rect 13597 14172 13661 14176
rect 13597 14116 13601 14172
rect 13601 14116 13657 14172
rect 13657 14116 13661 14172
rect 13597 14112 13661 14116
rect 4102 13628 4166 13632
rect 4102 13572 4106 13628
rect 4106 13572 4162 13628
rect 4162 13572 4166 13628
rect 4102 13568 4166 13572
rect 4182 13628 4246 13632
rect 4182 13572 4186 13628
rect 4186 13572 4242 13628
rect 4242 13572 4246 13628
rect 4182 13568 4246 13572
rect 4262 13628 4326 13632
rect 4262 13572 4266 13628
rect 4266 13572 4322 13628
rect 4322 13572 4326 13628
rect 4262 13568 4326 13572
rect 4342 13628 4406 13632
rect 4342 13572 4346 13628
rect 4346 13572 4402 13628
rect 4402 13572 4406 13628
rect 4342 13568 4406 13572
rect 7804 13628 7868 13632
rect 7804 13572 7808 13628
rect 7808 13572 7864 13628
rect 7864 13572 7868 13628
rect 7804 13568 7868 13572
rect 7884 13628 7948 13632
rect 7884 13572 7888 13628
rect 7888 13572 7944 13628
rect 7944 13572 7948 13628
rect 7884 13568 7948 13572
rect 7964 13628 8028 13632
rect 7964 13572 7968 13628
rect 7968 13572 8024 13628
rect 8024 13572 8028 13628
rect 7964 13568 8028 13572
rect 8044 13628 8108 13632
rect 8044 13572 8048 13628
rect 8048 13572 8104 13628
rect 8104 13572 8108 13628
rect 8044 13568 8108 13572
rect 11506 13628 11570 13632
rect 11506 13572 11510 13628
rect 11510 13572 11566 13628
rect 11566 13572 11570 13628
rect 11506 13568 11570 13572
rect 11586 13628 11650 13632
rect 11586 13572 11590 13628
rect 11590 13572 11646 13628
rect 11646 13572 11650 13628
rect 11586 13568 11650 13572
rect 11666 13628 11730 13632
rect 11666 13572 11670 13628
rect 11670 13572 11726 13628
rect 11726 13572 11730 13628
rect 11666 13568 11730 13572
rect 11746 13628 11810 13632
rect 11746 13572 11750 13628
rect 11750 13572 11806 13628
rect 11806 13572 11810 13628
rect 11746 13568 11810 13572
rect 15208 13628 15272 13632
rect 15208 13572 15212 13628
rect 15212 13572 15268 13628
rect 15268 13572 15272 13628
rect 15208 13568 15272 13572
rect 15288 13628 15352 13632
rect 15288 13572 15292 13628
rect 15292 13572 15348 13628
rect 15348 13572 15352 13628
rect 15288 13568 15352 13572
rect 15368 13628 15432 13632
rect 15368 13572 15372 13628
rect 15372 13572 15428 13628
rect 15428 13572 15432 13628
rect 15368 13568 15432 13572
rect 15448 13628 15512 13632
rect 15448 13572 15452 13628
rect 15452 13572 15508 13628
rect 15508 13572 15512 13628
rect 15448 13568 15512 13572
rect 2251 13084 2315 13088
rect 2251 13028 2255 13084
rect 2255 13028 2311 13084
rect 2311 13028 2315 13084
rect 2251 13024 2315 13028
rect 2331 13084 2395 13088
rect 2331 13028 2335 13084
rect 2335 13028 2391 13084
rect 2391 13028 2395 13084
rect 2331 13024 2395 13028
rect 2411 13084 2475 13088
rect 2411 13028 2415 13084
rect 2415 13028 2471 13084
rect 2471 13028 2475 13084
rect 2411 13024 2475 13028
rect 2491 13084 2555 13088
rect 2491 13028 2495 13084
rect 2495 13028 2551 13084
rect 2551 13028 2555 13084
rect 2491 13024 2555 13028
rect 5953 13084 6017 13088
rect 5953 13028 5957 13084
rect 5957 13028 6013 13084
rect 6013 13028 6017 13084
rect 5953 13024 6017 13028
rect 6033 13084 6097 13088
rect 6033 13028 6037 13084
rect 6037 13028 6093 13084
rect 6093 13028 6097 13084
rect 6033 13024 6097 13028
rect 6113 13084 6177 13088
rect 6113 13028 6117 13084
rect 6117 13028 6173 13084
rect 6173 13028 6177 13084
rect 6113 13024 6177 13028
rect 6193 13084 6257 13088
rect 6193 13028 6197 13084
rect 6197 13028 6253 13084
rect 6253 13028 6257 13084
rect 6193 13024 6257 13028
rect 9655 13084 9719 13088
rect 9655 13028 9659 13084
rect 9659 13028 9715 13084
rect 9715 13028 9719 13084
rect 9655 13024 9719 13028
rect 9735 13084 9799 13088
rect 9735 13028 9739 13084
rect 9739 13028 9795 13084
rect 9795 13028 9799 13084
rect 9735 13024 9799 13028
rect 9815 13084 9879 13088
rect 9815 13028 9819 13084
rect 9819 13028 9875 13084
rect 9875 13028 9879 13084
rect 9815 13024 9879 13028
rect 9895 13084 9959 13088
rect 9895 13028 9899 13084
rect 9899 13028 9955 13084
rect 9955 13028 9959 13084
rect 9895 13024 9959 13028
rect 13357 13084 13421 13088
rect 13357 13028 13361 13084
rect 13361 13028 13417 13084
rect 13417 13028 13421 13084
rect 13357 13024 13421 13028
rect 13437 13084 13501 13088
rect 13437 13028 13441 13084
rect 13441 13028 13497 13084
rect 13497 13028 13501 13084
rect 13437 13024 13501 13028
rect 13517 13084 13581 13088
rect 13517 13028 13521 13084
rect 13521 13028 13577 13084
rect 13577 13028 13581 13084
rect 13517 13024 13581 13028
rect 13597 13084 13661 13088
rect 13597 13028 13601 13084
rect 13601 13028 13657 13084
rect 13657 13028 13661 13084
rect 13597 13024 13661 13028
rect 4102 12540 4166 12544
rect 4102 12484 4106 12540
rect 4106 12484 4162 12540
rect 4162 12484 4166 12540
rect 4102 12480 4166 12484
rect 4182 12540 4246 12544
rect 4182 12484 4186 12540
rect 4186 12484 4242 12540
rect 4242 12484 4246 12540
rect 4182 12480 4246 12484
rect 4262 12540 4326 12544
rect 4262 12484 4266 12540
rect 4266 12484 4322 12540
rect 4322 12484 4326 12540
rect 4262 12480 4326 12484
rect 4342 12540 4406 12544
rect 4342 12484 4346 12540
rect 4346 12484 4402 12540
rect 4402 12484 4406 12540
rect 4342 12480 4406 12484
rect 7804 12540 7868 12544
rect 7804 12484 7808 12540
rect 7808 12484 7864 12540
rect 7864 12484 7868 12540
rect 7804 12480 7868 12484
rect 7884 12540 7948 12544
rect 7884 12484 7888 12540
rect 7888 12484 7944 12540
rect 7944 12484 7948 12540
rect 7884 12480 7948 12484
rect 7964 12540 8028 12544
rect 7964 12484 7968 12540
rect 7968 12484 8024 12540
rect 8024 12484 8028 12540
rect 7964 12480 8028 12484
rect 8044 12540 8108 12544
rect 8044 12484 8048 12540
rect 8048 12484 8104 12540
rect 8104 12484 8108 12540
rect 8044 12480 8108 12484
rect 11506 12540 11570 12544
rect 11506 12484 11510 12540
rect 11510 12484 11566 12540
rect 11566 12484 11570 12540
rect 11506 12480 11570 12484
rect 11586 12540 11650 12544
rect 11586 12484 11590 12540
rect 11590 12484 11646 12540
rect 11646 12484 11650 12540
rect 11586 12480 11650 12484
rect 11666 12540 11730 12544
rect 11666 12484 11670 12540
rect 11670 12484 11726 12540
rect 11726 12484 11730 12540
rect 11666 12480 11730 12484
rect 11746 12540 11810 12544
rect 11746 12484 11750 12540
rect 11750 12484 11806 12540
rect 11806 12484 11810 12540
rect 11746 12480 11810 12484
rect 15208 12540 15272 12544
rect 15208 12484 15212 12540
rect 15212 12484 15268 12540
rect 15268 12484 15272 12540
rect 15208 12480 15272 12484
rect 15288 12540 15352 12544
rect 15288 12484 15292 12540
rect 15292 12484 15348 12540
rect 15348 12484 15352 12540
rect 15288 12480 15352 12484
rect 15368 12540 15432 12544
rect 15368 12484 15372 12540
rect 15372 12484 15428 12540
rect 15428 12484 15432 12540
rect 15368 12480 15432 12484
rect 15448 12540 15512 12544
rect 15448 12484 15452 12540
rect 15452 12484 15508 12540
rect 15508 12484 15512 12540
rect 15448 12480 15512 12484
rect 2251 11996 2315 12000
rect 2251 11940 2255 11996
rect 2255 11940 2311 11996
rect 2311 11940 2315 11996
rect 2251 11936 2315 11940
rect 2331 11996 2395 12000
rect 2331 11940 2335 11996
rect 2335 11940 2391 11996
rect 2391 11940 2395 11996
rect 2331 11936 2395 11940
rect 2411 11996 2475 12000
rect 2411 11940 2415 11996
rect 2415 11940 2471 11996
rect 2471 11940 2475 11996
rect 2411 11936 2475 11940
rect 2491 11996 2555 12000
rect 2491 11940 2495 11996
rect 2495 11940 2551 11996
rect 2551 11940 2555 11996
rect 2491 11936 2555 11940
rect 5953 11996 6017 12000
rect 5953 11940 5957 11996
rect 5957 11940 6013 11996
rect 6013 11940 6017 11996
rect 5953 11936 6017 11940
rect 6033 11996 6097 12000
rect 6033 11940 6037 11996
rect 6037 11940 6093 11996
rect 6093 11940 6097 11996
rect 6033 11936 6097 11940
rect 6113 11996 6177 12000
rect 6113 11940 6117 11996
rect 6117 11940 6173 11996
rect 6173 11940 6177 11996
rect 6113 11936 6177 11940
rect 6193 11996 6257 12000
rect 6193 11940 6197 11996
rect 6197 11940 6253 11996
rect 6253 11940 6257 11996
rect 6193 11936 6257 11940
rect 9655 11996 9719 12000
rect 9655 11940 9659 11996
rect 9659 11940 9715 11996
rect 9715 11940 9719 11996
rect 9655 11936 9719 11940
rect 9735 11996 9799 12000
rect 9735 11940 9739 11996
rect 9739 11940 9795 11996
rect 9795 11940 9799 11996
rect 9735 11936 9799 11940
rect 9815 11996 9879 12000
rect 9815 11940 9819 11996
rect 9819 11940 9875 11996
rect 9875 11940 9879 11996
rect 9815 11936 9879 11940
rect 9895 11996 9959 12000
rect 9895 11940 9899 11996
rect 9899 11940 9955 11996
rect 9955 11940 9959 11996
rect 9895 11936 9959 11940
rect 13357 11996 13421 12000
rect 13357 11940 13361 11996
rect 13361 11940 13417 11996
rect 13417 11940 13421 11996
rect 13357 11936 13421 11940
rect 13437 11996 13501 12000
rect 13437 11940 13441 11996
rect 13441 11940 13497 11996
rect 13497 11940 13501 11996
rect 13437 11936 13501 11940
rect 13517 11996 13581 12000
rect 13517 11940 13521 11996
rect 13521 11940 13577 11996
rect 13577 11940 13581 11996
rect 13517 11936 13581 11940
rect 13597 11996 13661 12000
rect 13597 11940 13601 11996
rect 13601 11940 13657 11996
rect 13657 11940 13661 11996
rect 13597 11936 13661 11940
rect 4102 11452 4166 11456
rect 4102 11396 4106 11452
rect 4106 11396 4162 11452
rect 4162 11396 4166 11452
rect 4102 11392 4166 11396
rect 4182 11452 4246 11456
rect 4182 11396 4186 11452
rect 4186 11396 4242 11452
rect 4242 11396 4246 11452
rect 4182 11392 4246 11396
rect 4262 11452 4326 11456
rect 4262 11396 4266 11452
rect 4266 11396 4322 11452
rect 4322 11396 4326 11452
rect 4262 11392 4326 11396
rect 4342 11452 4406 11456
rect 4342 11396 4346 11452
rect 4346 11396 4402 11452
rect 4402 11396 4406 11452
rect 4342 11392 4406 11396
rect 7804 11452 7868 11456
rect 7804 11396 7808 11452
rect 7808 11396 7864 11452
rect 7864 11396 7868 11452
rect 7804 11392 7868 11396
rect 7884 11452 7948 11456
rect 7884 11396 7888 11452
rect 7888 11396 7944 11452
rect 7944 11396 7948 11452
rect 7884 11392 7948 11396
rect 7964 11452 8028 11456
rect 7964 11396 7968 11452
rect 7968 11396 8024 11452
rect 8024 11396 8028 11452
rect 7964 11392 8028 11396
rect 8044 11452 8108 11456
rect 8044 11396 8048 11452
rect 8048 11396 8104 11452
rect 8104 11396 8108 11452
rect 8044 11392 8108 11396
rect 11506 11452 11570 11456
rect 11506 11396 11510 11452
rect 11510 11396 11566 11452
rect 11566 11396 11570 11452
rect 11506 11392 11570 11396
rect 11586 11452 11650 11456
rect 11586 11396 11590 11452
rect 11590 11396 11646 11452
rect 11646 11396 11650 11452
rect 11586 11392 11650 11396
rect 11666 11452 11730 11456
rect 11666 11396 11670 11452
rect 11670 11396 11726 11452
rect 11726 11396 11730 11452
rect 11666 11392 11730 11396
rect 11746 11452 11810 11456
rect 11746 11396 11750 11452
rect 11750 11396 11806 11452
rect 11806 11396 11810 11452
rect 11746 11392 11810 11396
rect 15208 11452 15272 11456
rect 15208 11396 15212 11452
rect 15212 11396 15268 11452
rect 15268 11396 15272 11452
rect 15208 11392 15272 11396
rect 15288 11452 15352 11456
rect 15288 11396 15292 11452
rect 15292 11396 15348 11452
rect 15348 11396 15352 11452
rect 15288 11392 15352 11396
rect 15368 11452 15432 11456
rect 15368 11396 15372 11452
rect 15372 11396 15428 11452
rect 15428 11396 15432 11452
rect 15368 11392 15432 11396
rect 15448 11452 15512 11456
rect 15448 11396 15452 11452
rect 15452 11396 15508 11452
rect 15508 11396 15512 11452
rect 15448 11392 15512 11396
rect 2251 10908 2315 10912
rect 2251 10852 2255 10908
rect 2255 10852 2311 10908
rect 2311 10852 2315 10908
rect 2251 10848 2315 10852
rect 2331 10908 2395 10912
rect 2331 10852 2335 10908
rect 2335 10852 2391 10908
rect 2391 10852 2395 10908
rect 2331 10848 2395 10852
rect 2411 10908 2475 10912
rect 2411 10852 2415 10908
rect 2415 10852 2471 10908
rect 2471 10852 2475 10908
rect 2411 10848 2475 10852
rect 2491 10908 2555 10912
rect 2491 10852 2495 10908
rect 2495 10852 2551 10908
rect 2551 10852 2555 10908
rect 2491 10848 2555 10852
rect 5953 10908 6017 10912
rect 5953 10852 5957 10908
rect 5957 10852 6013 10908
rect 6013 10852 6017 10908
rect 5953 10848 6017 10852
rect 6033 10908 6097 10912
rect 6033 10852 6037 10908
rect 6037 10852 6093 10908
rect 6093 10852 6097 10908
rect 6033 10848 6097 10852
rect 6113 10908 6177 10912
rect 6113 10852 6117 10908
rect 6117 10852 6173 10908
rect 6173 10852 6177 10908
rect 6113 10848 6177 10852
rect 6193 10908 6257 10912
rect 6193 10852 6197 10908
rect 6197 10852 6253 10908
rect 6253 10852 6257 10908
rect 6193 10848 6257 10852
rect 9655 10908 9719 10912
rect 9655 10852 9659 10908
rect 9659 10852 9715 10908
rect 9715 10852 9719 10908
rect 9655 10848 9719 10852
rect 9735 10908 9799 10912
rect 9735 10852 9739 10908
rect 9739 10852 9795 10908
rect 9795 10852 9799 10908
rect 9735 10848 9799 10852
rect 9815 10908 9879 10912
rect 9815 10852 9819 10908
rect 9819 10852 9875 10908
rect 9875 10852 9879 10908
rect 9815 10848 9879 10852
rect 9895 10908 9959 10912
rect 9895 10852 9899 10908
rect 9899 10852 9955 10908
rect 9955 10852 9959 10908
rect 9895 10848 9959 10852
rect 13357 10908 13421 10912
rect 13357 10852 13361 10908
rect 13361 10852 13417 10908
rect 13417 10852 13421 10908
rect 13357 10848 13421 10852
rect 13437 10908 13501 10912
rect 13437 10852 13441 10908
rect 13441 10852 13497 10908
rect 13497 10852 13501 10908
rect 13437 10848 13501 10852
rect 13517 10908 13581 10912
rect 13517 10852 13521 10908
rect 13521 10852 13577 10908
rect 13577 10852 13581 10908
rect 13517 10848 13581 10852
rect 13597 10908 13661 10912
rect 13597 10852 13601 10908
rect 13601 10852 13657 10908
rect 13657 10852 13661 10908
rect 13597 10848 13661 10852
rect 4102 10364 4166 10368
rect 4102 10308 4106 10364
rect 4106 10308 4162 10364
rect 4162 10308 4166 10364
rect 4102 10304 4166 10308
rect 4182 10364 4246 10368
rect 4182 10308 4186 10364
rect 4186 10308 4242 10364
rect 4242 10308 4246 10364
rect 4182 10304 4246 10308
rect 4262 10364 4326 10368
rect 4262 10308 4266 10364
rect 4266 10308 4322 10364
rect 4322 10308 4326 10364
rect 4262 10304 4326 10308
rect 4342 10364 4406 10368
rect 4342 10308 4346 10364
rect 4346 10308 4402 10364
rect 4402 10308 4406 10364
rect 4342 10304 4406 10308
rect 7804 10364 7868 10368
rect 7804 10308 7808 10364
rect 7808 10308 7864 10364
rect 7864 10308 7868 10364
rect 7804 10304 7868 10308
rect 7884 10364 7948 10368
rect 7884 10308 7888 10364
rect 7888 10308 7944 10364
rect 7944 10308 7948 10364
rect 7884 10304 7948 10308
rect 7964 10364 8028 10368
rect 7964 10308 7968 10364
rect 7968 10308 8024 10364
rect 8024 10308 8028 10364
rect 7964 10304 8028 10308
rect 8044 10364 8108 10368
rect 8044 10308 8048 10364
rect 8048 10308 8104 10364
rect 8104 10308 8108 10364
rect 8044 10304 8108 10308
rect 11506 10364 11570 10368
rect 11506 10308 11510 10364
rect 11510 10308 11566 10364
rect 11566 10308 11570 10364
rect 11506 10304 11570 10308
rect 11586 10364 11650 10368
rect 11586 10308 11590 10364
rect 11590 10308 11646 10364
rect 11646 10308 11650 10364
rect 11586 10304 11650 10308
rect 11666 10364 11730 10368
rect 11666 10308 11670 10364
rect 11670 10308 11726 10364
rect 11726 10308 11730 10364
rect 11666 10304 11730 10308
rect 11746 10364 11810 10368
rect 11746 10308 11750 10364
rect 11750 10308 11806 10364
rect 11806 10308 11810 10364
rect 11746 10304 11810 10308
rect 15208 10364 15272 10368
rect 15208 10308 15212 10364
rect 15212 10308 15268 10364
rect 15268 10308 15272 10364
rect 15208 10304 15272 10308
rect 15288 10364 15352 10368
rect 15288 10308 15292 10364
rect 15292 10308 15348 10364
rect 15348 10308 15352 10364
rect 15288 10304 15352 10308
rect 15368 10364 15432 10368
rect 15368 10308 15372 10364
rect 15372 10308 15428 10364
rect 15428 10308 15432 10364
rect 15368 10304 15432 10308
rect 15448 10364 15512 10368
rect 15448 10308 15452 10364
rect 15452 10308 15508 10364
rect 15508 10308 15512 10364
rect 15448 10304 15512 10308
rect 2251 9820 2315 9824
rect 2251 9764 2255 9820
rect 2255 9764 2311 9820
rect 2311 9764 2315 9820
rect 2251 9760 2315 9764
rect 2331 9820 2395 9824
rect 2331 9764 2335 9820
rect 2335 9764 2391 9820
rect 2391 9764 2395 9820
rect 2331 9760 2395 9764
rect 2411 9820 2475 9824
rect 2411 9764 2415 9820
rect 2415 9764 2471 9820
rect 2471 9764 2475 9820
rect 2411 9760 2475 9764
rect 2491 9820 2555 9824
rect 2491 9764 2495 9820
rect 2495 9764 2551 9820
rect 2551 9764 2555 9820
rect 2491 9760 2555 9764
rect 5953 9820 6017 9824
rect 5953 9764 5957 9820
rect 5957 9764 6013 9820
rect 6013 9764 6017 9820
rect 5953 9760 6017 9764
rect 6033 9820 6097 9824
rect 6033 9764 6037 9820
rect 6037 9764 6093 9820
rect 6093 9764 6097 9820
rect 6033 9760 6097 9764
rect 6113 9820 6177 9824
rect 6113 9764 6117 9820
rect 6117 9764 6173 9820
rect 6173 9764 6177 9820
rect 6113 9760 6177 9764
rect 6193 9820 6257 9824
rect 6193 9764 6197 9820
rect 6197 9764 6253 9820
rect 6253 9764 6257 9820
rect 6193 9760 6257 9764
rect 9655 9820 9719 9824
rect 9655 9764 9659 9820
rect 9659 9764 9715 9820
rect 9715 9764 9719 9820
rect 9655 9760 9719 9764
rect 9735 9820 9799 9824
rect 9735 9764 9739 9820
rect 9739 9764 9795 9820
rect 9795 9764 9799 9820
rect 9735 9760 9799 9764
rect 9815 9820 9879 9824
rect 9815 9764 9819 9820
rect 9819 9764 9875 9820
rect 9875 9764 9879 9820
rect 9815 9760 9879 9764
rect 9895 9820 9959 9824
rect 9895 9764 9899 9820
rect 9899 9764 9955 9820
rect 9955 9764 9959 9820
rect 9895 9760 9959 9764
rect 13357 9820 13421 9824
rect 13357 9764 13361 9820
rect 13361 9764 13417 9820
rect 13417 9764 13421 9820
rect 13357 9760 13421 9764
rect 13437 9820 13501 9824
rect 13437 9764 13441 9820
rect 13441 9764 13497 9820
rect 13497 9764 13501 9820
rect 13437 9760 13501 9764
rect 13517 9820 13581 9824
rect 13517 9764 13521 9820
rect 13521 9764 13577 9820
rect 13577 9764 13581 9820
rect 13517 9760 13581 9764
rect 13597 9820 13661 9824
rect 13597 9764 13601 9820
rect 13601 9764 13657 9820
rect 13657 9764 13661 9820
rect 13597 9760 13661 9764
rect 4102 9276 4166 9280
rect 4102 9220 4106 9276
rect 4106 9220 4162 9276
rect 4162 9220 4166 9276
rect 4102 9216 4166 9220
rect 4182 9276 4246 9280
rect 4182 9220 4186 9276
rect 4186 9220 4242 9276
rect 4242 9220 4246 9276
rect 4182 9216 4246 9220
rect 4262 9276 4326 9280
rect 4262 9220 4266 9276
rect 4266 9220 4322 9276
rect 4322 9220 4326 9276
rect 4262 9216 4326 9220
rect 4342 9276 4406 9280
rect 4342 9220 4346 9276
rect 4346 9220 4402 9276
rect 4402 9220 4406 9276
rect 4342 9216 4406 9220
rect 7804 9276 7868 9280
rect 7804 9220 7808 9276
rect 7808 9220 7864 9276
rect 7864 9220 7868 9276
rect 7804 9216 7868 9220
rect 7884 9276 7948 9280
rect 7884 9220 7888 9276
rect 7888 9220 7944 9276
rect 7944 9220 7948 9276
rect 7884 9216 7948 9220
rect 7964 9276 8028 9280
rect 7964 9220 7968 9276
rect 7968 9220 8024 9276
rect 8024 9220 8028 9276
rect 7964 9216 8028 9220
rect 8044 9276 8108 9280
rect 8044 9220 8048 9276
rect 8048 9220 8104 9276
rect 8104 9220 8108 9276
rect 8044 9216 8108 9220
rect 11506 9276 11570 9280
rect 11506 9220 11510 9276
rect 11510 9220 11566 9276
rect 11566 9220 11570 9276
rect 11506 9216 11570 9220
rect 11586 9276 11650 9280
rect 11586 9220 11590 9276
rect 11590 9220 11646 9276
rect 11646 9220 11650 9276
rect 11586 9216 11650 9220
rect 11666 9276 11730 9280
rect 11666 9220 11670 9276
rect 11670 9220 11726 9276
rect 11726 9220 11730 9276
rect 11666 9216 11730 9220
rect 11746 9276 11810 9280
rect 11746 9220 11750 9276
rect 11750 9220 11806 9276
rect 11806 9220 11810 9276
rect 11746 9216 11810 9220
rect 15208 9276 15272 9280
rect 15208 9220 15212 9276
rect 15212 9220 15268 9276
rect 15268 9220 15272 9276
rect 15208 9216 15272 9220
rect 15288 9276 15352 9280
rect 15288 9220 15292 9276
rect 15292 9220 15348 9276
rect 15348 9220 15352 9276
rect 15288 9216 15352 9220
rect 15368 9276 15432 9280
rect 15368 9220 15372 9276
rect 15372 9220 15428 9276
rect 15428 9220 15432 9276
rect 15368 9216 15432 9220
rect 15448 9276 15512 9280
rect 15448 9220 15452 9276
rect 15452 9220 15508 9276
rect 15508 9220 15512 9276
rect 15448 9216 15512 9220
rect 2251 8732 2315 8736
rect 2251 8676 2255 8732
rect 2255 8676 2311 8732
rect 2311 8676 2315 8732
rect 2251 8672 2315 8676
rect 2331 8732 2395 8736
rect 2331 8676 2335 8732
rect 2335 8676 2391 8732
rect 2391 8676 2395 8732
rect 2331 8672 2395 8676
rect 2411 8732 2475 8736
rect 2411 8676 2415 8732
rect 2415 8676 2471 8732
rect 2471 8676 2475 8732
rect 2411 8672 2475 8676
rect 2491 8732 2555 8736
rect 2491 8676 2495 8732
rect 2495 8676 2551 8732
rect 2551 8676 2555 8732
rect 2491 8672 2555 8676
rect 5953 8732 6017 8736
rect 5953 8676 5957 8732
rect 5957 8676 6013 8732
rect 6013 8676 6017 8732
rect 5953 8672 6017 8676
rect 6033 8732 6097 8736
rect 6033 8676 6037 8732
rect 6037 8676 6093 8732
rect 6093 8676 6097 8732
rect 6033 8672 6097 8676
rect 6113 8732 6177 8736
rect 6113 8676 6117 8732
rect 6117 8676 6173 8732
rect 6173 8676 6177 8732
rect 6113 8672 6177 8676
rect 6193 8732 6257 8736
rect 6193 8676 6197 8732
rect 6197 8676 6253 8732
rect 6253 8676 6257 8732
rect 6193 8672 6257 8676
rect 9655 8732 9719 8736
rect 9655 8676 9659 8732
rect 9659 8676 9715 8732
rect 9715 8676 9719 8732
rect 9655 8672 9719 8676
rect 9735 8732 9799 8736
rect 9735 8676 9739 8732
rect 9739 8676 9795 8732
rect 9795 8676 9799 8732
rect 9735 8672 9799 8676
rect 9815 8732 9879 8736
rect 9815 8676 9819 8732
rect 9819 8676 9875 8732
rect 9875 8676 9879 8732
rect 9815 8672 9879 8676
rect 9895 8732 9959 8736
rect 9895 8676 9899 8732
rect 9899 8676 9955 8732
rect 9955 8676 9959 8732
rect 9895 8672 9959 8676
rect 13357 8732 13421 8736
rect 13357 8676 13361 8732
rect 13361 8676 13417 8732
rect 13417 8676 13421 8732
rect 13357 8672 13421 8676
rect 13437 8732 13501 8736
rect 13437 8676 13441 8732
rect 13441 8676 13497 8732
rect 13497 8676 13501 8732
rect 13437 8672 13501 8676
rect 13517 8732 13581 8736
rect 13517 8676 13521 8732
rect 13521 8676 13577 8732
rect 13577 8676 13581 8732
rect 13517 8672 13581 8676
rect 13597 8732 13661 8736
rect 13597 8676 13601 8732
rect 13601 8676 13657 8732
rect 13657 8676 13661 8732
rect 13597 8672 13661 8676
rect 4102 8188 4166 8192
rect 4102 8132 4106 8188
rect 4106 8132 4162 8188
rect 4162 8132 4166 8188
rect 4102 8128 4166 8132
rect 4182 8188 4246 8192
rect 4182 8132 4186 8188
rect 4186 8132 4242 8188
rect 4242 8132 4246 8188
rect 4182 8128 4246 8132
rect 4262 8188 4326 8192
rect 4262 8132 4266 8188
rect 4266 8132 4322 8188
rect 4322 8132 4326 8188
rect 4262 8128 4326 8132
rect 4342 8188 4406 8192
rect 4342 8132 4346 8188
rect 4346 8132 4402 8188
rect 4402 8132 4406 8188
rect 4342 8128 4406 8132
rect 7804 8188 7868 8192
rect 7804 8132 7808 8188
rect 7808 8132 7864 8188
rect 7864 8132 7868 8188
rect 7804 8128 7868 8132
rect 7884 8188 7948 8192
rect 7884 8132 7888 8188
rect 7888 8132 7944 8188
rect 7944 8132 7948 8188
rect 7884 8128 7948 8132
rect 7964 8188 8028 8192
rect 7964 8132 7968 8188
rect 7968 8132 8024 8188
rect 8024 8132 8028 8188
rect 7964 8128 8028 8132
rect 8044 8188 8108 8192
rect 8044 8132 8048 8188
rect 8048 8132 8104 8188
rect 8104 8132 8108 8188
rect 8044 8128 8108 8132
rect 11506 8188 11570 8192
rect 11506 8132 11510 8188
rect 11510 8132 11566 8188
rect 11566 8132 11570 8188
rect 11506 8128 11570 8132
rect 11586 8188 11650 8192
rect 11586 8132 11590 8188
rect 11590 8132 11646 8188
rect 11646 8132 11650 8188
rect 11586 8128 11650 8132
rect 11666 8188 11730 8192
rect 11666 8132 11670 8188
rect 11670 8132 11726 8188
rect 11726 8132 11730 8188
rect 11666 8128 11730 8132
rect 11746 8188 11810 8192
rect 11746 8132 11750 8188
rect 11750 8132 11806 8188
rect 11806 8132 11810 8188
rect 11746 8128 11810 8132
rect 15208 8188 15272 8192
rect 15208 8132 15212 8188
rect 15212 8132 15268 8188
rect 15268 8132 15272 8188
rect 15208 8128 15272 8132
rect 15288 8188 15352 8192
rect 15288 8132 15292 8188
rect 15292 8132 15348 8188
rect 15348 8132 15352 8188
rect 15288 8128 15352 8132
rect 15368 8188 15432 8192
rect 15368 8132 15372 8188
rect 15372 8132 15428 8188
rect 15428 8132 15432 8188
rect 15368 8128 15432 8132
rect 15448 8188 15512 8192
rect 15448 8132 15452 8188
rect 15452 8132 15508 8188
rect 15508 8132 15512 8188
rect 15448 8128 15512 8132
rect 2251 7644 2315 7648
rect 2251 7588 2255 7644
rect 2255 7588 2311 7644
rect 2311 7588 2315 7644
rect 2251 7584 2315 7588
rect 2331 7644 2395 7648
rect 2331 7588 2335 7644
rect 2335 7588 2391 7644
rect 2391 7588 2395 7644
rect 2331 7584 2395 7588
rect 2411 7644 2475 7648
rect 2411 7588 2415 7644
rect 2415 7588 2471 7644
rect 2471 7588 2475 7644
rect 2411 7584 2475 7588
rect 2491 7644 2555 7648
rect 2491 7588 2495 7644
rect 2495 7588 2551 7644
rect 2551 7588 2555 7644
rect 2491 7584 2555 7588
rect 5953 7644 6017 7648
rect 5953 7588 5957 7644
rect 5957 7588 6013 7644
rect 6013 7588 6017 7644
rect 5953 7584 6017 7588
rect 6033 7644 6097 7648
rect 6033 7588 6037 7644
rect 6037 7588 6093 7644
rect 6093 7588 6097 7644
rect 6033 7584 6097 7588
rect 6113 7644 6177 7648
rect 6113 7588 6117 7644
rect 6117 7588 6173 7644
rect 6173 7588 6177 7644
rect 6113 7584 6177 7588
rect 6193 7644 6257 7648
rect 6193 7588 6197 7644
rect 6197 7588 6253 7644
rect 6253 7588 6257 7644
rect 6193 7584 6257 7588
rect 9655 7644 9719 7648
rect 9655 7588 9659 7644
rect 9659 7588 9715 7644
rect 9715 7588 9719 7644
rect 9655 7584 9719 7588
rect 9735 7644 9799 7648
rect 9735 7588 9739 7644
rect 9739 7588 9795 7644
rect 9795 7588 9799 7644
rect 9735 7584 9799 7588
rect 9815 7644 9879 7648
rect 9815 7588 9819 7644
rect 9819 7588 9875 7644
rect 9875 7588 9879 7644
rect 9815 7584 9879 7588
rect 9895 7644 9959 7648
rect 9895 7588 9899 7644
rect 9899 7588 9955 7644
rect 9955 7588 9959 7644
rect 9895 7584 9959 7588
rect 13357 7644 13421 7648
rect 13357 7588 13361 7644
rect 13361 7588 13417 7644
rect 13417 7588 13421 7644
rect 13357 7584 13421 7588
rect 13437 7644 13501 7648
rect 13437 7588 13441 7644
rect 13441 7588 13497 7644
rect 13497 7588 13501 7644
rect 13437 7584 13501 7588
rect 13517 7644 13581 7648
rect 13517 7588 13521 7644
rect 13521 7588 13577 7644
rect 13577 7588 13581 7644
rect 13517 7584 13581 7588
rect 13597 7644 13661 7648
rect 13597 7588 13601 7644
rect 13601 7588 13657 7644
rect 13657 7588 13661 7644
rect 13597 7584 13661 7588
rect 4102 7100 4166 7104
rect 4102 7044 4106 7100
rect 4106 7044 4162 7100
rect 4162 7044 4166 7100
rect 4102 7040 4166 7044
rect 4182 7100 4246 7104
rect 4182 7044 4186 7100
rect 4186 7044 4242 7100
rect 4242 7044 4246 7100
rect 4182 7040 4246 7044
rect 4262 7100 4326 7104
rect 4262 7044 4266 7100
rect 4266 7044 4322 7100
rect 4322 7044 4326 7100
rect 4262 7040 4326 7044
rect 4342 7100 4406 7104
rect 4342 7044 4346 7100
rect 4346 7044 4402 7100
rect 4402 7044 4406 7100
rect 4342 7040 4406 7044
rect 7804 7100 7868 7104
rect 7804 7044 7808 7100
rect 7808 7044 7864 7100
rect 7864 7044 7868 7100
rect 7804 7040 7868 7044
rect 7884 7100 7948 7104
rect 7884 7044 7888 7100
rect 7888 7044 7944 7100
rect 7944 7044 7948 7100
rect 7884 7040 7948 7044
rect 7964 7100 8028 7104
rect 7964 7044 7968 7100
rect 7968 7044 8024 7100
rect 8024 7044 8028 7100
rect 7964 7040 8028 7044
rect 8044 7100 8108 7104
rect 8044 7044 8048 7100
rect 8048 7044 8104 7100
rect 8104 7044 8108 7100
rect 8044 7040 8108 7044
rect 11506 7100 11570 7104
rect 11506 7044 11510 7100
rect 11510 7044 11566 7100
rect 11566 7044 11570 7100
rect 11506 7040 11570 7044
rect 11586 7100 11650 7104
rect 11586 7044 11590 7100
rect 11590 7044 11646 7100
rect 11646 7044 11650 7100
rect 11586 7040 11650 7044
rect 11666 7100 11730 7104
rect 11666 7044 11670 7100
rect 11670 7044 11726 7100
rect 11726 7044 11730 7100
rect 11666 7040 11730 7044
rect 11746 7100 11810 7104
rect 11746 7044 11750 7100
rect 11750 7044 11806 7100
rect 11806 7044 11810 7100
rect 11746 7040 11810 7044
rect 15208 7100 15272 7104
rect 15208 7044 15212 7100
rect 15212 7044 15268 7100
rect 15268 7044 15272 7100
rect 15208 7040 15272 7044
rect 15288 7100 15352 7104
rect 15288 7044 15292 7100
rect 15292 7044 15348 7100
rect 15348 7044 15352 7100
rect 15288 7040 15352 7044
rect 15368 7100 15432 7104
rect 15368 7044 15372 7100
rect 15372 7044 15428 7100
rect 15428 7044 15432 7100
rect 15368 7040 15432 7044
rect 15448 7100 15512 7104
rect 15448 7044 15452 7100
rect 15452 7044 15508 7100
rect 15508 7044 15512 7100
rect 15448 7040 15512 7044
rect 2251 6556 2315 6560
rect 2251 6500 2255 6556
rect 2255 6500 2311 6556
rect 2311 6500 2315 6556
rect 2251 6496 2315 6500
rect 2331 6556 2395 6560
rect 2331 6500 2335 6556
rect 2335 6500 2391 6556
rect 2391 6500 2395 6556
rect 2331 6496 2395 6500
rect 2411 6556 2475 6560
rect 2411 6500 2415 6556
rect 2415 6500 2471 6556
rect 2471 6500 2475 6556
rect 2411 6496 2475 6500
rect 2491 6556 2555 6560
rect 2491 6500 2495 6556
rect 2495 6500 2551 6556
rect 2551 6500 2555 6556
rect 2491 6496 2555 6500
rect 5953 6556 6017 6560
rect 5953 6500 5957 6556
rect 5957 6500 6013 6556
rect 6013 6500 6017 6556
rect 5953 6496 6017 6500
rect 6033 6556 6097 6560
rect 6033 6500 6037 6556
rect 6037 6500 6093 6556
rect 6093 6500 6097 6556
rect 6033 6496 6097 6500
rect 6113 6556 6177 6560
rect 6113 6500 6117 6556
rect 6117 6500 6173 6556
rect 6173 6500 6177 6556
rect 6113 6496 6177 6500
rect 6193 6556 6257 6560
rect 6193 6500 6197 6556
rect 6197 6500 6253 6556
rect 6253 6500 6257 6556
rect 6193 6496 6257 6500
rect 9655 6556 9719 6560
rect 9655 6500 9659 6556
rect 9659 6500 9715 6556
rect 9715 6500 9719 6556
rect 9655 6496 9719 6500
rect 9735 6556 9799 6560
rect 9735 6500 9739 6556
rect 9739 6500 9795 6556
rect 9795 6500 9799 6556
rect 9735 6496 9799 6500
rect 9815 6556 9879 6560
rect 9815 6500 9819 6556
rect 9819 6500 9875 6556
rect 9875 6500 9879 6556
rect 9815 6496 9879 6500
rect 9895 6556 9959 6560
rect 9895 6500 9899 6556
rect 9899 6500 9955 6556
rect 9955 6500 9959 6556
rect 9895 6496 9959 6500
rect 13357 6556 13421 6560
rect 13357 6500 13361 6556
rect 13361 6500 13417 6556
rect 13417 6500 13421 6556
rect 13357 6496 13421 6500
rect 13437 6556 13501 6560
rect 13437 6500 13441 6556
rect 13441 6500 13497 6556
rect 13497 6500 13501 6556
rect 13437 6496 13501 6500
rect 13517 6556 13581 6560
rect 13517 6500 13521 6556
rect 13521 6500 13577 6556
rect 13577 6500 13581 6556
rect 13517 6496 13581 6500
rect 13597 6556 13661 6560
rect 13597 6500 13601 6556
rect 13601 6500 13657 6556
rect 13657 6500 13661 6556
rect 13597 6496 13661 6500
rect 4102 6012 4166 6016
rect 4102 5956 4106 6012
rect 4106 5956 4162 6012
rect 4162 5956 4166 6012
rect 4102 5952 4166 5956
rect 4182 6012 4246 6016
rect 4182 5956 4186 6012
rect 4186 5956 4242 6012
rect 4242 5956 4246 6012
rect 4182 5952 4246 5956
rect 4262 6012 4326 6016
rect 4262 5956 4266 6012
rect 4266 5956 4322 6012
rect 4322 5956 4326 6012
rect 4262 5952 4326 5956
rect 4342 6012 4406 6016
rect 4342 5956 4346 6012
rect 4346 5956 4402 6012
rect 4402 5956 4406 6012
rect 4342 5952 4406 5956
rect 7804 6012 7868 6016
rect 7804 5956 7808 6012
rect 7808 5956 7864 6012
rect 7864 5956 7868 6012
rect 7804 5952 7868 5956
rect 7884 6012 7948 6016
rect 7884 5956 7888 6012
rect 7888 5956 7944 6012
rect 7944 5956 7948 6012
rect 7884 5952 7948 5956
rect 7964 6012 8028 6016
rect 7964 5956 7968 6012
rect 7968 5956 8024 6012
rect 8024 5956 8028 6012
rect 7964 5952 8028 5956
rect 8044 6012 8108 6016
rect 8044 5956 8048 6012
rect 8048 5956 8104 6012
rect 8104 5956 8108 6012
rect 8044 5952 8108 5956
rect 11506 6012 11570 6016
rect 11506 5956 11510 6012
rect 11510 5956 11566 6012
rect 11566 5956 11570 6012
rect 11506 5952 11570 5956
rect 11586 6012 11650 6016
rect 11586 5956 11590 6012
rect 11590 5956 11646 6012
rect 11646 5956 11650 6012
rect 11586 5952 11650 5956
rect 11666 6012 11730 6016
rect 11666 5956 11670 6012
rect 11670 5956 11726 6012
rect 11726 5956 11730 6012
rect 11666 5952 11730 5956
rect 11746 6012 11810 6016
rect 11746 5956 11750 6012
rect 11750 5956 11806 6012
rect 11806 5956 11810 6012
rect 11746 5952 11810 5956
rect 15208 6012 15272 6016
rect 15208 5956 15212 6012
rect 15212 5956 15268 6012
rect 15268 5956 15272 6012
rect 15208 5952 15272 5956
rect 15288 6012 15352 6016
rect 15288 5956 15292 6012
rect 15292 5956 15348 6012
rect 15348 5956 15352 6012
rect 15288 5952 15352 5956
rect 15368 6012 15432 6016
rect 15368 5956 15372 6012
rect 15372 5956 15428 6012
rect 15428 5956 15432 6012
rect 15368 5952 15432 5956
rect 15448 6012 15512 6016
rect 15448 5956 15452 6012
rect 15452 5956 15508 6012
rect 15508 5956 15512 6012
rect 15448 5952 15512 5956
rect 2251 5468 2315 5472
rect 2251 5412 2255 5468
rect 2255 5412 2311 5468
rect 2311 5412 2315 5468
rect 2251 5408 2315 5412
rect 2331 5468 2395 5472
rect 2331 5412 2335 5468
rect 2335 5412 2391 5468
rect 2391 5412 2395 5468
rect 2331 5408 2395 5412
rect 2411 5468 2475 5472
rect 2411 5412 2415 5468
rect 2415 5412 2471 5468
rect 2471 5412 2475 5468
rect 2411 5408 2475 5412
rect 2491 5468 2555 5472
rect 2491 5412 2495 5468
rect 2495 5412 2551 5468
rect 2551 5412 2555 5468
rect 2491 5408 2555 5412
rect 5953 5468 6017 5472
rect 5953 5412 5957 5468
rect 5957 5412 6013 5468
rect 6013 5412 6017 5468
rect 5953 5408 6017 5412
rect 6033 5468 6097 5472
rect 6033 5412 6037 5468
rect 6037 5412 6093 5468
rect 6093 5412 6097 5468
rect 6033 5408 6097 5412
rect 6113 5468 6177 5472
rect 6113 5412 6117 5468
rect 6117 5412 6173 5468
rect 6173 5412 6177 5468
rect 6113 5408 6177 5412
rect 6193 5468 6257 5472
rect 6193 5412 6197 5468
rect 6197 5412 6253 5468
rect 6253 5412 6257 5468
rect 6193 5408 6257 5412
rect 9655 5468 9719 5472
rect 9655 5412 9659 5468
rect 9659 5412 9715 5468
rect 9715 5412 9719 5468
rect 9655 5408 9719 5412
rect 9735 5468 9799 5472
rect 9735 5412 9739 5468
rect 9739 5412 9795 5468
rect 9795 5412 9799 5468
rect 9735 5408 9799 5412
rect 9815 5468 9879 5472
rect 9815 5412 9819 5468
rect 9819 5412 9875 5468
rect 9875 5412 9879 5468
rect 9815 5408 9879 5412
rect 9895 5468 9959 5472
rect 9895 5412 9899 5468
rect 9899 5412 9955 5468
rect 9955 5412 9959 5468
rect 9895 5408 9959 5412
rect 13357 5468 13421 5472
rect 13357 5412 13361 5468
rect 13361 5412 13417 5468
rect 13417 5412 13421 5468
rect 13357 5408 13421 5412
rect 13437 5468 13501 5472
rect 13437 5412 13441 5468
rect 13441 5412 13497 5468
rect 13497 5412 13501 5468
rect 13437 5408 13501 5412
rect 13517 5468 13581 5472
rect 13517 5412 13521 5468
rect 13521 5412 13577 5468
rect 13577 5412 13581 5468
rect 13517 5408 13581 5412
rect 13597 5468 13661 5472
rect 13597 5412 13601 5468
rect 13601 5412 13657 5468
rect 13657 5412 13661 5468
rect 13597 5408 13661 5412
rect 4102 4924 4166 4928
rect 4102 4868 4106 4924
rect 4106 4868 4162 4924
rect 4162 4868 4166 4924
rect 4102 4864 4166 4868
rect 4182 4924 4246 4928
rect 4182 4868 4186 4924
rect 4186 4868 4242 4924
rect 4242 4868 4246 4924
rect 4182 4864 4246 4868
rect 4262 4924 4326 4928
rect 4262 4868 4266 4924
rect 4266 4868 4322 4924
rect 4322 4868 4326 4924
rect 4262 4864 4326 4868
rect 4342 4924 4406 4928
rect 4342 4868 4346 4924
rect 4346 4868 4402 4924
rect 4402 4868 4406 4924
rect 4342 4864 4406 4868
rect 7804 4924 7868 4928
rect 7804 4868 7808 4924
rect 7808 4868 7864 4924
rect 7864 4868 7868 4924
rect 7804 4864 7868 4868
rect 7884 4924 7948 4928
rect 7884 4868 7888 4924
rect 7888 4868 7944 4924
rect 7944 4868 7948 4924
rect 7884 4864 7948 4868
rect 7964 4924 8028 4928
rect 7964 4868 7968 4924
rect 7968 4868 8024 4924
rect 8024 4868 8028 4924
rect 7964 4864 8028 4868
rect 8044 4924 8108 4928
rect 8044 4868 8048 4924
rect 8048 4868 8104 4924
rect 8104 4868 8108 4924
rect 8044 4864 8108 4868
rect 11506 4924 11570 4928
rect 11506 4868 11510 4924
rect 11510 4868 11566 4924
rect 11566 4868 11570 4924
rect 11506 4864 11570 4868
rect 11586 4924 11650 4928
rect 11586 4868 11590 4924
rect 11590 4868 11646 4924
rect 11646 4868 11650 4924
rect 11586 4864 11650 4868
rect 11666 4924 11730 4928
rect 11666 4868 11670 4924
rect 11670 4868 11726 4924
rect 11726 4868 11730 4924
rect 11666 4864 11730 4868
rect 11746 4924 11810 4928
rect 11746 4868 11750 4924
rect 11750 4868 11806 4924
rect 11806 4868 11810 4924
rect 11746 4864 11810 4868
rect 15208 4924 15272 4928
rect 15208 4868 15212 4924
rect 15212 4868 15268 4924
rect 15268 4868 15272 4924
rect 15208 4864 15272 4868
rect 15288 4924 15352 4928
rect 15288 4868 15292 4924
rect 15292 4868 15348 4924
rect 15348 4868 15352 4924
rect 15288 4864 15352 4868
rect 15368 4924 15432 4928
rect 15368 4868 15372 4924
rect 15372 4868 15428 4924
rect 15428 4868 15432 4924
rect 15368 4864 15432 4868
rect 15448 4924 15512 4928
rect 15448 4868 15452 4924
rect 15452 4868 15508 4924
rect 15508 4868 15512 4924
rect 15448 4864 15512 4868
rect 2251 4380 2315 4384
rect 2251 4324 2255 4380
rect 2255 4324 2311 4380
rect 2311 4324 2315 4380
rect 2251 4320 2315 4324
rect 2331 4380 2395 4384
rect 2331 4324 2335 4380
rect 2335 4324 2391 4380
rect 2391 4324 2395 4380
rect 2331 4320 2395 4324
rect 2411 4380 2475 4384
rect 2411 4324 2415 4380
rect 2415 4324 2471 4380
rect 2471 4324 2475 4380
rect 2411 4320 2475 4324
rect 2491 4380 2555 4384
rect 2491 4324 2495 4380
rect 2495 4324 2551 4380
rect 2551 4324 2555 4380
rect 2491 4320 2555 4324
rect 5953 4380 6017 4384
rect 5953 4324 5957 4380
rect 5957 4324 6013 4380
rect 6013 4324 6017 4380
rect 5953 4320 6017 4324
rect 6033 4380 6097 4384
rect 6033 4324 6037 4380
rect 6037 4324 6093 4380
rect 6093 4324 6097 4380
rect 6033 4320 6097 4324
rect 6113 4380 6177 4384
rect 6113 4324 6117 4380
rect 6117 4324 6173 4380
rect 6173 4324 6177 4380
rect 6113 4320 6177 4324
rect 6193 4380 6257 4384
rect 6193 4324 6197 4380
rect 6197 4324 6253 4380
rect 6253 4324 6257 4380
rect 6193 4320 6257 4324
rect 9655 4380 9719 4384
rect 9655 4324 9659 4380
rect 9659 4324 9715 4380
rect 9715 4324 9719 4380
rect 9655 4320 9719 4324
rect 9735 4380 9799 4384
rect 9735 4324 9739 4380
rect 9739 4324 9795 4380
rect 9795 4324 9799 4380
rect 9735 4320 9799 4324
rect 9815 4380 9879 4384
rect 9815 4324 9819 4380
rect 9819 4324 9875 4380
rect 9875 4324 9879 4380
rect 9815 4320 9879 4324
rect 9895 4380 9959 4384
rect 9895 4324 9899 4380
rect 9899 4324 9955 4380
rect 9955 4324 9959 4380
rect 9895 4320 9959 4324
rect 13357 4380 13421 4384
rect 13357 4324 13361 4380
rect 13361 4324 13417 4380
rect 13417 4324 13421 4380
rect 13357 4320 13421 4324
rect 13437 4380 13501 4384
rect 13437 4324 13441 4380
rect 13441 4324 13497 4380
rect 13497 4324 13501 4380
rect 13437 4320 13501 4324
rect 13517 4380 13581 4384
rect 13517 4324 13521 4380
rect 13521 4324 13577 4380
rect 13577 4324 13581 4380
rect 13517 4320 13581 4324
rect 13597 4380 13661 4384
rect 13597 4324 13601 4380
rect 13601 4324 13657 4380
rect 13657 4324 13661 4380
rect 13597 4320 13661 4324
rect 4102 3836 4166 3840
rect 4102 3780 4106 3836
rect 4106 3780 4162 3836
rect 4162 3780 4166 3836
rect 4102 3776 4166 3780
rect 4182 3836 4246 3840
rect 4182 3780 4186 3836
rect 4186 3780 4242 3836
rect 4242 3780 4246 3836
rect 4182 3776 4246 3780
rect 4262 3836 4326 3840
rect 4262 3780 4266 3836
rect 4266 3780 4322 3836
rect 4322 3780 4326 3836
rect 4262 3776 4326 3780
rect 4342 3836 4406 3840
rect 4342 3780 4346 3836
rect 4346 3780 4402 3836
rect 4402 3780 4406 3836
rect 4342 3776 4406 3780
rect 7804 3836 7868 3840
rect 7804 3780 7808 3836
rect 7808 3780 7864 3836
rect 7864 3780 7868 3836
rect 7804 3776 7868 3780
rect 7884 3836 7948 3840
rect 7884 3780 7888 3836
rect 7888 3780 7944 3836
rect 7944 3780 7948 3836
rect 7884 3776 7948 3780
rect 7964 3836 8028 3840
rect 7964 3780 7968 3836
rect 7968 3780 8024 3836
rect 8024 3780 8028 3836
rect 7964 3776 8028 3780
rect 8044 3836 8108 3840
rect 8044 3780 8048 3836
rect 8048 3780 8104 3836
rect 8104 3780 8108 3836
rect 8044 3776 8108 3780
rect 11506 3836 11570 3840
rect 11506 3780 11510 3836
rect 11510 3780 11566 3836
rect 11566 3780 11570 3836
rect 11506 3776 11570 3780
rect 11586 3836 11650 3840
rect 11586 3780 11590 3836
rect 11590 3780 11646 3836
rect 11646 3780 11650 3836
rect 11586 3776 11650 3780
rect 11666 3836 11730 3840
rect 11666 3780 11670 3836
rect 11670 3780 11726 3836
rect 11726 3780 11730 3836
rect 11666 3776 11730 3780
rect 11746 3836 11810 3840
rect 11746 3780 11750 3836
rect 11750 3780 11806 3836
rect 11806 3780 11810 3836
rect 11746 3776 11810 3780
rect 15208 3836 15272 3840
rect 15208 3780 15212 3836
rect 15212 3780 15268 3836
rect 15268 3780 15272 3836
rect 15208 3776 15272 3780
rect 15288 3836 15352 3840
rect 15288 3780 15292 3836
rect 15292 3780 15348 3836
rect 15348 3780 15352 3836
rect 15288 3776 15352 3780
rect 15368 3836 15432 3840
rect 15368 3780 15372 3836
rect 15372 3780 15428 3836
rect 15428 3780 15432 3836
rect 15368 3776 15432 3780
rect 15448 3836 15512 3840
rect 15448 3780 15452 3836
rect 15452 3780 15508 3836
rect 15508 3780 15512 3836
rect 15448 3776 15512 3780
rect 2251 3292 2315 3296
rect 2251 3236 2255 3292
rect 2255 3236 2311 3292
rect 2311 3236 2315 3292
rect 2251 3232 2315 3236
rect 2331 3292 2395 3296
rect 2331 3236 2335 3292
rect 2335 3236 2391 3292
rect 2391 3236 2395 3292
rect 2331 3232 2395 3236
rect 2411 3292 2475 3296
rect 2411 3236 2415 3292
rect 2415 3236 2471 3292
rect 2471 3236 2475 3292
rect 2411 3232 2475 3236
rect 2491 3292 2555 3296
rect 2491 3236 2495 3292
rect 2495 3236 2551 3292
rect 2551 3236 2555 3292
rect 2491 3232 2555 3236
rect 5953 3292 6017 3296
rect 5953 3236 5957 3292
rect 5957 3236 6013 3292
rect 6013 3236 6017 3292
rect 5953 3232 6017 3236
rect 6033 3292 6097 3296
rect 6033 3236 6037 3292
rect 6037 3236 6093 3292
rect 6093 3236 6097 3292
rect 6033 3232 6097 3236
rect 6113 3292 6177 3296
rect 6113 3236 6117 3292
rect 6117 3236 6173 3292
rect 6173 3236 6177 3292
rect 6113 3232 6177 3236
rect 6193 3292 6257 3296
rect 6193 3236 6197 3292
rect 6197 3236 6253 3292
rect 6253 3236 6257 3292
rect 6193 3232 6257 3236
rect 9655 3292 9719 3296
rect 9655 3236 9659 3292
rect 9659 3236 9715 3292
rect 9715 3236 9719 3292
rect 9655 3232 9719 3236
rect 9735 3292 9799 3296
rect 9735 3236 9739 3292
rect 9739 3236 9795 3292
rect 9795 3236 9799 3292
rect 9735 3232 9799 3236
rect 9815 3292 9879 3296
rect 9815 3236 9819 3292
rect 9819 3236 9875 3292
rect 9875 3236 9879 3292
rect 9815 3232 9879 3236
rect 9895 3292 9959 3296
rect 9895 3236 9899 3292
rect 9899 3236 9955 3292
rect 9955 3236 9959 3292
rect 9895 3232 9959 3236
rect 13357 3292 13421 3296
rect 13357 3236 13361 3292
rect 13361 3236 13417 3292
rect 13417 3236 13421 3292
rect 13357 3232 13421 3236
rect 13437 3292 13501 3296
rect 13437 3236 13441 3292
rect 13441 3236 13497 3292
rect 13497 3236 13501 3292
rect 13437 3232 13501 3236
rect 13517 3292 13581 3296
rect 13517 3236 13521 3292
rect 13521 3236 13577 3292
rect 13577 3236 13581 3292
rect 13517 3232 13581 3236
rect 13597 3292 13661 3296
rect 13597 3236 13601 3292
rect 13601 3236 13657 3292
rect 13657 3236 13661 3292
rect 13597 3232 13661 3236
rect 4102 2748 4166 2752
rect 4102 2692 4106 2748
rect 4106 2692 4162 2748
rect 4162 2692 4166 2748
rect 4102 2688 4166 2692
rect 4182 2748 4246 2752
rect 4182 2692 4186 2748
rect 4186 2692 4242 2748
rect 4242 2692 4246 2748
rect 4182 2688 4246 2692
rect 4262 2748 4326 2752
rect 4262 2692 4266 2748
rect 4266 2692 4322 2748
rect 4322 2692 4326 2748
rect 4262 2688 4326 2692
rect 4342 2748 4406 2752
rect 4342 2692 4346 2748
rect 4346 2692 4402 2748
rect 4402 2692 4406 2748
rect 4342 2688 4406 2692
rect 7804 2748 7868 2752
rect 7804 2692 7808 2748
rect 7808 2692 7864 2748
rect 7864 2692 7868 2748
rect 7804 2688 7868 2692
rect 7884 2748 7948 2752
rect 7884 2692 7888 2748
rect 7888 2692 7944 2748
rect 7944 2692 7948 2748
rect 7884 2688 7948 2692
rect 7964 2748 8028 2752
rect 7964 2692 7968 2748
rect 7968 2692 8024 2748
rect 8024 2692 8028 2748
rect 7964 2688 8028 2692
rect 8044 2748 8108 2752
rect 8044 2692 8048 2748
rect 8048 2692 8104 2748
rect 8104 2692 8108 2748
rect 8044 2688 8108 2692
rect 11506 2748 11570 2752
rect 11506 2692 11510 2748
rect 11510 2692 11566 2748
rect 11566 2692 11570 2748
rect 11506 2688 11570 2692
rect 11586 2748 11650 2752
rect 11586 2692 11590 2748
rect 11590 2692 11646 2748
rect 11646 2692 11650 2748
rect 11586 2688 11650 2692
rect 11666 2748 11730 2752
rect 11666 2692 11670 2748
rect 11670 2692 11726 2748
rect 11726 2692 11730 2748
rect 11666 2688 11730 2692
rect 11746 2748 11810 2752
rect 11746 2692 11750 2748
rect 11750 2692 11806 2748
rect 11806 2692 11810 2748
rect 11746 2688 11810 2692
rect 15208 2748 15272 2752
rect 15208 2692 15212 2748
rect 15212 2692 15268 2748
rect 15268 2692 15272 2748
rect 15208 2688 15272 2692
rect 15288 2748 15352 2752
rect 15288 2692 15292 2748
rect 15292 2692 15348 2748
rect 15348 2692 15352 2748
rect 15288 2688 15352 2692
rect 15368 2748 15432 2752
rect 15368 2692 15372 2748
rect 15372 2692 15428 2748
rect 15428 2692 15432 2748
rect 15368 2688 15432 2692
rect 15448 2748 15512 2752
rect 15448 2692 15452 2748
rect 15452 2692 15508 2748
rect 15508 2692 15512 2748
rect 15448 2688 15512 2692
rect 2251 2204 2315 2208
rect 2251 2148 2255 2204
rect 2255 2148 2311 2204
rect 2311 2148 2315 2204
rect 2251 2144 2315 2148
rect 2331 2204 2395 2208
rect 2331 2148 2335 2204
rect 2335 2148 2391 2204
rect 2391 2148 2395 2204
rect 2331 2144 2395 2148
rect 2411 2204 2475 2208
rect 2411 2148 2415 2204
rect 2415 2148 2471 2204
rect 2471 2148 2475 2204
rect 2411 2144 2475 2148
rect 2491 2204 2555 2208
rect 2491 2148 2495 2204
rect 2495 2148 2551 2204
rect 2551 2148 2555 2204
rect 2491 2144 2555 2148
rect 5953 2204 6017 2208
rect 5953 2148 5957 2204
rect 5957 2148 6013 2204
rect 6013 2148 6017 2204
rect 5953 2144 6017 2148
rect 6033 2204 6097 2208
rect 6033 2148 6037 2204
rect 6037 2148 6093 2204
rect 6093 2148 6097 2204
rect 6033 2144 6097 2148
rect 6113 2204 6177 2208
rect 6113 2148 6117 2204
rect 6117 2148 6173 2204
rect 6173 2148 6177 2204
rect 6113 2144 6177 2148
rect 6193 2204 6257 2208
rect 6193 2148 6197 2204
rect 6197 2148 6253 2204
rect 6253 2148 6257 2204
rect 6193 2144 6257 2148
rect 9655 2204 9719 2208
rect 9655 2148 9659 2204
rect 9659 2148 9715 2204
rect 9715 2148 9719 2204
rect 9655 2144 9719 2148
rect 9735 2204 9799 2208
rect 9735 2148 9739 2204
rect 9739 2148 9795 2204
rect 9795 2148 9799 2204
rect 9735 2144 9799 2148
rect 9815 2204 9879 2208
rect 9815 2148 9819 2204
rect 9819 2148 9875 2204
rect 9875 2148 9879 2204
rect 9815 2144 9879 2148
rect 9895 2204 9959 2208
rect 9895 2148 9899 2204
rect 9899 2148 9955 2204
rect 9955 2148 9959 2204
rect 9895 2144 9959 2148
rect 13357 2204 13421 2208
rect 13357 2148 13361 2204
rect 13361 2148 13417 2204
rect 13417 2148 13421 2204
rect 13357 2144 13421 2148
rect 13437 2204 13501 2208
rect 13437 2148 13441 2204
rect 13441 2148 13497 2204
rect 13497 2148 13501 2204
rect 13437 2144 13501 2148
rect 13517 2204 13581 2208
rect 13517 2148 13521 2204
rect 13521 2148 13577 2204
rect 13577 2148 13581 2204
rect 13517 2144 13581 2148
rect 13597 2204 13661 2208
rect 13597 2148 13601 2204
rect 13601 2148 13657 2204
rect 13657 2148 13661 2204
rect 13597 2144 13661 2148
rect 4102 1660 4166 1664
rect 4102 1604 4106 1660
rect 4106 1604 4162 1660
rect 4162 1604 4166 1660
rect 4102 1600 4166 1604
rect 4182 1660 4246 1664
rect 4182 1604 4186 1660
rect 4186 1604 4242 1660
rect 4242 1604 4246 1660
rect 4182 1600 4246 1604
rect 4262 1660 4326 1664
rect 4262 1604 4266 1660
rect 4266 1604 4322 1660
rect 4322 1604 4326 1660
rect 4262 1600 4326 1604
rect 4342 1660 4406 1664
rect 4342 1604 4346 1660
rect 4346 1604 4402 1660
rect 4402 1604 4406 1660
rect 4342 1600 4406 1604
rect 7804 1660 7868 1664
rect 7804 1604 7808 1660
rect 7808 1604 7864 1660
rect 7864 1604 7868 1660
rect 7804 1600 7868 1604
rect 7884 1660 7948 1664
rect 7884 1604 7888 1660
rect 7888 1604 7944 1660
rect 7944 1604 7948 1660
rect 7884 1600 7948 1604
rect 7964 1660 8028 1664
rect 7964 1604 7968 1660
rect 7968 1604 8024 1660
rect 8024 1604 8028 1660
rect 7964 1600 8028 1604
rect 8044 1660 8108 1664
rect 8044 1604 8048 1660
rect 8048 1604 8104 1660
rect 8104 1604 8108 1660
rect 8044 1600 8108 1604
rect 11506 1660 11570 1664
rect 11506 1604 11510 1660
rect 11510 1604 11566 1660
rect 11566 1604 11570 1660
rect 11506 1600 11570 1604
rect 11586 1660 11650 1664
rect 11586 1604 11590 1660
rect 11590 1604 11646 1660
rect 11646 1604 11650 1660
rect 11586 1600 11650 1604
rect 11666 1660 11730 1664
rect 11666 1604 11670 1660
rect 11670 1604 11726 1660
rect 11726 1604 11730 1660
rect 11666 1600 11730 1604
rect 11746 1660 11810 1664
rect 11746 1604 11750 1660
rect 11750 1604 11806 1660
rect 11806 1604 11810 1660
rect 11746 1600 11810 1604
rect 15208 1660 15272 1664
rect 15208 1604 15212 1660
rect 15212 1604 15268 1660
rect 15268 1604 15272 1660
rect 15208 1600 15272 1604
rect 15288 1660 15352 1664
rect 15288 1604 15292 1660
rect 15292 1604 15348 1660
rect 15348 1604 15352 1660
rect 15288 1600 15352 1604
rect 15368 1660 15432 1664
rect 15368 1604 15372 1660
rect 15372 1604 15428 1660
rect 15428 1604 15432 1660
rect 15368 1600 15432 1604
rect 15448 1660 15512 1664
rect 15448 1604 15452 1660
rect 15452 1604 15508 1660
rect 15508 1604 15512 1660
rect 15448 1600 15512 1604
rect 2251 1116 2315 1120
rect 2251 1060 2255 1116
rect 2255 1060 2311 1116
rect 2311 1060 2315 1116
rect 2251 1056 2315 1060
rect 2331 1116 2395 1120
rect 2331 1060 2335 1116
rect 2335 1060 2391 1116
rect 2391 1060 2395 1116
rect 2331 1056 2395 1060
rect 2411 1116 2475 1120
rect 2411 1060 2415 1116
rect 2415 1060 2471 1116
rect 2471 1060 2475 1116
rect 2411 1056 2475 1060
rect 2491 1116 2555 1120
rect 2491 1060 2495 1116
rect 2495 1060 2551 1116
rect 2551 1060 2555 1116
rect 2491 1056 2555 1060
rect 5953 1116 6017 1120
rect 5953 1060 5957 1116
rect 5957 1060 6013 1116
rect 6013 1060 6017 1116
rect 5953 1056 6017 1060
rect 6033 1116 6097 1120
rect 6033 1060 6037 1116
rect 6037 1060 6093 1116
rect 6093 1060 6097 1116
rect 6033 1056 6097 1060
rect 6113 1116 6177 1120
rect 6113 1060 6117 1116
rect 6117 1060 6173 1116
rect 6173 1060 6177 1116
rect 6113 1056 6177 1060
rect 6193 1116 6257 1120
rect 6193 1060 6197 1116
rect 6197 1060 6253 1116
rect 6253 1060 6257 1116
rect 6193 1056 6257 1060
rect 9655 1116 9719 1120
rect 9655 1060 9659 1116
rect 9659 1060 9715 1116
rect 9715 1060 9719 1116
rect 9655 1056 9719 1060
rect 9735 1116 9799 1120
rect 9735 1060 9739 1116
rect 9739 1060 9795 1116
rect 9795 1060 9799 1116
rect 9735 1056 9799 1060
rect 9815 1116 9879 1120
rect 9815 1060 9819 1116
rect 9819 1060 9875 1116
rect 9875 1060 9879 1116
rect 9815 1056 9879 1060
rect 9895 1116 9959 1120
rect 9895 1060 9899 1116
rect 9899 1060 9955 1116
rect 9955 1060 9959 1116
rect 9895 1056 9959 1060
rect 13357 1116 13421 1120
rect 13357 1060 13361 1116
rect 13361 1060 13417 1116
rect 13417 1060 13421 1116
rect 13357 1056 13421 1060
rect 13437 1116 13501 1120
rect 13437 1060 13441 1116
rect 13441 1060 13497 1116
rect 13497 1060 13501 1116
rect 13437 1056 13501 1060
rect 13517 1116 13581 1120
rect 13517 1060 13521 1116
rect 13521 1060 13577 1116
rect 13577 1060 13581 1116
rect 13517 1056 13581 1060
rect 13597 1116 13661 1120
rect 13597 1060 13601 1116
rect 13601 1060 13657 1116
rect 13657 1060 13661 1116
rect 13597 1056 13661 1060
rect 4102 572 4166 576
rect 4102 516 4106 572
rect 4106 516 4162 572
rect 4162 516 4166 572
rect 4102 512 4166 516
rect 4182 572 4246 576
rect 4182 516 4186 572
rect 4186 516 4242 572
rect 4242 516 4246 572
rect 4182 512 4246 516
rect 4262 572 4326 576
rect 4262 516 4266 572
rect 4266 516 4322 572
rect 4322 516 4326 572
rect 4262 512 4326 516
rect 4342 572 4406 576
rect 4342 516 4346 572
rect 4346 516 4402 572
rect 4402 516 4406 572
rect 4342 512 4406 516
rect 7804 572 7868 576
rect 7804 516 7808 572
rect 7808 516 7864 572
rect 7864 516 7868 572
rect 7804 512 7868 516
rect 7884 572 7948 576
rect 7884 516 7888 572
rect 7888 516 7944 572
rect 7944 516 7948 572
rect 7884 512 7948 516
rect 7964 572 8028 576
rect 7964 516 7968 572
rect 7968 516 8024 572
rect 8024 516 8028 572
rect 7964 512 8028 516
rect 8044 572 8108 576
rect 8044 516 8048 572
rect 8048 516 8104 572
rect 8104 516 8108 572
rect 8044 512 8108 516
rect 11506 572 11570 576
rect 11506 516 11510 572
rect 11510 516 11566 572
rect 11566 516 11570 572
rect 11506 512 11570 516
rect 11586 572 11650 576
rect 11586 516 11590 572
rect 11590 516 11646 572
rect 11646 516 11650 572
rect 11586 512 11650 516
rect 11666 572 11730 576
rect 11666 516 11670 572
rect 11670 516 11726 572
rect 11726 516 11730 572
rect 11666 512 11730 516
rect 11746 572 11810 576
rect 11746 516 11750 572
rect 11750 516 11806 572
rect 11806 516 11810 572
rect 11746 512 11810 516
rect 15208 572 15272 576
rect 15208 516 15212 572
rect 15212 516 15268 572
rect 15268 516 15272 572
rect 15208 512 15272 516
rect 15288 572 15352 576
rect 15288 516 15292 572
rect 15292 516 15348 572
rect 15348 516 15352 572
rect 15288 512 15352 516
rect 15368 572 15432 576
rect 15368 516 15372 572
rect 15372 516 15428 572
rect 15428 516 15432 572
rect 15368 512 15432 516
rect 15448 572 15512 576
rect 15448 516 15452 572
rect 15452 516 15508 572
rect 15508 516 15512 572
rect 15448 512 15512 516
<< metal4 >>
rect 2243 15264 2563 15280
rect 2243 15200 2251 15264
rect 2315 15200 2331 15264
rect 2395 15200 2411 15264
rect 2475 15200 2491 15264
rect 2555 15200 2563 15264
rect 2243 14176 2563 15200
rect 2243 14112 2251 14176
rect 2315 14112 2331 14176
rect 2395 14112 2411 14176
rect 2475 14112 2491 14176
rect 2555 14112 2563 14176
rect 2243 13088 2563 14112
rect 2243 13024 2251 13088
rect 2315 13024 2331 13088
rect 2395 13024 2411 13088
rect 2475 13024 2491 13088
rect 2555 13024 2563 13088
rect 2243 12000 2563 13024
rect 2243 11936 2251 12000
rect 2315 11936 2331 12000
rect 2395 11936 2411 12000
rect 2475 11936 2491 12000
rect 2555 11936 2563 12000
rect 2243 10912 2563 11936
rect 2243 10848 2251 10912
rect 2315 10848 2331 10912
rect 2395 10848 2411 10912
rect 2475 10848 2491 10912
rect 2555 10848 2563 10912
rect 2243 9824 2563 10848
rect 2243 9760 2251 9824
rect 2315 9760 2331 9824
rect 2395 9760 2411 9824
rect 2475 9760 2491 9824
rect 2555 9760 2563 9824
rect 2243 8736 2563 9760
rect 2243 8672 2251 8736
rect 2315 8672 2331 8736
rect 2395 8672 2411 8736
rect 2475 8672 2491 8736
rect 2555 8672 2563 8736
rect 2243 7648 2563 8672
rect 2243 7584 2251 7648
rect 2315 7584 2331 7648
rect 2395 7584 2411 7648
rect 2475 7584 2491 7648
rect 2555 7584 2563 7648
rect 2243 6560 2563 7584
rect 2243 6496 2251 6560
rect 2315 6496 2331 6560
rect 2395 6496 2411 6560
rect 2475 6496 2491 6560
rect 2555 6496 2563 6560
rect 2243 5472 2563 6496
rect 2243 5408 2251 5472
rect 2315 5408 2331 5472
rect 2395 5408 2411 5472
rect 2475 5408 2491 5472
rect 2555 5408 2563 5472
rect 2243 4384 2563 5408
rect 2243 4320 2251 4384
rect 2315 4320 2331 4384
rect 2395 4320 2411 4384
rect 2475 4320 2491 4384
rect 2555 4320 2563 4384
rect 2243 3296 2563 4320
rect 2243 3232 2251 3296
rect 2315 3232 2331 3296
rect 2395 3232 2411 3296
rect 2475 3232 2491 3296
rect 2555 3232 2563 3296
rect 2243 2208 2563 3232
rect 2243 2144 2251 2208
rect 2315 2144 2331 2208
rect 2395 2144 2411 2208
rect 2475 2144 2491 2208
rect 2555 2144 2563 2208
rect 2243 1120 2563 2144
rect 2243 1056 2251 1120
rect 2315 1056 2331 1120
rect 2395 1056 2411 1120
rect 2475 1056 2491 1120
rect 2555 1056 2563 1120
rect 2243 496 2563 1056
rect 4094 14720 4414 15280
rect 4094 14656 4102 14720
rect 4166 14656 4182 14720
rect 4246 14656 4262 14720
rect 4326 14656 4342 14720
rect 4406 14656 4414 14720
rect 4094 13632 4414 14656
rect 4094 13568 4102 13632
rect 4166 13568 4182 13632
rect 4246 13568 4262 13632
rect 4326 13568 4342 13632
rect 4406 13568 4414 13632
rect 4094 12544 4414 13568
rect 4094 12480 4102 12544
rect 4166 12480 4182 12544
rect 4246 12480 4262 12544
rect 4326 12480 4342 12544
rect 4406 12480 4414 12544
rect 4094 11456 4414 12480
rect 4094 11392 4102 11456
rect 4166 11392 4182 11456
rect 4246 11392 4262 11456
rect 4326 11392 4342 11456
rect 4406 11392 4414 11456
rect 4094 10368 4414 11392
rect 4094 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4342 10368
rect 4406 10304 4414 10368
rect 4094 9280 4414 10304
rect 4094 9216 4102 9280
rect 4166 9216 4182 9280
rect 4246 9216 4262 9280
rect 4326 9216 4342 9280
rect 4406 9216 4414 9280
rect 4094 8192 4414 9216
rect 4094 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4342 8192
rect 4406 8128 4414 8192
rect 4094 7104 4414 8128
rect 4094 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4342 7104
rect 4406 7040 4414 7104
rect 4094 6016 4414 7040
rect 4094 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4342 6016
rect 4406 5952 4414 6016
rect 4094 4928 4414 5952
rect 4094 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4342 4928
rect 4406 4864 4414 4928
rect 4094 3840 4414 4864
rect 4094 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4342 3840
rect 4406 3776 4414 3840
rect 4094 2752 4414 3776
rect 4094 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4342 2752
rect 4406 2688 4414 2752
rect 4094 1664 4414 2688
rect 4094 1600 4102 1664
rect 4166 1600 4182 1664
rect 4246 1600 4262 1664
rect 4326 1600 4342 1664
rect 4406 1600 4414 1664
rect 4094 576 4414 1600
rect 4094 512 4102 576
rect 4166 512 4182 576
rect 4246 512 4262 576
rect 4326 512 4342 576
rect 4406 512 4414 576
rect 4094 496 4414 512
rect 5945 15264 6265 15280
rect 5945 15200 5953 15264
rect 6017 15200 6033 15264
rect 6097 15200 6113 15264
rect 6177 15200 6193 15264
rect 6257 15200 6265 15264
rect 5945 14176 6265 15200
rect 5945 14112 5953 14176
rect 6017 14112 6033 14176
rect 6097 14112 6113 14176
rect 6177 14112 6193 14176
rect 6257 14112 6265 14176
rect 5945 13088 6265 14112
rect 5945 13024 5953 13088
rect 6017 13024 6033 13088
rect 6097 13024 6113 13088
rect 6177 13024 6193 13088
rect 6257 13024 6265 13088
rect 5945 12000 6265 13024
rect 5945 11936 5953 12000
rect 6017 11936 6033 12000
rect 6097 11936 6113 12000
rect 6177 11936 6193 12000
rect 6257 11936 6265 12000
rect 5945 10912 6265 11936
rect 5945 10848 5953 10912
rect 6017 10848 6033 10912
rect 6097 10848 6113 10912
rect 6177 10848 6193 10912
rect 6257 10848 6265 10912
rect 5945 9824 6265 10848
rect 5945 9760 5953 9824
rect 6017 9760 6033 9824
rect 6097 9760 6113 9824
rect 6177 9760 6193 9824
rect 6257 9760 6265 9824
rect 5945 8736 6265 9760
rect 5945 8672 5953 8736
rect 6017 8672 6033 8736
rect 6097 8672 6113 8736
rect 6177 8672 6193 8736
rect 6257 8672 6265 8736
rect 5945 7648 6265 8672
rect 5945 7584 5953 7648
rect 6017 7584 6033 7648
rect 6097 7584 6113 7648
rect 6177 7584 6193 7648
rect 6257 7584 6265 7648
rect 5945 6560 6265 7584
rect 5945 6496 5953 6560
rect 6017 6496 6033 6560
rect 6097 6496 6113 6560
rect 6177 6496 6193 6560
rect 6257 6496 6265 6560
rect 5945 5472 6265 6496
rect 5945 5408 5953 5472
rect 6017 5408 6033 5472
rect 6097 5408 6113 5472
rect 6177 5408 6193 5472
rect 6257 5408 6265 5472
rect 5945 4384 6265 5408
rect 5945 4320 5953 4384
rect 6017 4320 6033 4384
rect 6097 4320 6113 4384
rect 6177 4320 6193 4384
rect 6257 4320 6265 4384
rect 5945 3296 6265 4320
rect 5945 3232 5953 3296
rect 6017 3232 6033 3296
rect 6097 3232 6113 3296
rect 6177 3232 6193 3296
rect 6257 3232 6265 3296
rect 5945 2208 6265 3232
rect 5945 2144 5953 2208
rect 6017 2144 6033 2208
rect 6097 2144 6113 2208
rect 6177 2144 6193 2208
rect 6257 2144 6265 2208
rect 5945 1120 6265 2144
rect 5945 1056 5953 1120
rect 6017 1056 6033 1120
rect 6097 1056 6113 1120
rect 6177 1056 6193 1120
rect 6257 1056 6265 1120
rect 5945 496 6265 1056
rect 7796 14720 8116 15280
rect 7796 14656 7804 14720
rect 7868 14656 7884 14720
rect 7948 14656 7964 14720
rect 8028 14656 8044 14720
rect 8108 14656 8116 14720
rect 7796 13632 8116 14656
rect 7796 13568 7804 13632
rect 7868 13568 7884 13632
rect 7948 13568 7964 13632
rect 8028 13568 8044 13632
rect 8108 13568 8116 13632
rect 7796 12544 8116 13568
rect 7796 12480 7804 12544
rect 7868 12480 7884 12544
rect 7948 12480 7964 12544
rect 8028 12480 8044 12544
rect 8108 12480 8116 12544
rect 7796 11456 8116 12480
rect 7796 11392 7804 11456
rect 7868 11392 7884 11456
rect 7948 11392 7964 11456
rect 8028 11392 8044 11456
rect 8108 11392 8116 11456
rect 7796 10368 8116 11392
rect 7796 10304 7804 10368
rect 7868 10304 7884 10368
rect 7948 10304 7964 10368
rect 8028 10304 8044 10368
rect 8108 10304 8116 10368
rect 7796 9280 8116 10304
rect 7796 9216 7804 9280
rect 7868 9216 7884 9280
rect 7948 9216 7964 9280
rect 8028 9216 8044 9280
rect 8108 9216 8116 9280
rect 7796 8192 8116 9216
rect 7796 8128 7804 8192
rect 7868 8128 7884 8192
rect 7948 8128 7964 8192
rect 8028 8128 8044 8192
rect 8108 8128 8116 8192
rect 7796 7104 8116 8128
rect 7796 7040 7804 7104
rect 7868 7040 7884 7104
rect 7948 7040 7964 7104
rect 8028 7040 8044 7104
rect 8108 7040 8116 7104
rect 7796 6016 8116 7040
rect 7796 5952 7804 6016
rect 7868 5952 7884 6016
rect 7948 5952 7964 6016
rect 8028 5952 8044 6016
rect 8108 5952 8116 6016
rect 7796 4928 8116 5952
rect 7796 4864 7804 4928
rect 7868 4864 7884 4928
rect 7948 4864 7964 4928
rect 8028 4864 8044 4928
rect 8108 4864 8116 4928
rect 7796 3840 8116 4864
rect 7796 3776 7804 3840
rect 7868 3776 7884 3840
rect 7948 3776 7964 3840
rect 8028 3776 8044 3840
rect 8108 3776 8116 3840
rect 7796 2752 8116 3776
rect 7796 2688 7804 2752
rect 7868 2688 7884 2752
rect 7948 2688 7964 2752
rect 8028 2688 8044 2752
rect 8108 2688 8116 2752
rect 7796 1664 8116 2688
rect 7796 1600 7804 1664
rect 7868 1600 7884 1664
rect 7948 1600 7964 1664
rect 8028 1600 8044 1664
rect 8108 1600 8116 1664
rect 7796 576 8116 1600
rect 7796 512 7804 576
rect 7868 512 7884 576
rect 7948 512 7964 576
rect 8028 512 8044 576
rect 8108 512 8116 576
rect 7796 496 8116 512
rect 9647 15264 9967 15280
rect 9647 15200 9655 15264
rect 9719 15200 9735 15264
rect 9799 15200 9815 15264
rect 9879 15200 9895 15264
rect 9959 15200 9967 15264
rect 9647 14176 9967 15200
rect 9647 14112 9655 14176
rect 9719 14112 9735 14176
rect 9799 14112 9815 14176
rect 9879 14112 9895 14176
rect 9959 14112 9967 14176
rect 9647 13088 9967 14112
rect 9647 13024 9655 13088
rect 9719 13024 9735 13088
rect 9799 13024 9815 13088
rect 9879 13024 9895 13088
rect 9959 13024 9967 13088
rect 9647 12000 9967 13024
rect 9647 11936 9655 12000
rect 9719 11936 9735 12000
rect 9799 11936 9815 12000
rect 9879 11936 9895 12000
rect 9959 11936 9967 12000
rect 9647 10912 9967 11936
rect 9647 10848 9655 10912
rect 9719 10848 9735 10912
rect 9799 10848 9815 10912
rect 9879 10848 9895 10912
rect 9959 10848 9967 10912
rect 9647 9824 9967 10848
rect 9647 9760 9655 9824
rect 9719 9760 9735 9824
rect 9799 9760 9815 9824
rect 9879 9760 9895 9824
rect 9959 9760 9967 9824
rect 9647 8736 9967 9760
rect 9647 8672 9655 8736
rect 9719 8672 9735 8736
rect 9799 8672 9815 8736
rect 9879 8672 9895 8736
rect 9959 8672 9967 8736
rect 9647 7648 9967 8672
rect 9647 7584 9655 7648
rect 9719 7584 9735 7648
rect 9799 7584 9815 7648
rect 9879 7584 9895 7648
rect 9959 7584 9967 7648
rect 9647 6560 9967 7584
rect 9647 6496 9655 6560
rect 9719 6496 9735 6560
rect 9799 6496 9815 6560
rect 9879 6496 9895 6560
rect 9959 6496 9967 6560
rect 9647 5472 9967 6496
rect 9647 5408 9655 5472
rect 9719 5408 9735 5472
rect 9799 5408 9815 5472
rect 9879 5408 9895 5472
rect 9959 5408 9967 5472
rect 9647 4384 9967 5408
rect 9647 4320 9655 4384
rect 9719 4320 9735 4384
rect 9799 4320 9815 4384
rect 9879 4320 9895 4384
rect 9959 4320 9967 4384
rect 9647 3296 9967 4320
rect 9647 3232 9655 3296
rect 9719 3232 9735 3296
rect 9799 3232 9815 3296
rect 9879 3232 9895 3296
rect 9959 3232 9967 3296
rect 9647 2208 9967 3232
rect 9647 2144 9655 2208
rect 9719 2144 9735 2208
rect 9799 2144 9815 2208
rect 9879 2144 9895 2208
rect 9959 2144 9967 2208
rect 9647 1120 9967 2144
rect 9647 1056 9655 1120
rect 9719 1056 9735 1120
rect 9799 1056 9815 1120
rect 9879 1056 9895 1120
rect 9959 1056 9967 1120
rect 9647 496 9967 1056
rect 11498 14720 11818 15280
rect 11498 14656 11506 14720
rect 11570 14656 11586 14720
rect 11650 14656 11666 14720
rect 11730 14656 11746 14720
rect 11810 14656 11818 14720
rect 11498 13632 11818 14656
rect 11498 13568 11506 13632
rect 11570 13568 11586 13632
rect 11650 13568 11666 13632
rect 11730 13568 11746 13632
rect 11810 13568 11818 13632
rect 11498 12544 11818 13568
rect 11498 12480 11506 12544
rect 11570 12480 11586 12544
rect 11650 12480 11666 12544
rect 11730 12480 11746 12544
rect 11810 12480 11818 12544
rect 11498 11456 11818 12480
rect 11498 11392 11506 11456
rect 11570 11392 11586 11456
rect 11650 11392 11666 11456
rect 11730 11392 11746 11456
rect 11810 11392 11818 11456
rect 11498 10368 11818 11392
rect 11498 10304 11506 10368
rect 11570 10304 11586 10368
rect 11650 10304 11666 10368
rect 11730 10304 11746 10368
rect 11810 10304 11818 10368
rect 11498 9280 11818 10304
rect 11498 9216 11506 9280
rect 11570 9216 11586 9280
rect 11650 9216 11666 9280
rect 11730 9216 11746 9280
rect 11810 9216 11818 9280
rect 11498 8192 11818 9216
rect 11498 8128 11506 8192
rect 11570 8128 11586 8192
rect 11650 8128 11666 8192
rect 11730 8128 11746 8192
rect 11810 8128 11818 8192
rect 11498 7104 11818 8128
rect 11498 7040 11506 7104
rect 11570 7040 11586 7104
rect 11650 7040 11666 7104
rect 11730 7040 11746 7104
rect 11810 7040 11818 7104
rect 11498 6016 11818 7040
rect 11498 5952 11506 6016
rect 11570 5952 11586 6016
rect 11650 5952 11666 6016
rect 11730 5952 11746 6016
rect 11810 5952 11818 6016
rect 11498 4928 11818 5952
rect 11498 4864 11506 4928
rect 11570 4864 11586 4928
rect 11650 4864 11666 4928
rect 11730 4864 11746 4928
rect 11810 4864 11818 4928
rect 11498 3840 11818 4864
rect 11498 3776 11506 3840
rect 11570 3776 11586 3840
rect 11650 3776 11666 3840
rect 11730 3776 11746 3840
rect 11810 3776 11818 3840
rect 11498 2752 11818 3776
rect 11498 2688 11506 2752
rect 11570 2688 11586 2752
rect 11650 2688 11666 2752
rect 11730 2688 11746 2752
rect 11810 2688 11818 2752
rect 11498 1664 11818 2688
rect 11498 1600 11506 1664
rect 11570 1600 11586 1664
rect 11650 1600 11666 1664
rect 11730 1600 11746 1664
rect 11810 1600 11818 1664
rect 11498 576 11818 1600
rect 11498 512 11506 576
rect 11570 512 11586 576
rect 11650 512 11666 576
rect 11730 512 11746 576
rect 11810 512 11818 576
rect 11498 496 11818 512
rect 13349 15264 13669 15280
rect 13349 15200 13357 15264
rect 13421 15200 13437 15264
rect 13501 15200 13517 15264
rect 13581 15200 13597 15264
rect 13661 15200 13669 15264
rect 13349 14176 13669 15200
rect 13349 14112 13357 14176
rect 13421 14112 13437 14176
rect 13501 14112 13517 14176
rect 13581 14112 13597 14176
rect 13661 14112 13669 14176
rect 13349 13088 13669 14112
rect 13349 13024 13357 13088
rect 13421 13024 13437 13088
rect 13501 13024 13517 13088
rect 13581 13024 13597 13088
rect 13661 13024 13669 13088
rect 13349 12000 13669 13024
rect 13349 11936 13357 12000
rect 13421 11936 13437 12000
rect 13501 11936 13517 12000
rect 13581 11936 13597 12000
rect 13661 11936 13669 12000
rect 13349 10912 13669 11936
rect 13349 10848 13357 10912
rect 13421 10848 13437 10912
rect 13501 10848 13517 10912
rect 13581 10848 13597 10912
rect 13661 10848 13669 10912
rect 13349 9824 13669 10848
rect 13349 9760 13357 9824
rect 13421 9760 13437 9824
rect 13501 9760 13517 9824
rect 13581 9760 13597 9824
rect 13661 9760 13669 9824
rect 13349 8736 13669 9760
rect 13349 8672 13357 8736
rect 13421 8672 13437 8736
rect 13501 8672 13517 8736
rect 13581 8672 13597 8736
rect 13661 8672 13669 8736
rect 13349 7648 13669 8672
rect 13349 7584 13357 7648
rect 13421 7584 13437 7648
rect 13501 7584 13517 7648
rect 13581 7584 13597 7648
rect 13661 7584 13669 7648
rect 13349 6560 13669 7584
rect 13349 6496 13357 6560
rect 13421 6496 13437 6560
rect 13501 6496 13517 6560
rect 13581 6496 13597 6560
rect 13661 6496 13669 6560
rect 13349 5472 13669 6496
rect 13349 5408 13357 5472
rect 13421 5408 13437 5472
rect 13501 5408 13517 5472
rect 13581 5408 13597 5472
rect 13661 5408 13669 5472
rect 13349 4384 13669 5408
rect 13349 4320 13357 4384
rect 13421 4320 13437 4384
rect 13501 4320 13517 4384
rect 13581 4320 13597 4384
rect 13661 4320 13669 4384
rect 13349 3296 13669 4320
rect 13349 3232 13357 3296
rect 13421 3232 13437 3296
rect 13501 3232 13517 3296
rect 13581 3232 13597 3296
rect 13661 3232 13669 3296
rect 13349 2208 13669 3232
rect 13349 2144 13357 2208
rect 13421 2144 13437 2208
rect 13501 2144 13517 2208
rect 13581 2144 13597 2208
rect 13661 2144 13669 2208
rect 13349 1120 13669 2144
rect 13349 1056 13357 1120
rect 13421 1056 13437 1120
rect 13501 1056 13517 1120
rect 13581 1056 13597 1120
rect 13661 1056 13669 1120
rect 13349 496 13669 1056
rect 15200 14720 15520 15280
rect 15200 14656 15208 14720
rect 15272 14656 15288 14720
rect 15352 14656 15368 14720
rect 15432 14656 15448 14720
rect 15512 14656 15520 14720
rect 15200 13632 15520 14656
rect 15200 13568 15208 13632
rect 15272 13568 15288 13632
rect 15352 13568 15368 13632
rect 15432 13568 15448 13632
rect 15512 13568 15520 13632
rect 15200 12544 15520 13568
rect 15200 12480 15208 12544
rect 15272 12480 15288 12544
rect 15352 12480 15368 12544
rect 15432 12480 15448 12544
rect 15512 12480 15520 12544
rect 15200 11456 15520 12480
rect 15200 11392 15208 11456
rect 15272 11392 15288 11456
rect 15352 11392 15368 11456
rect 15432 11392 15448 11456
rect 15512 11392 15520 11456
rect 15200 10368 15520 11392
rect 15200 10304 15208 10368
rect 15272 10304 15288 10368
rect 15352 10304 15368 10368
rect 15432 10304 15448 10368
rect 15512 10304 15520 10368
rect 15200 9280 15520 10304
rect 15200 9216 15208 9280
rect 15272 9216 15288 9280
rect 15352 9216 15368 9280
rect 15432 9216 15448 9280
rect 15512 9216 15520 9280
rect 15200 8192 15520 9216
rect 15200 8128 15208 8192
rect 15272 8128 15288 8192
rect 15352 8128 15368 8192
rect 15432 8128 15448 8192
rect 15512 8128 15520 8192
rect 15200 7104 15520 8128
rect 15200 7040 15208 7104
rect 15272 7040 15288 7104
rect 15352 7040 15368 7104
rect 15432 7040 15448 7104
rect 15512 7040 15520 7104
rect 15200 6016 15520 7040
rect 15200 5952 15208 6016
rect 15272 5952 15288 6016
rect 15352 5952 15368 6016
rect 15432 5952 15448 6016
rect 15512 5952 15520 6016
rect 15200 4928 15520 5952
rect 15200 4864 15208 4928
rect 15272 4864 15288 4928
rect 15352 4864 15368 4928
rect 15432 4864 15448 4928
rect 15512 4864 15520 4928
rect 15200 3840 15520 4864
rect 15200 3776 15208 3840
rect 15272 3776 15288 3840
rect 15352 3776 15368 3840
rect 15432 3776 15448 3840
rect 15512 3776 15520 3840
rect 15200 2752 15520 3776
rect 15200 2688 15208 2752
rect 15272 2688 15288 2752
rect 15352 2688 15368 2752
rect 15432 2688 15448 2752
rect 15512 2688 15520 2752
rect 15200 1664 15520 2688
rect 15200 1600 15208 1664
rect 15272 1600 15288 1664
rect 15352 1600 15368 1664
rect 15432 1600 15448 1664
rect 15512 1600 15520 1664
rect 15200 576 15520 1600
rect 15200 512 15208 576
rect 15272 512 15288 576
rect 15352 512 15368 576
rect 15432 512 15448 576
rect 15512 512 15520 576
rect 15200 496 15520 512
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1685868990
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1685868990
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1685868990
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1685868990
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1685868990
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1685868990
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1685868990
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1685868990
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1685868990
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1685868990
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1685868990
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1685868990
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1685868990
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 14628 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_157
timestamp 1685868990
transform 1 0 14996 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1685868990
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1685868990
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1685868990
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1685868990
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1685868990
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1685868990
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1685868990
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1685868990
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1685868990
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1685868990
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1685868990
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1685868990
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1685868990
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1685868990
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_149 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 14260 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_157
timestamp 1685868990
transform 1 0 14996 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1685868990
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1685868990
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1685868990
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1685868990
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1685868990
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1685868990
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1685868990
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1685868990
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1685868990
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1685868990
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1685868990
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1685868990
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1685868990
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1685868990
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1685868990
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1685868990
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_153
timestamp 1685868990
transform 1 0 14628 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_157
timestamp 1685868990
transform 1 0 14996 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1685868990
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1685868990
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1685868990
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1685868990
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1685868990
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1685868990
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1685868990
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1685868990
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1685868990
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1685868990
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1685868990
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1685868990
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1685868990
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1685868990
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1685868990
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_149
timestamp 1685868990
transform 1 0 14260 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_157
timestamp 1685868990
transform 1 0 14996 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1685868990
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1685868990
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1685868990
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1685868990
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1685868990
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1685868990
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1685868990
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1685868990
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1685868990
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1685868990
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1685868990
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1685868990
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1685868990
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1685868990
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1685868990
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1685868990
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_153
timestamp 1685868990
transform 1 0 14628 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_157
timestamp 1685868990
transform 1 0 14996 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1685868990
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1685868990
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1685868990
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1685868990
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1685868990
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1685868990
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1685868990
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1685868990
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1685868990
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1685868990
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1685868990
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1685868990
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1685868990
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1685868990
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1685868990
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_149
timestamp 1685868990
transform 1 0 14260 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_157
timestamp 1685868990
transform 1 0 14996 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1685868990
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1685868990
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1685868990
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1685868990
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1685868990
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1685868990
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1685868990
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1685868990
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1685868990
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1685868990
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_97 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_118
timestamp 1685868990
transform 1 0 11408 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_130
timestamp 1685868990
transform 1 0 12512 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1685868990
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1685868990
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_153
timestamp 1685868990
transform 1 0 14628 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_157
timestamp 1685868990
transform 1 0 14996 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1685868990
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1685868990
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1685868990
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1685868990
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1685868990
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1685868990
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1685868990
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1685868990
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1685868990
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1685868990
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1685868990
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1685868990
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1685868990
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1685868990
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1685868990
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_149
timestamp 1685868990
transform 1 0 14260 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_157
timestamp 1685868990
transform 1 0 14996 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1685868990
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1685868990
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1685868990
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_29
timestamp 1685868990
transform 1 0 3220 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_46
timestamp 1685868990
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_64
timestamp 1685868990
transform 1 0 6440 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_85
timestamp 1685868990
transform 1 0 8372 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_107
timestamp 1685868990
transform 1 0 10396 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_115
timestamp 1685868990
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_136
timestamp 1685868990
transform 1 0 13064 0 1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1685868990
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_153
timestamp 1685868990
transform 1 0 14628 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_157
timestamp 1685868990
transform 1 0 14996 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1685868990
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1685868990
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_27
timestamp 1685868990
transform 1 0 3036 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_33
timestamp 1685868990
transform 1 0 3588 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_41
timestamp 1685868990
transform 1 0 4324 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 1685868990
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_57
timestamp 1685868990
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_99
timestamp 1685868990
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1685868990
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_113
timestamp 1685868990
transform 1 0 10948 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_120
timestamp 1685868990
transform 1 0 11592 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_130
timestamp 1685868990
transform 1 0 12512 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_152
timestamp 1685868990
transform 1 0 14536 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_3
timestamp 1685868990
transform 1 0 828 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_29
timestamp 1685868990
transform 1 0 3220 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_35
timestamp 1685868990
transform 1 0 3772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_46
timestamp 1685868990
transform 1 0 4784 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_54
timestamp 1685868990
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_75
timestamp 1685868990
transform 1 0 7452 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1685868990
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_93
timestamp 1685868990
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_105
timestamp 1685868990
transform 1 0 10212 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_111
timestamp 1685868990
transform 1 0 10764 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_119
timestamp 1685868990
transform 1 0 11500 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_127
timestamp 1685868990
transform 1 0 12236 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1685868990
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_156
timestamp 1685868990
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1685868990
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_15
timestamp 1685868990
transform 1 0 1932 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_23
timestamp 1685868990
transform 1 0 2668 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_42
timestamp 1685868990
transform 1 0 4416 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_50
timestamp 1685868990
transform 1 0 5152 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1685868990
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_57
timestamp 1685868990
transform 1 0 5796 0 -1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_72
timestamp 1685868990
transform 1 0 7176 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_84
timestamp 1685868990
transform 1 0 8280 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_96
timestamp 1685868990
transform 1 0 9384 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_108
timestamp 1685868990
transform 1 0 10488 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_113
timestamp 1685868990
transform 1 0 10948 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_121
timestamp 1685868990
transform 1 0 11684 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_128
timestamp 1685868990
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_135
timestamp 1685868990
transform 1 0 12972 0 -1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1685868990
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1685868990
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1685868990
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_29
timestamp 1685868990
transform 1 0 3220 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_47
timestamp 1685868990
transform 1 0 4876 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_64
timestamp 1685868990
transform 1 0 6440 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_76
timestamp 1685868990
transform 1 0 7544 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1685868990
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1685868990
transform 1 0 8372 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_93
timestamp 1685868990
transform 1 0 9108 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_108
timestamp 1685868990
transform 1 0 10488 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_121
timestamp 1685868990
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_132
timestamp 1685868990
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1685868990
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_149
timestamp 1685868990
transform 1 0 14260 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_157
timestamp 1685868990
transform 1 0 14996 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1685868990
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_15
timestamp 1685868990
transform 1 0 1932 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_49
timestamp 1685868990
transform 1 0 5060 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1685868990
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1685868990
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_69
timestamp 1685868990
transform 1 0 6900 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_73
timestamp 1685868990
transform 1 0 7268 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1685868990
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1685868990
transform 1 0 10212 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1685868990
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_113
timestamp 1685868990
transform 1 0 10948 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_121
timestamp 1685868990
transform 1 0 11684 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_142
timestamp 1685868990
transform 1 0 13616 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_154
timestamp 1685868990
transform 1 0 14720 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_3
timestamp 1685868990
transform 1 0 828 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_9
timestamp 1685868990
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1685868990
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_33
timestamp 1685868990
transform 1 0 3588 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_51
timestamp 1685868990
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_57
timestamp 1685868990
transform 1 0 5796 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_61
timestamp 1685868990
transform 1 0 6164 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_67
timestamp 1685868990
transform 1 0 6716 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_79
timestamp 1685868990
transform 1 0 7820 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1685868990
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_100
timestamp 1685868990
transform 1 0 9752 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_117
timestamp 1685868990
transform 1 0 11316 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_129
timestamp 1685868990
transform 1 0 12420 0 1 8160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_144
timestamp 1685868990
transform 1 0 13800 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_156
timestamp 1685868990
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1685868990
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_23
timestamp 1685868990
transform 1 0 2668 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_32
timestamp 1685868990
transform 1 0 3496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_39
timestamp 1685868990
transform 1 0 4140 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_45
timestamp 1685868990
transform 1 0 4692 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_49
timestamp 1685868990
transform 1 0 5060 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1685868990
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1685868990
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_129
timestamp 1685868990
transform 1 0 12420 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_3
timestamp 1685868990
transform 1 0 828 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_11
timestamp 1685868990
transform 1 0 1564 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_50
timestamp 1685868990
transform 1 0 5152 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_60
timestamp 1685868990
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_65
timestamp 1685868990
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1685868990
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_101
timestamp 1685868990
transform 1 0 9844 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_109
timestamp 1685868990
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_138
timestamp 1685868990
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_153
timestamp 1685868990
transform 1 0 14628 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_157
timestamp 1685868990
transform 1 0 14996 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1685868990
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1685868990
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1685868990
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_39
timestamp 1685868990
transform 1 0 4140 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_46
timestamp 1685868990
transform 1 0 4784 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_50
timestamp 1685868990
transform 1 0 5152 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1685868990
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1685868990
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1685868990
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_81
timestamp 1685868990
transform 1 0 8004 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_101
timestamp 1685868990
transform 1 0 9844 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1685868990
transform 1 0 10580 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_113
timestamp 1685868990
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_122
timestamp 1685868990
transform 1 0 11776 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_134
timestamp 1685868990
transform 1 0 12880 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_146
timestamp 1685868990
transform 1 0 13984 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1685868990
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_15
timestamp 1685868990
transform 1 0 1932 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_26
timestamp 1685868990
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_72
timestamp 1685868990
transform 1 0 7176 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_80
timestamp 1685868990
transform 1 0 7912 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_105
timestamp 1685868990
transform 1 0 10212 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_122
timestamp 1685868990
transform 1 0 11776 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_154
timestamp 1685868990
transform 1 0 14720 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_3
timestamp 1685868990
transform 1 0 828 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1685868990
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_57
timestamp 1685868990
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_75
timestamp 1685868990
transform 1 0 7452 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_87
timestamp 1685868990
transform 1 0 8556 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_105
timestamp 1685868990
transform 1 0 10212 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_127
timestamp 1685868990
transform 1 0 12236 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1685868990
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_15
timestamp 1685868990
transform 1 0 1932 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_24
timestamp 1685868990
transform 1 0 2760 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_29
timestamp 1685868990
transform 1 0 3220 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_40
timestamp 1685868990
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_49
timestamp 1685868990
transform 1 0 5060 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_59
timestamp 1685868990
transform 1 0 5980 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_66
timestamp 1685868990
transform 1 0 6624 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_74
timestamp 1685868990
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_108
timestamp 1685868990
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_119
timestamp 1685868990
transform 1 0 11500 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_126
timestamp 1685868990
transform 1 0 12144 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1685868990
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1685868990
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_153
timestamp 1685868990
transform 1 0 14628 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_157
timestamp 1685868990
transform 1 0 14996 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1685868990
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_15
timestamp 1685868990
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_33
timestamp 1685868990
transform 1 0 3588 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_37
timestamp 1685868990
transform 1 0 3956 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_43
timestamp 1685868990
transform 1 0 4508 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1685868990
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_57
timestamp 1685868990
transform 1 0 5796 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_66
timestamp 1685868990
transform 1 0 6624 0 -1 12512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_79
timestamp 1685868990
transform 1 0 7820 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_91
timestamp 1685868990
transform 1 0 8924 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_102
timestamp 1685868990
transform 1 0 9936 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1685868990
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_113
timestamp 1685868990
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_122
timestamp 1685868990
transform 1 0 11776 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_134
timestamp 1685868990
transform 1 0 12880 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_138
timestamp 1685868990
transform 1 0 13248 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1685868990
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1685868990
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1685868990
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_29
timestamp 1685868990
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_47
timestamp 1685868990
transform 1 0 4876 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_63
timestamp 1685868990
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1685868990
transform 1 0 8004 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_85
timestamp 1685868990
transform 1 0 8372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_107
timestamp 1685868990
transform 1 0 10396 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_127
timestamp 1685868990
transform 1 0 12236 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_152
timestamp 1685868990
transform 1 0 14536 0 1 12512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1685868990
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1685868990
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1685868990
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1685868990
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1685868990
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1685868990
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_57
timestamp 1685868990
transform 1 0 5796 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_63
timestamp 1685868990
transform 1 0 6348 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_67
timestamp 1685868990
transform 1 0 6716 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_75
timestamp 1685868990
transform 1 0 7452 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_91
timestamp 1685868990
transform 1 0 8924 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_107
timestamp 1685868990
transform 1 0 10396 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1685868990
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_113
timestamp 1685868990
transform 1 0 10948 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_124
timestamp 1685868990
transform 1 0 11960 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_132
timestamp 1685868990
transform 1 0 12696 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_151
timestamp 1685868990
transform 1 0 14444 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_157
timestamp 1685868990
transform 1 0 14996 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1685868990
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_15
timestamp 1685868990
transform 1 0 1932 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_24
timestamp 1685868990
transform 1 0 2760 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_29
timestamp 1685868990
transform 1 0 3220 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_48
timestamp 1685868990
transform 1 0 4968 0 1 13600
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_69
timestamp 1685868990
transform 1 0 6900 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1685868990
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_93
timestamp 1685868990
transform 1 0 9108 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_97
timestamp 1685868990
transform 1 0 9476 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_106
timestamp 1685868990
transform 1 0 10304 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_114
timestamp 1685868990
transform 1 0 11040 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_125
timestamp 1685868990
transform 1 0 12052 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_133
timestamp 1685868990
transform 1 0 12788 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1685868990
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_145
timestamp 1685868990
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_155
timestamp 1685868990
transform 1 0 14812 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_3
timestamp 1685868990
transform 1 0 828 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_11
timestamp 1685868990
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_57
timestamp 1685868990
transform 1 0 5796 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_86
timestamp 1685868990
transform 1 0 8464 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_90
timestamp 1685868990
transform 1 0 8832 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_107
timestamp 1685868990
transform 1 0 10396 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1685868990
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_129
timestamp 1685868990
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1685868990
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_15
timestamp 1685868990
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_23
timestamp 1685868990
transform 1 0 2668 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1685868990
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_29
timestamp 1685868990
transform 1 0 3220 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_36
timestamp 1685868990
transform 1 0 3864 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_44
timestamp 1685868990
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_50
timestamp 1685868990
transform 1 0 5152 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_67
timestamp 1685868990
transform 1 0 6716 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_73
timestamp 1685868990
transform 1 0 7268 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1685868990
transform 1 0 7636 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1685868990
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_95
timestamp 1685868990
transform 1 0 9292 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_108
timestamp 1685868990
transform 1 0 10488 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_113
timestamp 1685868990
transform 1 0 10948 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_127
timestamp 1685868990
transform 1 0 12236 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_133
timestamp 1685868990
transform 1 0 12788 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_141
timestamp 1685868990
transform 1 0 13524 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_147
timestamp 1685868990
transform 1 0 14076 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1685868990
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1685868990
transform -1 0 15364 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1685868990
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1685868990
transform -1 0 15364 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1685868990
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1685868990
transform -1 0 15364 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1685868990
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1685868990
transform -1 0 15364 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1685868990
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1685868990
transform -1 0 15364 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1685868990
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1685868990
transform -1 0 15364 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1685868990
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1685868990
transform -1 0 15364 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1685868990
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1685868990
transform -1 0 15364 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1685868990
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1685868990
transform -1 0 15364 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1685868990
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1685868990
transform -1 0 15364 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1685868990
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1685868990
transform -1 0 15364 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1685868990
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1685868990
transform -1 0 15364 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1685868990
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1685868990
transform -1 0 15364 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1685868990
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1685868990
transform -1 0 15364 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1685868990
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1685868990
transform -1 0 15364 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1685868990
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1685868990
transform -1 0 15364 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1685868990
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1685868990
transform -1 0 15364 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1685868990
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1685868990
transform -1 0 15364 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1685868990
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1685868990
transform -1 0 15364 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1685868990
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1685868990
transform -1 0 15364 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1685868990
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1685868990
transform -1 0 15364 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1685868990
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1685868990
transform -1 0 15364 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1685868990
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1685868990
transform -1 0 15364 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1685868990
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1685868990
transform -1 0 15364 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1685868990
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1685868990
transform -1 0 15364 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1685868990
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1685868990
transform -1 0 15364 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1685868990
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1685868990
transform -1 0 15364 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1685868990
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1685868990
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1685868990
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1685868990
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1685868990
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1685868990
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1685868990
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1685868990
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1685868990
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1685868990
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1685868990
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1685868990
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1685868990
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1685868990
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1685868990
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1685868990
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1685868990
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1685868990
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1685868990
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1685868990
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1685868990
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1685868990
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1685868990
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1685868990
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1685868990
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1685868990
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1685868990
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1685868990
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1685868990
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1685868990
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1685868990
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1685868990
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1685868990
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1685868990
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1685868990
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1685868990
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1685868990
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1685868990
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1685868990
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1685868990
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1685868990
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1685868990
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1685868990
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1685868990
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1685868990
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1685868990
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1685868990
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1685868990
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1685868990
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1685868990
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1685868990
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1685868990
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1685868990
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1685868990
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1685868990
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1685868990
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1685868990
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1685868990
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1685868990
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1685868990
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1685868990
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1685868990
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1685868990
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1685868990
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1685868990
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1685868990
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1685868990
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1685868990
transform 1 0 5704 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1685868990
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1685868990
transform 1 0 10856 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1685868990
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12880 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _166_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 14352 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11224 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13524 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12512 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12880 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14720 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _172_
timestamp 1685868990
transform -1 0 12604 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _173_
timestamp 1676037725
transform 1 0 12604 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _174_
timestamp 1685868990
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _175_
timestamp 1685868990
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 12512 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 13984 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _179_
timestamp 1685868990
transform -1 0 13984 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _180_
timestamp 1685868990
transform -1 0 13248 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13340 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _182_
timestamp 1685868990
transform 1 0 13156 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _183_
timestamp 1685868990
transform -1 0 13432 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _184_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12880 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13524 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _186_
timestamp 1676037725
transform 1 0 9844 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 9292 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _188_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 5704 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7544 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9108 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _191_
timestamp 1685868990
transform -1 0 7820 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _192_
timestamp 1676037725
transform -1 0 6808 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _193_
timestamp 1676037725
transform 1 0 5980 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 7452 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5704 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _196_
timestamp 1685868990
transform -1 0 5520 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6440 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _198_
timestamp 1685868990
transform 1 0 6164 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp 1685868990
transform 1 0 7912 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _200_
timestamp 1676037725
transform 1 0 6440 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _201_
timestamp 1685868990
transform -1 0 5520 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _202_
timestamp 1685868990
transform -1 0 4324 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _203_
timestamp 1685868990
transform 1 0 4508 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _204_
timestamp 1685868990
transform -1 0 4416 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4508 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _206_
timestamp 1676037725
transform 1 0 3680 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4140 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _208_
timestamp 1676037725
transform 1 0 2760 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _209_
timestamp 1685868990
transform 1 0 2852 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _210_
timestamp 1685868990
transform 1 0 2300 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5060 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _213_
timestamp 1676037725
transform -1 0 4600 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _214_
timestamp 1676037725
transform 1 0 3220 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _215_
timestamp 1685868990
transform -1 0 4140 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _216_
timestamp 1685868990
transform 1 0 4416 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _217_
timestamp 1676037725
transform 1 0 4600 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1685868990
transform 1 0 4784 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _219_
timestamp 1676037725
transform 1 0 3220 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _220_
timestamp 1685868990
transform 1 0 3220 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _221_
timestamp 1685868990
transform 1 0 5520 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _222_
timestamp 1685868990
transform -1 0 5520 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _223_
timestamp 1676037725
transform 1 0 6440 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _224_
timestamp 1685868990
transform 1 0 5980 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 6348 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1685868990
transform -1 0 5520 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _227_
timestamp 1685868990
transform -1 0 5520 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _228_
timestamp 1676037725
transform -1 0 4784 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _229_
timestamp 1676037725
transform 1 0 4140 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _230_
timestamp 1685868990
transform -1 0 3956 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _231_
timestamp 1685868990
transform 1 0 2668 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _232_
timestamp 1685868990
transform 1 0 3864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 3220 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _234_
timestamp 1676037725
transform 1 0 2300 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _235_
timestamp 1676037725
transform 1 0 4876 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _236_
timestamp 1676037725
transform 1 0 4416 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _237_
timestamp 1676037725
transform 1 0 4692 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _238_
timestamp 1676037725
transform 1 0 3496 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _239_
timestamp 1685868990
transform 1 0 2484 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _240_
timestamp 1685868990
transform -1 0 7912 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _241_
timestamp 1685868990
transform 1 0 5244 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _242_
timestamp 1685868990
transform -1 0 8188 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _243_
timestamp 1676037725
transform 1 0 6716 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _244_
timestamp 1685868990
transform -1 0 6716 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _245_
timestamp 1685868990
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _246_
timestamp 1676037725
transform -1 0 9476 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _247_
timestamp 1676037725
transform 1 0 8372 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _248_
timestamp 1676037725
transform 1 0 8372 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _249_
timestamp 1685868990
transform -1 0 7912 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _250_
timestamp 1676037725
transform 1 0 10396 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _251_
timestamp 1676037725
transform 1 0 8832 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _252_
timestamp 1676037725
transform -1 0 9660 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _253_
timestamp 1685868990
transform -1 0 10396 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1685868990
transform -1 0 11040 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _255_
timestamp 1676037725
transform -1 0 11776 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1685868990
transform -1 0 2760 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _258_
timestamp 1685868990
transform 1 0 6624 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _259_
timestamp 1676037725
transform 1 0 3680 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _260_
timestamp 1676037725
transform -1 0 6900 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6256 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _262_
timestamp 1676037725
transform -1 0 6440 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _263_
timestamp 1676037725
transform 1 0 5888 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _264_
timestamp 1676037725
transform -1 0 8924 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _265_
timestamp 1676037725
transform -1 0 8280 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _266_
timestamp 1676037725
transform 1 0 8372 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _267_
timestamp 1676037725
transform -1 0 9108 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _268_
timestamp 1676037725
transform -1 0 10212 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _269_
timestamp 1676037725
transform 1 0 9568 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1685868990
transform -1 0 8924 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9476 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _272_
timestamp 1676037725
transform -1 0 10396 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _273_
timestamp 1676037725
transform -1 0 11776 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _274_
timestamp 1676037725
transform 1 0 11224 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _275_
timestamp 1676037725
transform -1 0 11960 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _276_
timestamp 1676037725
transform 1 0 11316 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1685868990
transform 1 0 5704 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 5244 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 5152 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _280_
timestamp 1685868990
transform 1 0 5796 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _281_
timestamp 1676037725
transform 1 0 5888 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1685868990
transform 1 0 4232 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7820 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _284_
timestamp 1685868990
transform 1 0 10672 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _285_
timestamp 1676037725
transform -1 0 12236 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _286_
timestamp 1685868990
transform 1 0 10304 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _287_
timestamp 1676037725
transform -1 0 11592 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1685868990
transform -1 0 8280 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _289_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9200 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _290_
timestamp 1685868990
transform -1 0 10488 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _291_
timestamp 1676037725
transform 1 0 7544 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _292_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9200 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1685868990
transform -1 0 9752 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _294_
timestamp 1676037725
transform -1 0 9568 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1685868990
transform -1 0 11500 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _296_
timestamp 1685868990
transform -1 0 12144 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _297_
timestamp 1685868990
transform 1 0 10488 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9568 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _299_
timestamp 1685868990
transform -1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _300_
timestamp 1676037725
transform 1 0 9292 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _301_
timestamp 1676037725
transform -1 0 12420 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _302_
timestamp 1685868990
transform 1 0 11408 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _303_
timestamp 1676037725
transform -1 0 9752 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1685868990
transform 1 0 6440 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _305_
timestamp 1676037725
transform 1 0 9752 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _306_
timestamp 1676037725
transform 1 0 10120 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _307_
timestamp 1685868990
transform -1 0 9016 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _308_
timestamp 1676037725
transform 1 0 9292 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _309_
timestamp 1676037725
transform 1 0 10856 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _310_
timestamp 1685868990
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11408 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _312_
timestamp 1685868990
transform 1 0 11224 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _313_
timestamp 1676037725
transform 1 0 11960 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _314_
timestamp 1676037725
transform -1 0 11592 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _315_
timestamp 1685868990
transform 1 0 5428 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _316_
timestamp 1685868990
transform 1 0 8832 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _317_
timestamp 1676037725
transform -1 0 12328 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _318_
timestamp 1676037725
transform -1 0 12972 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _319_
timestamp 1676037725
transform -1 0 12880 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _320_
timestamp 1676037725
transform -1 0 12420 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _321_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12512 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _322_
timestamp 1676037725
transform -1 0 14904 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _323_
timestamp 1685868990
transform 1 0 13524 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _324_
timestamp 1685868990
transform 1 0 12880 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4232 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _326_
timestamp 1676037725
transform 1 0 3496 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _327_
timestamp 1676037725
transform -1 0 8004 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _328_
timestamp 1676037725
transform -1 0 8464 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _329_
timestamp 1676037725
transform -1 0 10396 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _330_
timestamp 1676037725
transform -1 0 10396 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _331_
timestamp 1676037725
transform -1 0 12236 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _332_
timestamp 1676037725
transform -1 0 12420 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _333_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9660 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _334_
timestamp 1676037725
transform 1 0 11316 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _335_
timestamp 1676037725
transform 1 0 12788 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _336_
timestamp 1676037725
transform 1 0 13340 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _337_
timestamp 1676037725
transform 1 0 13340 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _338_
timestamp 1676037725
transform 1 0 13340 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _339_
timestamp 1676037725
transform 1 0 13340 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _340_
timestamp 1676037725
transform 1 0 13340 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _341_
timestamp 1676037725
transform 1 0 8924 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _342_
timestamp 1676037725
transform -1 0 8280 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _343_
timestamp 1676037725
transform 1 0 4968 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _344_
timestamp 1676037725
transform 1 0 4968 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _345_
timestamp 1676037725
transform 1 0 3312 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _346_
timestamp 1676037725
transform 1 0 1380 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _347_
timestamp 1676037725
transform 1 0 1472 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _348_
timestamp 1676037725
transform 1 0 1656 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _349_
timestamp 1676037725
transform 1 0 5980 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _350_
timestamp 1676037725
transform 1 0 3404 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _351_
timestamp 1676037725
transform -1 0 2484 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _352_
timestamp 1676037725
transform 1 0 2116 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _353_
timestamp 1676037725
transform 1 0 5796 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _354_
timestamp 1676037725
transform 1 0 7360 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _355_
timestamp 1676037725
transform 1 0 9844 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _356_
timestamp 1676037725
transform 1 0 11040 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _357__12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 2116 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _357_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1748 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7268 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1676037725
transform -1 0 5060 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1676037725
transform 1 0 7820 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1676037725
transform 1 0 8372 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2668 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1676037725
transform -1 0 5244 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1676037725
transform -1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1676037725
transform 1 0 6808 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1676037725
transform 1 0 6808 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1676037725
transform 1 0 3956 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1676037725
transform -1 0 13248 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1676037725
transform -1 0 10764 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1676037725
transform -1 0 14260 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1676037725
transform -1 0 14812 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1676037725
transform 1 0 4876 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1676037725
transform -1 0 11684 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1676037725
transform 1 0 7360 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1676037725
transform -1 0 9292 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1676037725
transform 1 0 10212 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1676037725
transform 1 0 11960 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1676037725
transform 1 0 12512 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1685868990
transform -1 0 14076 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1676037725
transform -1 0 15088 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1676037725
transform 1 0 4784 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1685868990
transform -1 0 2668 0 1 14688
box -38 -48 314 592
<< labels >>
flabel metal4 s 4094 496 4414 15280 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7796 496 8116 15280 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11498 496 11818 15280 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15200 496 15520 15280 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2243 496 2563 15280 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5945 496 6265 15280 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9647 496 9967 15280 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13349 496 13669 15280 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 846 15600 902 16000 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal2 s 5998 15600 6054 16000 0 FreeSans 224 90 0 0 data[0]
port 3 nsew signal input
flabel metal2 s 7286 15600 7342 16000 0 FreeSans 224 90 0 0 data[1]
port 4 nsew signal input
flabel metal2 s 8574 15600 8630 16000 0 FreeSans 224 90 0 0 data[2]
port 5 nsew signal input
flabel metal2 s 9862 15600 9918 16000 0 FreeSans 224 90 0 0 data[3]
port 6 nsew signal input
flabel metal2 s 11150 15600 11206 16000 0 FreeSans 224 90 0 0 data[4]
port 7 nsew signal input
flabel metal2 s 12438 15600 12494 16000 0 FreeSans 224 90 0 0 data[5]
port 8 nsew signal input
flabel metal2 s 13726 15600 13782 16000 0 FreeSans 224 90 0 0 data[6]
port 9 nsew signal input
flabel metal2 s 15014 15600 15070 16000 0 FreeSans 224 90 0 0 data[7]
port 10 nsew signal input
flabel metal2 s 3422 15600 3478 16000 0 FreeSans 224 90 0 0 ext_data
port 11 nsew signal input
flabel metal2 s 4710 15600 4766 16000 0 FreeSans 224 90 0 0 load_divider
port 12 nsew signal input
flabel metal2 s 2134 15600 2190 16000 0 FreeSans 224 90 0 0 n_rst
port 13 nsew signal input
flabel metal3 s 15600 1096 16000 1216 0 FreeSans 480 0 0 0 r2r_out[0]
port 14 nsew signal tristate
flabel metal3 s 15600 3000 16000 3120 0 FreeSans 480 0 0 0 r2r_out[1]
port 15 nsew signal tristate
flabel metal3 s 15600 4904 16000 5024 0 FreeSans 480 0 0 0 r2r_out[2]
port 16 nsew signal tristate
flabel metal3 s 15600 6808 16000 6928 0 FreeSans 480 0 0 0 r2r_out[3]
port 17 nsew signal tristate
flabel metal3 s 15600 8712 16000 8832 0 FreeSans 480 0 0 0 r2r_out[4]
port 18 nsew signal tristate
flabel metal3 s 15600 10616 16000 10736 0 FreeSans 480 0 0 0 r2r_out[5]
port 19 nsew signal tristate
flabel metal3 s 15600 12520 16000 12640 0 FreeSans 480 0 0 0 r2r_out[6]
port 20 nsew signal tristate
flabel metal3 s 15600 14424 16000 14544 0 FreeSans 480 0 0 0 r2r_out[7]
port 21 nsew signal tristate
rlabel via1 8036 14688 8036 14688 0 VGND
rlabel metal1 7958 15232 7958 15232 0 VPWR
rlabel metal1 2714 13974 2714 13974 0 _000_
rlabel metal2 5566 14144 5566 14144 0 _001_
rlabel metal1 4503 13838 4503 13838 0 _002_
rlabel via1 7686 12750 7686 12750 0 _003_
rlabel metal1 8372 14042 8372 14042 0 _004_
rlabel metal2 10258 14246 10258 14246 0 _005_
rlabel via1 10078 12682 10078 12682 0 _006_
rlabel via1 11918 12682 11918 12682 0 _007_
rlabel metal1 12052 14042 12052 14042 0 _008_
rlabel metal2 10074 4148 10074 4148 0 _009_
rlabel metal2 11638 5338 11638 5338 0 _010_
rlabel metal1 12834 5746 12834 5746 0 _011_
rlabel metal1 13616 7174 13616 7174 0 _012_
rlabel metal1 13478 9010 13478 9010 0 _013_
rlabel metal1 13662 10778 13662 10778 0 _014_
rlabel metal1 13800 12274 13800 12274 0 _015_
rlabel metal1 13708 14382 13708 14382 0 _016_
rlabel metal1 9287 5066 9287 5066 0 _017_
rlabel via1 7962 5134 7962 5134 0 _018_
rlabel via1 5285 5134 5285 5134 0 _019_
rlabel metal2 5382 7106 5382 7106 0 _020_
rlabel metal1 3675 5066 3675 5066 0 _021_
rlabel metal1 2341 6154 2341 6154 0 _022_
rlabel metal1 2990 8364 2990 8364 0 _023_
rlabel metal2 3358 9282 3358 9282 0 _024_
rlabel metal1 6343 11254 6343 11254 0 _025_
rlabel metal1 3767 12682 3767 12682 0 _026_
rlabel via1 2166 11186 2166 11186 0 _027_
rlabel metal1 2576 11866 2576 11866 0 _028_
rlabel metal1 6205 9078 6205 9078 0 _029_
rlabel metal1 7774 7514 7774 7514 0 _030_
rlabel via1 10161 8398 10161 8398 0 _031_
rlabel metal1 11592 9146 11592 9146 0 _032_
rlabel metal2 5934 12444 5934 12444 0 _033_
rlabel metal1 7866 11526 7866 11526 0 _034_
rlabel metal1 4278 11662 4278 11662 0 _035_
rlabel metal1 8326 11662 8326 11662 0 _036_
rlabel metal2 11178 11356 11178 11356 0 _037_
rlabel metal1 10810 10608 10810 10608 0 _038_
rlabel metal2 10902 10846 10902 10846 0 _039_
rlabel metal1 9798 11254 9798 11254 0 _040_
rlabel metal1 8142 11594 8142 11594 0 _041_
rlabel metal1 9016 11798 9016 11798 0 _042_
rlabel metal1 9614 11526 9614 11526 0 _043_
rlabel metal1 8556 11866 8556 11866 0 _044_
rlabel metal1 9108 10098 9108 10098 0 _045_
rlabel metal1 9016 8398 9016 8398 0 _046_
rlabel metal1 9706 11050 9706 11050 0 _047_
rlabel metal1 10994 10540 10994 10540 0 _048_
rlabel metal1 11316 10574 11316 10574 0 _049_
rlabel metal1 10304 10710 10304 10710 0 _050_
rlabel metal1 9292 10098 9292 10098 0 _051_
rlabel metal1 5106 8568 5106 8568 0 _052_
rlabel metal1 10534 9010 10534 9010 0 _053_
rlabel metal2 9522 7072 9522 7072 0 _054_
rlabel metal1 9614 7446 9614 7446 0 _055_
rlabel metal1 9798 7446 9798 7446 0 _056_
rlabel metal1 6118 10608 6118 10608 0 _057_
rlabel metal1 10120 7242 10120 7242 0 _058_
rlabel metal2 6992 9486 6992 9486 0 _059_
rlabel metal1 9292 9010 9292 9010 0 _060_
rlabel metal1 11362 5712 11362 5712 0 _061_
rlabel metal1 11178 7378 11178 7378 0 _062_
rlabel metal1 11040 7174 11040 7174 0 _063_
rlabel metal1 11270 5780 11270 5780 0 _064_
rlabel metal1 3680 12274 3680 12274 0 _065_
rlabel metal1 2852 10574 2852 10574 0 _066_
rlabel metal1 12098 7820 12098 7820 0 _067_
rlabel metal1 12466 6698 12466 6698 0 _068_
rlabel metal1 12742 7242 12742 7242 0 _069_
rlabel metal1 12190 7820 12190 7820 0 _070_
rlabel metal1 12558 6222 12558 6222 0 _071_
rlabel metal1 13570 8364 13570 8364 0 _072_
rlabel metal1 13202 8432 13202 8432 0 _073_
rlabel metal1 13202 7514 13202 7514 0 _074_
rlabel metal2 14030 7514 14030 7514 0 _075_
rlabel metal1 13064 8602 13064 8602 0 _076_
rlabel metal1 14260 9350 14260 9350 0 _077_
rlabel metal2 3726 9214 3726 9214 0 _078_
rlabel metal1 12742 9044 12742 9044 0 _079_
rlabel metal2 12926 10982 12926 10982 0 _080_
rlabel via1 14309 12750 14309 12750 0 _081_
rlabel viali 12742 11186 12742 11186 0 _082_
rlabel metal1 13662 10982 13662 10982 0 _083_
rlabel metal1 13846 12648 13846 12648 0 _084_
rlabel metal2 13754 12682 13754 12682 0 _085_
rlabel metal2 14214 12959 14214 12959 0 _086_
rlabel metal1 13662 12954 13662 12954 0 _087_
rlabel metal1 13156 14042 13156 14042 0 _088_
rlabel metal1 13248 14586 13248 14586 0 _089_
rlabel metal1 13524 13838 13524 13838 0 _090_
rlabel metal2 13018 13056 13018 13056 0 _091_
rlabel metal1 13524 13498 13524 13498 0 _092_
rlabel metal1 9614 6222 9614 6222 0 _093_
rlabel metal1 4370 6392 4370 6392 0 _094_
rlabel metal1 8326 6358 8326 6358 0 _095_
rlabel metal1 8418 5746 8418 5746 0 _096_
rlabel metal2 6026 6052 6026 6052 0 _097_
rlabel metal1 6072 5610 6072 5610 0 _098_
rlabel metal1 6854 6222 6854 6222 0 _099_
rlabel metal2 5750 5916 5750 5916 0 _100_
rlabel metal2 4554 6324 4554 6324 0 _101_
rlabel metal1 6578 6766 6578 6766 0 _102_
rlabel metal1 7360 6834 7360 6834 0 _103_
rlabel metal1 5474 6766 5474 6766 0 _104_
rlabel metal1 4048 5678 4048 5678 0 _105_
rlabel metal1 4416 6290 4416 6290 0 _106_
rlabel metal1 4370 6630 4370 6630 0 _107_
rlabel metal1 4002 5780 4002 5780 0 _108_
rlabel metal1 3450 6630 3450 6630 0 _109_
rlabel metal1 2852 6222 2852 6222 0 _110_
rlabel metal2 3450 8160 3450 8160 0 _111_
rlabel metal1 4278 9010 4278 9010 0 _112_
rlabel metal1 4784 7718 4784 7718 0 _113_
rlabel metal1 3772 8398 3772 8398 0 _114_
rlabel metal1 3772 9146 3772 9146 0 _115_
rlabel metal2 4830 7956 4830 7956 0 _116_
rlabel metal2 5290 9044 5290 9044 0 _117_
rlabel metal2 4922 9350 4922 9350 0 _118_
rlabel metal1 3266 9078 3266 9078 0 _119_
rlabel metal1 6348 10506 6348 10506 0 _120_
rlabel metal1 5290 10540 5290 10540 0 _121_
rlabel metal1 6348 10574 6348 10574 0 _122_
rlabel metal1 6486 10778 6486 10778 0 _123_
rlabel metal1 5152 10982 5152 10982 0 _124_
rlabel metal1 4784 10778 4784 10778 0 _125_
rlabel via2 4554 11101 4554 11101 0 _126_
rlabel metal1 4048 11322 4048 11322 0 _127_
rlabel metal1 2668 10438 2668 10438 0 _128_
rlabel metal1 3726 11084 3726 11084 0 _129_
rlabel metal1 2622 10608 2622 10608 0 _130_
rlabel metal1 4695 11322 4695 11322 0 _131_
rlabel metal1 4884 9350 4884 9350 0 _132_
rlabel metal1 5060 9554 5060 9554 0 _133_
rlabel metal1 2530 11696 2530 11696 0 _134_
rlabel metal1 7038 9384 7038 9384 0 _135_
rlabel metal1 8142 9554 8142 9554 0 _136_
rlabel metal1 6946 9520 6946 9520 0 _137_
rlabel metal1 6532 8398 6532 8398 0 _138_
rlabel metal1 6394 8602 6394 8602 0 _139_
rlabel metal1 9062 8534 9062 8534 0 _140_
rlabel metal1 10764 9010 10764 9010 0 _141_
rlabel metal1 7866 7276 7866 7276 0 _142_
rlabel metal2 9982 8942 9982 8942 0 _143_
rlabel metal1 9154 9044 9154 9044 0 _144_
rlabel metal1 9890 9044 9890 9044 0 _145_
rlabel metal2 10902 9180 10902 9180 0 _146_
rlabel metal1 12098 9010 12098 9010 0 _147_
rlabel metal2 9982 13600 9982 13600 0 _148_
rlabel metal1 3588 14314 3588 14314 0 _149_
rlabel metal1 6256 13702 6256 13702 0 _150_
rlabel metal1 5888 14586 5888 14586 0 _151_
rlabel metal1 8280 13498 8280 13498 0 _152_
rlabel metal1 9016 13906 9016 13906 0 _153_
rlabel metal1 9568 13906 9568 13906 0 _154_
rlabel metal1 9154 12070 9154 12070 0 _155_
rlabel metal1 10028 12410 10028 12410 0 _156_
rlabel metal1 11224 12410 11224 12410 0 _157_
rlabel metal2 11362 14348 11362 14348 0 _158_
rlabel metal2 6302 12070 6302 12070 0 _159_
rlabel metal1 5980 12342 5980 12342 0 _160_
rlabel metal2 5658 12036 5658 12036 0 _161_
rlabel metal2 874 14052 874 14052 0 clk
rlabel metal1 5014 10608 5014 10608 0 clknet_0_clk
rlabel metal2 1426 6595 1426 6595 0 clknet_2_0__leaf_clk
rlabel metal1 4048 10778 4048 10778 0 clknet_2_1__leaf_clk
rlabel metal1 9246 5134 9246 5134 0 clknet_2_2__leaf_clk
rlabel metal1 10350 14484 10350 14484 0 clknet_2_3__leaf_clk
rlabel metal1 10488 5678 10488 5678 0 counter\[0\]
rlabel metal1 2760 11118 2760 11118 0 counter\[10\]
rlabel metal1 4462 11832 4462 11832 0 counter\[11\]
rlabel metal2 9062 8976 9062 8976 0 counter\[12\]
rlabel metal1 10166 11594 10166 11594 0 counter\[13\]
rlabel metal1 10534 11186 10534 11186 0 counter\[14\]
rlabel metal1 11638 10098 11638 10098 0 counter\[15\]
rlabel metal1 6808 5338 6808 5338 0 counter\[1\]
rlabel metal1 6348 5338 6348 5338 0 counter\[2\]
rlabel metal1 6624 7446 6624 7446 0 counter\[3\]
rlabel metal2 4738 8092 4738 8092 0 counter\[4\]
rlabel metal1 2944 6970 2944 6970 0 counter\[5\]
rlabel metal2 2898 8772 2898 8772 0 counter\[6\]
rlabel metal1 4094 9452 4094 9452 0 counter\[7\]
rlabel metal1 5336 11594 5336 11594 0 counter\[8\]
rlabel metal1 4784 12614 4784 12614 0 counter\[9\]
rlabel metal1 6486 14960 6486 14960 0 data[0]
rlabel metal1 7360 14926 7360 14926 0 data[1]
rlabel metal1 9246 14892 9246 14892 0 data[2]
rlabel metal1 10258 14960 10258 14960 0 data[3]
rlabel metal1 12006 14994 12006 14994 0 data[4]
rlabel metal1 12512 14926 12512 14926 0 data[5]
rlabel metal1 13800 14926 13800 14926 0 data[6]
rlabel metal2 15042 15310 15042 15310 0 data[7]
rlabel metal1 5750 14246 5750 14246 0 divider\[0\]
rlabel metal2 6394 14450 6394 14450 0 divider\[1\]
rlabel metal1 8234 12274 8234 12274 0 divider\[2\]
rlabel metal1 7728 14586 7728 14586 0 divider\[3\]
rlabel metal1 9568 14586 9568 14586 0 divider\[4\]
rlabel metal1 9016 12614 9016 12614 0 divider\[5\]
rlabel metal1 10810 11798 10810 11798 0 divider\[6\]
rlabel metal2 11914 11492 11914 11492 0 divider\[7\]
rlabel metal1 3542 14926 3542 14926 0 ext_data
rlabel metal1 4830 14926 4830 14926 0 load_divider
rlabel metal1 2300 14926 2300 14926 0 n_rst
rlabel metal2 5750 13396 5750 13396 0 net1
rlabel metal1 6348 14450 6348 14450 0 net10
rlabel metal1 2668 13838 2668 13838 0 net11
rlabel metal1 2116 14518 2116 14518 0 net12
rlabel metal1 2162 7922 2162 7922 0 net13
rlabel metal1 4416 5746 4416 5746 0 net14
rlabel metal2 2714 10778 2714 10778 0 net15
rlabel metal1 7958 7344 7958 7344 0 net16
rlabel metal1 7452 5882 7452 5882 0 net17
rlabel metal1 4738 9010 4738 9010 0 net18
rlabel metal1 10994 9520 10994 9520 0 net19
rlabel metal2 7590 14246 7590 14246 0 net2
rlabel metal1 9936 5882 9936 5882 0 net20
rlabel metal1 13386 6222 13386 6222 0 net21
rlabel metal1 13294 13294 13294 13294 0 net22
rlabel metal2 5566 11628 5566 11628 0 net23
rlabel metal1 9430 8976 9430 8976 0 net24
rlabel metal1 7774 13260 7774 13260 0 net3
rlabel metal2 10442 11424 10442 11424 0 net4
rlabel metal1 10074 13940 10074 13940 0 net5
rlabel metal1 9890 13430 9890 13430 0 net6
rlabel metal1 14214 13294 14214 13294 0 net7
rlabel via1 12821 14450 12821 14450 0 net8
rlabel metal1 4416 14858 4416 14858 0 net9
rlabel metal3 13133 1292 13133 1292 0 r2r_out[0]
rlabel metal1 12282 6970 12282 6970 0 r2r_out[1]
rlabel metal1 12926 6936 12926 6936 0 r2r_out[2]
rlabel metal1 13846 7344 13846 7344 0 r2r_out[3]
rlabel metal1 14996 8806 14996 8806 0 r2r_out[4]
rlabel metal2 14950 10829 14950 10829 0 r2r_out[5]
rlabel via2 15042 12325 15042 12325 0 r2r_out[6]
rlabel via2 15042 14467 15042 14467 0 r2r_out[7]
rlabel metal1 3542 14552 3542 14552 0 rst
<< properties >>
string FIXED_BBOX 0 0 16000 16000
<< end >>
