magic
tech sky130A
magscale 1 2
timestamp 1708461036
<< metal1 >>
rect 160 1880 360 2080
rect 480 1880 680 2080
rect 780 1880 980 2080
rect 1100 1880 1300 2080
rect 1420 1880 1620 2080
rect 1740 1880 1940 2080
rect 2060 1880 2260 2080
rect 2400 2002 2600 2080
rect 2398 1880 2600 2002
rect 274 1622 334 1880
rect 568 1754 628 1880
rect 910 1830 970 1880
rect 910 1770 1068 1830
rect 568 1694 868 1754
rect 274 1562 664 1622
rect 808 1568 868 1694
rect 1008 1562 1068 1770
rect 1206 1586 1266 1880
rect 1466 1792 1526 1880
rect 1758 1848 1818 1880
rect 1406 1732 1526 1792
rect 1664 1788 1818 1848
rect 2098 1842 2158 1880
rect 1664 1764 1724 1788
rect 1406 1584 1466 1732
rect 1612 1704 1724 1764
rect 1928 1782 2158 1842
rect 1928 1756 1988 1782
rect 1612 1586 1672 1704
rect 1810 1696 1988 1756
rect 1810 1592 1870 1696
rect 2398 1650 2458 1880
rect 2000 1590 2458 1650
rect 784 802 952 804
rect 610 344 670 802
rect 784 600 968 802
rect 592 188 876 344
rect 280 -462 480 -400
rect 906 -424 968 600
rect 1004 350 1074 794
rect 1208 628 1362 832
rect 1000 194 1284 350
rect 806 -430 968 -424
rect 1312 -426 1362 628
rect 1404 366 1474 810
rect 1598 642 1766 846
rect 1702 636 1764 642
rect 1394 210 1652 366
rect 1710 -418 1764 636
rect 1804 368 1874 814
rect 1988 668 2072 770
rect 1988 560 2306 668
rect 1988 462 2500 560
rect 2002 460 2500 462
rect 2156 396 2500 460
rect 1794 212 2078 368
rect 1604 -420 1652 -418
rect 1710 -420 1870 -418
rect 1312 -428 1374 -426
rect 280 -552 656 -462
rect 280 -600 480 -552
rect 806 -570 1074 -430
rect 1206 -568 1472 -428
rect 1604 -558 1870 -420
rect 2166 -422 2252 396
rect 2300 360 2500 396
rect 1996 -562 2262 -422
rect 806 -584 956 -570
use sky130_fd_pr__res_high_po_0p35_JK9DHS  XR1
timestamp 1708459662
transform 1 0 637 0 1 1132
box -37 -532 37 532
use sky130_fd_pr__res_high_po_0p35_JK9DHS  XR2
timestamp 1708459662
transform 1 0 837 0 1 1132
box -37 -532 37 532
use sky130_fd_pr__res_high_po_0p35_JK9DHS  XR3
timestamp 1708459662
transform 1 0 1037 0 1 1132
box -37 -532 37 532
use sky130_fd_pr__res_high_po_0p35_JK9DHS  XR4
timestamp 1708459662
transform 1 0 1237 0 1 1132
box -37 -532 37 532
use sky130_fd_pr__res_high_po_0p35_JK9DHS  XR5
timestamp 1708459662
transform 1 0 1437 0 1 1132
box -37 -532 37 532
use sky130_fd_pr__res_high_po_0p35_JK9DHS  XR6
timestamp 1708459662
transform 1 0 1637 0 1 1132
box -37 -532 37 532
use sky130_fd_pr__res_high_po_0p35_JK9DHS  XR7
timestamp 1708459662
transform 1 0 1837 0 1 1132
box -37 -532 37 532
use sky130_fd_pr__res_high_po_0p35_JK9DHS  XR8
timestamp 1708459662
transform 1 0 2037 0 1 1132
box -37 -532 37 532
use sky130_fd_pr__res_high_po_0p35_B8JXJA  XR9
timestamp 1708459662
transform 1 0 837 0 1 -118
box -37 -482 37 482
use sky130_fd_pr__res_high_po_0p35_B8JXJA  XR10
timestamp 1708459662
transform 1 0 1037 0 1 -118
box -37 -482 37 482
use sky130_fd_pr__res_high_po_0p35_B8JXJA  XR11
timestamp 1708459662
transform 1 0 1237 0 1 -118
box -37 -482 37 482
use sky130_fd_pr__res_high_po_0p35_B8JXJA  XR12
timestamp 1708459662
transform 1 0 1437 0 1 -118
box -37 -482 37 482
use sky130_fd_pr__res_high_po_0p35_B8JXJA  XR13
timestamp 1708459662
transform 1 0 1637 0 1 -118
box -37 -482 37 482
use sky130_fd_pr__res_high_po_0p35_B8JXJA  XR14
timestamp 1708459662
transform 1 0 1837 0 1 -118
box -37 -482 37 482
use sky130_fd_pr__res_high_po_0p35_B8JXJA  sky130_fd_pr__res_high_po_0p35_B8JXJA_0
timestamp 1708459662
transform 1 0 2037 0 1 -118
box -37 -482 37 482
use sky130_fd_pr__res_high_po_0p35_JK9DHS  sky130_fd_pr__res_high_po_0p35_JK9DHS_0
timestamp 1708459662
transform 1 0 637 0 1 -68
box -37 -532 37 532
<< labels >>
flabel metal1 480 1880 680 2080 0 FreeSans 256 0 0 0 b1
port 1 nsew
flabel metal1 160 1880 360 2080 0 FreeSans 256 0 0 0 b0
port 0 nsew
flabel metal1 780 1880 980 2080 0 FreeSans 256 0 0 0 b2
port 2 nsew
flabel metal1 1100 1880 1300 2080 0 FreeSans 256 0 0 0 b3
port 3 nsew
flabel metal1 1420 1880 1620 2080 0 FreeSans 256 0 0 0 b4
port 4 nsew
flabel metal1 1740 1880 1940 2080 0 FreeSans 256 0 0 0 b5
port 5 nsew
flabel metal1 2060 1880 2260 2080 0 FreeSans 256 0 0 0 b6
port 6 nsew
flabel metal1 2400 1880 2600 2080 0 FreeSans 256 0 0 0 b7
port 7 nsew
flabel metal1 2300 360 2500 560 0 FreeSans 256 0 0 0 out
port 8 nsew
flabel metal1 280 -600 480 -400 0 FreeSans 256 0 0 0 B
port 9 nsew
<< end >>
