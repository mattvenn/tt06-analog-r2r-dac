** sch_path: /home/matt/work/asic-workshop/shuttle-2404/tt06-analog-r2r-dac/xschem/r2r.sch
.subckt r2r b0 b1 b2 b3 b4 b5 b6 b7 out VSUBS GND
*.PININFO b0:I b1:I b2:I b3:I b4:I b5:I b6:I b7:I out:O VSUBS:I GND:B
XR1 net1 b0 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR2 net2 b1 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR3 net3 b2 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR4 net4 b3 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR5 net5 b4 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR6 net6 b5 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR7 net7 b6 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR8 out b7 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR9 net2 net1 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR10 net3 net2 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR11 net4 net3 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR12 net5 net4 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR13 net6 net5 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR14 net7 net6 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR15 out net7 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR16 GND net1 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
.ends
.end
