magic
tech sky130A
magscale 1 2
timestamp 1709129632
<< pwell >>
rect -2480 2660 -1760 2740
<< metal1 >>
rect -1200 17400 -960 17600
rect -600 17400 -360 17600
rect 0 17400 240 17600
rect 600 17400 840 17600
rect 1200 17400 1440 17600
rect 1800 17400 2040 17600
rect 2400 17400 2640 17600
rect 3000 17400 3240 17600
rect -1040 16460 -960 17400
rect -440 16460 -360 17400
rect 160 16460 240 17400
rect 760 16460 840 17400
rect 1360 16460 1440 17400
rect 1960 16460 2040 17400
rect 2560 16460 2640 17400
rect 3160 16460 3240 17400
rect -1840 11620 -1380 11700
rect -1840 11060 -1760 11620
rect -1460 8200 -1380 11620
rect -1460 8120 -960 8200
rect -1040 7040 -960 8120
rect -740 8120 -360 8200
rect -2600 2740 -2400 2800
rect -1840 2740 -1760 2920
rect -740 2740 -660 8120
rect 160 7260 240 8200
rect -440 7180 240 7260
rect 160 7040 240 7180
rect 460 8120 840 8200
rect 460 2740 540 8120
rect 1360 7260 1440 8200
rect 760 7180 1440 7260
rect 1360 7040 1440 7180
rect 1660 8120 2040 8200
rect 1660 2740 1740 8120
rect 2560 7260 2640 8220
rect 1960 7180 2640 7260
rect 2560 7060 2640 7180
rect 3160 7540 3240 8220
rect 4000 8000 4200 8200
rect 4000 7540 4080 8000
rect 3160 7460 4080 7540
rect 2560 2760 2640 2900
rect 3160 2760 3240 7460
rect -2600 2660 -1760 2740
rect -1040 2660 -360 2740
rect 160 2660 840 2740
rect 1360 2660 2040 2740
rect 2560 2680 3240 2760
rect -2600 2600 -2400 2660
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR1
timestamp 1709128825
transform 1 0 -999 0 1 12398
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR2
timestamp 1709128825
transform 1 0 -399 0 1 12398
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR3
timestamp 1709128825
transform 1 0 201 0 1 12398
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR4
timestamp 1709128825
transform 1 0 801 0 1 12398
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR5
timestamp 1709128825
transform 1 0 1401 0 1 12398
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR6
timestamp 1709128825
transform 1 0 2001 0 1 12398
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR7
timestamp 1709128825
transform 1 0 2601 0 1 12398
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR8
timestamp 1709128825
transform 1 0 3201 0 1 12398
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR9
timestamp 1709128825
transform 1 0 -999 0 1 4998
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR10
timestamp 1709128825
transform 1 0 -399 0 1 4998
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR11
timestamp 1709128825
transform 1 0 201 0 1 4998
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR12
timestamp 1709128825
transform 1 0 801 0 1 4998
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR13
timestamp 1709128825
transform 1 0 1401 0 1 4998
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR14
timestamp 1709128825
transform 1 0 2001 0 1 4998
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR15
timestamp 1709128825
transform 1 0 2601 0 1 4998
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR16
timestamp 1709128825
transform 1 0 -1799 0 1 6998
box -201 -4598 201 4598
<< labels >>
flabel metal1 4000 8000 4200 8200 0 FreeSans 256 0 0 0 out
port 8 nsew
flabel metal1 -600 17400 -400 17600 0 FreeSans 256 0 0 0 b1
port 1 nsew
flabel metal1 0 17400 200 17600 0 FreeSans 256 0 0 0 b2
port 2 nsew
flabel metal1 600 17400 800 17600 0 FreeSans 256 0 0 0 b3
port 3 nsew
flabel metal1 1200 17400 1400 17600 0 FreeSans 256 0 0 0 b4
port 4 nsew
flabel metal1 1800 17400 2000 17600 0 FreeSans 256 0 0 0 b5
port 5 nsew
flabel metal1 2400 17400 2600 17600 0 FreeSans 256 0 0 0 b6
port 6 nsew
flabel metal1 3000 17400 3200 17600 0 FreeSans 256 0 0 0 b7
port 7 nsew
flabel metal1 -1200 17400 -1000 17600 0 FreeSans 256 0 0 0 b0
port 0 nsew
flabel metal1 -2600 2600 -2400 2800 0 FreeSans 256 0 0 0 GND
port 10 nsew
<< end >>
