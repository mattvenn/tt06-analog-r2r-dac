** sch_path: /home/matt/work/asic-workshop/shuttle-2404/tt06-analog-r2r-dac/xschem/testbench.sch
**.subckt testbench
x1 b0 b1 b2 b3 out r2r
V1 b3 GND pulse(0 1.8 0 0 0 8u 16u)
V2 b2 GND pulse(0 1.8 0 0 0 4u 8u)
V3 b1 GND pulse(0 1.8 0 0 0 2u 4u)
V4 b0 GND pulse(0 1.8 0 0 0 1u 2u)
**** begin user architecture code


.tran 1n 20u uic
.save all


**** end user architecture code
**.ends

* expanding   symbol:  r2r.sym # of pins=5
** sym_path: /home/matt/work/asic-workshop/shuttle-2404/tt06-analog-r2r-dac/xschem/r2r.sym
** sch_path: /home/matt/work/asic-workshop/shuttle-2404/tt06-analog-r2r-dac/xschem/r2r.sch
.subckt r2r b0 b1 b2 b3 out
*.ipin b1
*.opin out
*.ipin b0
*.ipin b2
*.ipin b3
R1 b0 net1 1k m=1
R2 b1 net2 1k m=1
R3 b2 net3 1k m=1
R4 net1 GND 1k m=1
R5 b3 out 1k m=1
R6 net2 net1 500 m=1
R7 net3 net2 500 m=1
R8 out net3 500 m=1
.ends

.GLOBAL GND
.end
