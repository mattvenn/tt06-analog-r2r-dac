* NGSPICE file created from tt_um_mattvenn_r2r_dac.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X a_78_199# a_215_47#
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.141375 ps=1.41 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=2.003333 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=10400,504
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
**devattr s=9400,294 d=4200,242
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=2.003333 as=0.28 ps=2.56 w=1 l=0.15
**devattr s=11200,512 d=14900,349
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.141375 ps=1.41 w=0.65 l=0.15
**devattr s=4550,200 d=3510,184
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
**devattr s=4700,247 d=9400,294
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.141375 pd=1.41 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.141375 pd=1.41 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=4550,200
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.335 ps=2.003333 w=1 l=0.15
**devattr s=14900,349 d=4700,247
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
C0 B2 VGND 0.010267f
C1 B2 a_78_199# 0.081601f
C2 A1 VPB 0.031899f
C3 a_78_199# VPB 0.05169f
C4 B2 a_215_47# 0.020719f
C5 B1 VGND 0.011856f
C6 a_78_199# B1 0.147802f
C7 A1 VPWR 0.05704f
C8 VGND VPWR 0.066763f
C9 a_78_199# VPWR 0.211049f
C10 a_493_297# A2 0.010465f
C11 B2 VPB 0.028066f
C12 a_78_199# a_292_297# 0.012951f
C13 B2 B1 0.081466f
C14 B1 VPB 0.038762f
C15 A1 A2 0.087859f
C16 A2 VGND 0.015286f
C17 B2 VPWR 0.010367f
C18 a_78_199# A2 0.070688f
C19 VPWR VPB 0.074428f
C20 X VGND 0.047175f
C21 a_78_199# X 0.104588f
C22 A2 a_215_47# 0.043898f
C23 B1 VPWR 0.022722f
C24 B2 A2 0.06759f
C25 A2 VPB 0.034104f
C26 X VPB 0.010691f
C27 A1 VGND 0.014626f
C28 A2 VPWR 0.120404f
C29 a_78_199# VGND 0.068403f
C30 A1 a_215_47# 0.049793f
C31 X VPWR 0.091108f
C32 VGND a_215_47# 0.257828f
C33 a_78_199# a_215_47# 0.090715f
C34 VGND VNB 0.402531f
C35 VPWR VNB 0.35911f
C36 X VNB 0.088397f
C37 A1 VNB 0.132282f
C38 A2 VNB 0.097054f
C39 B2 VNB 0.091305f
C40 B1 VNB 0.109674f
C41 VPB VNB 0.69336f
C42 a_215_47# VNB 0.035725f
C43 a_78_199# VNB 0.15408f
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=4.73
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=4.73
**devattr d=5720,324
C0 VPWR VGND 1.56539f
C1 VPB VGND 0.349732f
C2 VPWR VPB 0.136888f
C3 VPWR VNB 1.67352f
C4 VGND VNB 1.46552f
C5 VPB VNB 1.13634f
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q a_891_413# a_466_413# a_1059_315#
+ a_193_47# a_634_159# a_381_47# a_27_47#
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12054 ps=1.304827 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12353 pd=1.162647 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.193015 ps=1.816635 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.081066 ps=0.762987 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.077887 pd=0.843119 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193015 pd=1.816635 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.081066 pd=0.762987 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0.118685 ps=1.284752 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0.144761 ps=1.362476 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.077887 pd=0.843119 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.077887 ps=0.843119 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.081066 pd=0.762987 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.12353 ps=1.162647 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.12054 pd=1.304827 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0.077887 ps=0.843119 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.077887 pd=0.843119 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
C0 a_193_47# a_381_47# 0.101638f
C1 D VGND 0.038993f
C2 VPWR CLK 0.019411f
C3 VPB D 0.096334f
C4 a_891_413# VGND 0.131537f
C5 VPB a_891_413# 0.069773f
C6 a_466_413# a_27_47# 0.273138f
C7 a_27_47# a_381_47# 0.062224f
C8 VPWR a_193_47# 0.117215f
C9 Q a_1059_315# 0.081249f
C10 D a_381_47# 0.112186f
C11 a_27_47# CLK 0.213838f
C12 VPWR a_27_47# 0.379856f
C13 a_634_159# VGND 0.124877f
C14 VPB a_634_159# 0.07647f
C15 a_193_47# a_27_47# 0.974525f
C16 a_1059_315# VGND 0.155119f
C17 VPB a_1059_315# 0.154738f
C18 VPWR D 0.025067f
C19 Q VGND 0.076612f
C20 VPWR a_891_413# 0.115323f
C21 Q VPB 0.013828f
C22 a_466_413# a_634_159# 0.239923f
C23 a_193_47# D 0.175777f
C24 a_193_47# a_891_413# 0.196846f
C25 D a_27_47# 0.065857f
C26 VPB VGND 0.012227f
C27 a_27_47# a_891_413# 0.032244f
C28 VPWR a_634_159# 0.102126f
C29 a_193_47# a_634_159# 0.127288f
C30 VPWR a_1059_315# 0.232446f
C31 a_466_413# VGND 0.088802f
C32 a_466_413# VPB 0.074456f
C33 VPWR Q 0.110929f
C34 a_381_47# VGND 0.052221f
C35 VPB a_381_47# 0.014142f
C36 a_193_47# a_1059_315# 0.034054f
C37 a_634_159# a_27_47# 0.141453f
C38 VGND CLK 0.019463f
C39 VPB CLK 0.070057f
C40 a_466_413# a_381_47# 0.037333f
C41 a_1059_315# a_27_47# 0.048748f
C42 VPWR VGND 0.063886f
C43 VPWR VPB 0.168181f
C44 a_634_159# a_891_413# 0.036838f
C45 a_193_47# VGND 0.200101f
C46 a_193_47# VPB 0.176133f
C47 a_1059_315# a_891_413# 0.310858f
C48 VPWR a_466_413# 0.170985f
C49 VPWR a_381_47# 0.061283f
C50 a_27_47# VGND 0.136686f
C51 VPB a_27_47# 0.247821f
C52 a_466_413# a_193_47# 0.083013f
C53 Q VNB 0.088256f
C54 VGND VNB 0.84362f
C55 VPWR VNB 0.681368f
C56 D VNB 0.142509f
C57 CLK VNB 0.195983f
C58 VPB VNB 1.49072f
C59 a_381_47# VNB 0.015369f
C60 a_891_413# VNB 0.161052f
C61 a_1059_315# VNB 0.248849f
C62 a_466_413# VNB 0.133203f
C63 a_634_159# VNB 0.142309f
C64 a_193_47# VNB 0.284262f
C65 a_27_47# VNB 0.449511f
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
C0 VPWR VGND 0.042274f
C1 Y A 0.089386f
C2 VPB VPWR 0.052063f
C3 VPWR A 0.06305f
C4 Y VPWR 0.209105f
C5 VGND A 0.063754f
C6 VPB A 0.074183f
C7 Y VGND 0.154601f
C8 VGND VNB 0.266187f
C9 Y VNB 0.03316f
C10 VPWR VNB 0.246044f
C11 A VNB 0.262807f
C12 VPB VNB 0.338976f
.ends

.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X a_227_47# a_77_199#
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.1313 ps=1.184 w=0.65 l=0.15
**devattr s=5070,208 d=5330,212
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=7800,278
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.186667 ps=1.706667 w=1 l=0.15
**devattr s=5400,254 d=6600,266
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1313 pd=1.184 as=0.13325 ps=1.06 w=0.65 l=0.15
**devattr s=5330,212 d=7540,376
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186667 pd=1.706667 as=0.205 ps=1.41 w=1 l=0.15
**devattr s=8200,282 d=11600,516
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1313 pd=1.184 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=5070,208 d=5070,208
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186667 pd=1.706667 as=0.335 ps=2.67 w=1 l=0.15
**devattr s=13400,534 d=5400,254
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
**devattr s=7800,278 d=7800,278
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1313 ps=1.184 w=0.65 l=0.15
**devattr s=4290,196 d=5070,208
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1313 pd=1.184 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=3510,184 d=4290,196
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
**devattr s=7800,278 d=8200,282
C0 A2 A1 0.075092f
C1 B2 VPWR 0.012246f
C2 X VPWR 0.102456f
C3 a_227_47# VGND 0.326249f
C4 A1 VPWR 0.018718f
C5 VPB A3 0.033035f
C6 A2 a_323_297# 0.011623f
C7 a_227_297# a_77_199# 0.018661f
C8 A2 VGND 0.016397f
C9 a_227_47# A2 0.041255f
C10 B2 B1 0.04397f
C11 VGND VPWR 0.072113f
C12 B2 a_77_199# 0.116444f
C13 a_77_199# X 0.092774f
C14 A2 VPWR 0.013495f
C15 A1 a_77_199# 0.123952f
C16 VGND B1 0.010652f
C17 a_227_47# B1 0.03409f
C18 a_77_199# a_323_297# 0.014272f
C19 B2 A3 0.102249f
C20 VGND a_77_199# 0.038735f
C21 a_227_47# a_77_199# 0.085098f
C22 A2 a_77_199# 0.113015f
C23 B1 VPWR 0.046731f
C24 B2 VPB 0.033813f
C25 VPB X 0.015707f
C26 a_77_199# VPWR 0.360105f
C27 VPB A1 0.029013f
C28 VGND A3 0.013109f
C29 a_227_47# A3 0.037584f
C30 A2 A3 0.106179f
C31 a_539_297# a_77_199# 0.022925f
C32 a_77_199# B1 0.046787f
C33 A2 VPB 0.033537f
C34 VPB VPWR 0.083235f
C35 A3 a_77_199# 0.030617f
C36 B2 VGND 0.010524f
C37 VPB B1 0.041119f
C38 a_227_47# B2 0.027482f
C39 VGND X 0.103165f
C40 VPB a_77_199# 0.047656f
C41 VGND A1 0.019687f
C42 a_227_47# A1 0.015082f
C43 VGND VNB 0.437857f
C44 VPWR VNB 0.404492f
C45 X VNB 0.100953f
C46 B1 VNB 0.150231f
C47 B2 VNB 0.097709f
C48 A3 VNB 0.096505f
C49 A2 VNB 0.096218f
C50 A1 VNB 0.094556f
C51 VPB VNB 0.781956f
C52 a_227_47# VNB 0.030865f
C53 a_77_199# VNB 0.146762f
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=0.59
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=0.59
**devattr d=5720,324
C0 VGND VPWR 0.352999f
C1 VGND VPB 0.079664f
C2 VPB VPWR 0.062496f
C3 VPWR VNB 0.469966f
C4 VGND VNB 0.427318f
C5 VPB VNB 0.338976f
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=1.05
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=1.05
**devattr d=5720,324
C0 VGND VPWR 0.545943f
C1 VGND VPB 0.116247f
C2 VPB VPWR 0.078686f
C3 VPWR VNB 0.61942f
C4 VGND VNB 0.553666f
C5 VPB VNB 0.427572f
.ends

.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X a_215_297# a_27_413#
+ a_298_297#
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178333 pd=1.69 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=5400,254
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.216269 ps=1.395992 w=0.65 l=0.15
**devattr s=5436,220 d=3510,184
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178333 pd=1.69 as=0.189825 ps=1.883041 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.216269 ps=1.395992 w=0.65 l=0.15
**devattr s=10335,289 d=6760,364
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.079726 pd=0.790877 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.189825 ps=1.883041 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3640,186
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.139743 pd=0.902025 as=0.1113 ps=1.37 w=0.42 l=0.15
**devattr s=4452,274 d=5436,220
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.189825 pd=1.883041 as=0.178333 ps=1.69 w=1 l=0.15
**devattr s=5400,254 d=5600,256
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.216269 pd=1.395992 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=10335,289
C0 a_27_413# A1 0.057273f
C1 B1_N VGND 0.049226f
C2 a_298_297# VPWR 0.196264f
C3 A1 VPB 0.027656f
C4 a_27_413# VGND 0.098153f
C5 A1 VPWR 0.021516f
C6 a_27_413# B1_N 0.237073f
C7 VPB VGND 0.011706f
C8 B1_N VPB 0.103238f
C9 VPWR VGND 0.07888f
C10 B1_N VPWR 0.018972f
C11 a_27_413# VPB 0.098696f
C12 a_27_413# VPWR 0.107226f
C13 a_298_297# A2 0.035704f
C14 X VGND 0.057294f
C15 VPWR VPB 0.097622f
C16 a_298_297# a_215_297# 0.071778f
C17 A2 A1 0.111772f
C18 A1 a_215_297# 0.092984f
C19 A2 VGND 0.019667f
C20 a_215_297# VGND 0.271787f
C21 X VPB 0.011733f
C22 VPWR X 0.114913f
C23 a_27_413# a_215_297# 0.141213f
C24 A2 VPB 0.041742f
C25 a_215_297# VPB 0.05456f
C26 A2 VPWR 0.030697f
C27 a_215_297# VPWR 0.129868f
C28 a_298_297# A1 0.049414f
C29 a_215_297# a_382_47# 0.01048f
C30 a_215_297# X 0.080241f
C31 A1 VGND 0.01436f
C32 A2 a_215_297# 0.094911f
C33 VGND VNB 0.439582f
C34 X VNB 0.089001f
C35 VPWR VNB 0.36562f
C36 A2 VNB 0.107548f
C37 A1 VNB 0.089279f
C38 B1_N VNB 0.290462f
C39 VPB VNB 0.781956f
C40 a_215_297# VNB 0.152836f
C41 a_27_413# VNB 0.171579f
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.564 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=6600,266
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.07602 pd=0.866 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=4872,284
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.07602 pd=0.866 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.182 ps=1.564 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07602 ps=0.866 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07602 pd=0.866 as=0.1113 ps=1.37 w=0.42 l=0.15
**devattr s=4452,274 d=2814,151
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.564 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=12000,520
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07602 ps=0.866 w=0.42 l=0.15
**devattr s=2814,151 d=2352,140
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.182 ps=1.564 w=1 l=0.15
**devattr s=6600,266 d=5600,256
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.564 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
C0 VPWR A 0.021953f
C1 VGND a_27_47# 0.148483f
C2 VPB X 0.012159f
C3 a_27_47# X 0.327705f
C4 VGND X 0.21559f
C5 VPB A 0.032139f
C6 VPWR VPB 0.063172f
C7 a_27_47# A 0.195005f
C8 VPWR a_27_47# 0.219243f
C9 VGND A 0.043094f
C10 VPWR VGND 0.057043f
C11 X A 0.013951f
C12 VPWR X 0.316967f
C13 a_27_47# VPB 0.138763f
C14 VGND VNB 0.357713f
C15 X VNB 0.067008f
C16 VPWR VNB 0.307647f
C17 A VNB 0.147639f
C18 VPB VNB 0.604764f
C19 a_27_47# VNB 0.542977f
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=1.97
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=1.97
**devattr d=5720,324
C0 VPB VPWR 0.085759f
C1 VGND VPWR 0.903312f
C2 VPB VGND 0.161065f
C3 VPWR VNB 0.867393f
C4 VGND VNB 0.761362f
C5 VPB VNB 0.604764f
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=2.89
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=2.89
**devattr d=5720,324
C0 VPB VPWR 0.104823f
C1 VGND VPWR 1.27274f
C2 VPB VGND 0.219503f
C3 VPWR VNB 1.14152f
C4 VGND VNB 0.991595f
C5 VPB VNB 0.781956f
.ends

.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X a_516_297# a_85_193#
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19435 pd=1.378 as=0.082875 ps=0.905 w=0.65 l=0.15
**devattr s=3315,181 d=7540,376
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.19435 pd=1.378 as=0.143 ps=1.09 w=0.65 l=0.15
**devattr s=4030,192 d=4680,202
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
**devattr s=5000,250 d=7200,272
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0.19435 pd=1.378 as=0.2145 ps=1.96 w=0.65 l=0.15
**devattr s=8580,392 d=10985,299
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
**devattr s=15400,554 d=5000,250
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.283333 pd=1.9 as=0.18 ps=1.36 w=1 l=0.15
**devattr s=7200,272 d=11200,312
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.283333 pd=1.9 as=0.178333 ps=1.69 w=1 l=0.15
**devattr s=5400,254 d=11600,516
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.143 ps=1.09 w=0.65 l=0.15
**devattr s=7410,244 d=3315,181
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.19435 ps=1.378 w=0.65 l=0.15
**devattr s=10985,299 d=4030,192
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178333 pd=1.69 as=0.283333 ps=1.9 w=1 l=0.15
**devattr s=11200,312 d=5400,254
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.19435 ps=1.378 w=0.65 l=0.15
**devattr s=4680,202 d=7410,244
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178333 pd=1.69 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=10600,506
C0 C1 D1 0.169347f
C1 A1 VPWR 0.02157f
C2 VPB a_85_193# 0.066264f
C3 X VPWR 0.094258f
C4 D1 VPWR 0.036977f
C5 VPB B1 0.036936f
C6 C1 VGND 0.016422f
C7 VPWR a_516_297# 0.217239f
C8 A1 A2 0.083244f
C9 VGND VPWR 0.087252f
C10 C1 VPWR 0.04987f
C11 A2 a_516_297# 0.056021f
C12 VGND A2 0.046422f
C13 A1 a_85_193# 0.056088f
C14 a_85_193# X 0.106854f
C15 A1 B1 0.068882f
C16 a_85_193# D1 0.184988f
C17 C1 a_414_297# 0.01365f
C18 A2 VPWR 0.021508f
C19 A1 VPB 0.033363f
C20 a_85_193# VGND 0.292376f
C21 VPB X 0.010929f
C22 B1 a_516_297# 0.087957f
C23 VPB D1 0.038109f
C24 VGND B1 0.014558f
C25 C1 a_85_193# 0.037306f
C26 VPB a_516_297# 0.010413f
C27 C1 B1 0.164685f
C28 VPB VGND 0.0102f
C29 a_85_193# VPWR 0.14392f
C30 B1 VPWR 0.043795f
C31 C1 VPB 0.030173f
C32 VPB VPWR 0.098773f
C33 A1 a_516_297# 0.05885f
C34 VPB A2 0.033731f
C35 A1 VGND 0.116703f
C36 VGND X 0.068497f
C37 VGND D1 0.015289f
C38 a_85_193# B1 0.039821f
C39 VGND VNB 0.505453f
C40 VPWR VNB 0.405283f
C41 X VNB 0.088362f
C42 A2 VNB 0.136216f
C43 A1 VNB 0.114026f
C44 B1 VNB 0.101766f
C45 C1 VNB 0.09306f
C46 D1 VNB 0.10506f
C47 VPB VNB 0.870552f
C48 a_516_297# VNB 0.035006f
C49 a_85_193# VNB 0.166604f
.ends

.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X a_215_53# a_109_93#
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.076267 ps=0.849013 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.913333 as=0.076267 ps=0.849013 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.076267 pd=0.849013 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.076267 pd=0.849013 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.092605 pd=0.922174 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=5930,268
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2730,149
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.220489 ps=2.195652 w=1 l=0.15
**devattr s=5930,268 d=11000,510
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.092605 ps=0.922174 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.118032 ps=1.313948 w=0.65 l=0.15
**devattr s=4010,197 d=7150,370
C0 a_215_53# B 0.120778f
C1 VPWR VGND 0.06567f
C2 B VPB 0.110475f
C3 a_215_53# VGND 0.232049f
C4 B A 0.079275f
C5 a_215_53# VPWR 0.085727f
C6 VPB VGND 0.010346f
C7 VPWR VPB 0.109107f
C8 A VGND 0.018847f
C9 a_215_53# VPB 0.049294f
C10 a_215_53# A 0.245132f
C11 X VGND 0.035902f
C12 A VPB 0.03757f
C13 VPWR X 0.088522f
C14 B a_109_93# 0.099724f
C15 a_215_53# X 0.099129f
C16 C_N VGND 0.042739f
C17 C_N VPWR 0.037773f
C18 a_109_93# VGND 0.084353f
C19 X VPB 0.010957f
C20 VPWR a_109_93# 0.0369f
C21 a_215_53# a_109_93# 0.13675f
C22 C_N VPB 0.046442f
C23 a_109_93# VPB 0.053437f
C24 a_109_93# A 0.036898f
C25 B VGND 0.015735f
C26 VPWR B 0.234984f
C27 C_N a_109_93# 0.05842f
C28 VGND VNB 0.439259f
C29 X VNB 0.08839f
C30 A VNB 0.112741f
C31 C_N VNB 0.150085f
C32 B VNB 0.103426f
C33 VPWR VNB 0.362977f
C34 VPB VNB 0.69336f
C35 a_109_93# VNB 0.160708f
C36 a_215_53# VNB 0.142592f
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213258 pd=1.962121 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10600,506
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.213258 ps=1.962121 w=1 l=0.15
**devattr s=5960,265 d=5400,254
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.136485 pd=1.255758 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=5960,265
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.138408 ps=1.428488 w=0.65 l=0.15
**devattr s=3880,195 d=3510,184
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.138408 pd=1.428488 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6890,366
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.089433 pd=0.923023 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
C0 VPWR A 0.022108f
C1 VGND a_27_47# 0.12719f
C2 a_27_47# X 0.148785f
C3 VGND X 0.111264f
C4 VPB A 0.069727f
C5 VPWR VPB 0.05279f
C6 a_27_47# A 0.157874f
C7 VPWR a_27_47# 0.153302f
C8 VGND A 0.019887f
C9 VPWR VGND 0.051753f
C10 VPWR X 0.168994f
C11 a_27_47# VPB 0.074969f
C12 VGND VNB 0.284185f
C13 X VNB 0.021498f
C14 VPWR VNB 0.249629f
C15 A VNB 0.187471f
C16 VPB VNB 0.427572f
C17 a_27_47# VNB 0.28447f
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y a_47_47# a_285_47#
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.3475 ps=2.195 w=1 l=0.15
**devattr s=14600,346 d=4200,242
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3475 ps=2.195 w=1 l=0.15
**devattr s=12000,520 d=5400,254
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=2730,172
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=7800,380
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.06825 ps=0.86 w=0.65 l=0.15
**devattr s=2730,172 d=3510,184
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3475 pd=2.195 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=14600,346
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3475 pd=2.195 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=14400,544
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=6600,266
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
C0 VPWR A 0.034894f
C1 B a_47_47# 0.35554f
C2 a_47_47# VPB 0.044386f
C3 VGND a_47_47# 0.103529f
C4 B VPB 0.064326f
C5 VGND Y 0.038107f
C6 a_47_47# A 0.030704f
C7 VGND B 0.038916f
C8 a_47_47# a_285_47# 0.017546f
C9 Y a_285_47# 0.043869f
C10 B A 0.23582f
C11 VPWR a_47_47# 0.272937f
C12 B a_285_47# 0.066964f
C13 VPWR Y 0.107281f
C14 A VPB 0.082204f
C15 VPWR B 0.040822f
C16 VGND A 0.063473f
C17 VPWR VPB 0.071773f
C18 VGND a_285_47# 0.210545f
C19 A a_285_47# 0.035318f
C20 a_47_47# Y 0.142676f
C21 VGND VPWR 0.066517f
C22 VGND VNB 0.399812f
C23 Y VNB 0.078329f
C24 VPWR VNB 0.351939f
C25 A VNB 0.216579f
C26 B VNB 0.212328f
C27 VPB VNB 0.69336f
C28 a_285_47# VNB 0.017425f
C29 a_47_47# VNB 0.199276f
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X a_49_47# a_285_47# a_391_47#
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.073388 pd=0.748938 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.067596 pd=0.732251 as=0.1092 ps=1.36 w=0.42 l=0.5
**devattr s=4368,272 d=3880,195
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.174735 ps=1.783186 w=1 l=0.15
**devattr s=5630,265 d=10400,504
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.067596 pd=0.732251 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.073388 pd=0.748938 as=0.1092 ps=1.36 w=0.42 l=0.5
**devattr s=4368,272 d=5630,265
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.067596 ps=0.732251 w=0.42 l=0.5
**devattr s=2268,138 d=4368,272
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.073388 ps=0.748938 w=0.42 l=0.5
**devattr s=2268,138 d=4368,272
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.104613 ps=1.133246 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
C0 a_49_47# VPB 0.125413f
C1 VPB A 0.082837f
C2 a_49_47# VPWR 0.144268f
C3 VPWR A 0.020643f
C4 a_49_47# A 0.279977f
C5 a_391_47# VGND 0.130239f
C6 a_391_47# a_285_47# 0.419086f
C7 VGND X 0.07961f
C8 a_285_47# VPB 0.156427f
C9 VGND VPWR 0.071507f
C10 VPWR a_285_47# 0.119832f
C11 a_49_47# VGND 0.143546f
C12 a_49_47# a_285_47# 0.22264f
C13 VGND A 0.021393f
C14 a_391_47# VPB 0.044127f
C15 a_391_47# X 0.128943f
C16 X VPB 0.015496f
C17 a_391_47# VPWR 0.134775f
C18 VPWR VPB 0.0787f
C19 VPWR X 0.080229f
C20 VGND a_285_47# 0.120945f
C21 VGND VNB 0.43965f
C22 X VNB 0.095447f
C23 VPWR VNB 0.367348f
C24 A VNB 0.178652f
C25 VPB VNB 0.781956f
C26 a_391_47# VNB 0.127705f
C27 a_285_47# VNB 0.29867f
C28 a_49_47# VNB 0.306903f
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X a_193_297# a_109_297#
+ a_27_47#
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4290,196
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.191667 ps=1.716667 w=1 l=0.15
**devattr s=6300,263 d=10400,504
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.15 ps=1.3 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.104813 ps=0.9725 w=0.65 l=0.15
**devattr s=4095,193 d=6760,364
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.104813 ps=0.9725 w=0.65 l=0.15
**devattr s=4290,196 d=2730,172
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.191667 pd=1.716667 as=0.15 ps=1.3 w=1 l=0.15
**devattr s=6600,266 d=6300,263
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.191667 ps=1.716667 w=1 l=0.15
**devattr s=10400,504 d=6600,266
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
**devattr s=2730,172 d=6760,364
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104813 pd=0.9725 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4290,196
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104813 pd=0.9725 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=4095,193
C0 B2 C1 0.072571f
C1 VPB a_27_47# 0.05124f
C2 VPWR X 0.089708f
C3 VPB B1 0.032075f
C4 a_109_297# VPWR 0.150131f
C5 B2 VGND 0.017443f
C6 A1 A2 0.069236f
C7 VGND X 0.061021f
C8 VPWR A2 0.020928f
C9 A1 a_193_297# 0.010869f
C10 a_193_297# VPWR 0.169243f
C11 B2 a_109_297# 0.013349f
C12 VGND A2 0.016752f
C13 A1 a_27_47# 0.09838f
C14 a_27_47# VPWR 0.099007f
C15 A1 B1 0.060935f
C16 a_27_47# C1 0.07922f
C17 A1 VPB 0.034297f
C18 a_27_47# VGND 0.395423f
C19 VPB VPWR 0.079908f
C20 a_465_47# a_27_47# 0.013015f
C21 VPB C1 0.036702f
C22 VGND B1 0.013269f
C23 a_109_297# a_193_297# 0.092725f
C24 B2 a_27_47# 0.09593f
C25 B2 B1 0.078429f
C26 a_27_47# X 0.09209f
C27 a_27_47# a_109_297# 0.096132f
C28 B2 VPB 0.025561f
C29 VPB X 0.011274f
C30 a_27_47# A2 0.152957f
C31 A1 VPWR 0.01613f
C32 a_27_47# a_193_297# 0.143754f
C33 C1 VPWR 0.013943f
C34 A1 VGND 0.012567f
C35 VPB A2 0.026961f
C36 VGND VPWR 0.072225f
C37 VGND C1 0.019615f
C38 a_27_47# B1 0.11237f
C39 VGND VNB 0.437277f
C40 X VNB 0.091856f
C41 VPWR VNB 0.363959f
C42 A2 VNB 0.089572f
C43 A1 VNB 0.105908f
C44 B1 VNB 0.108471f
C45 B2 VNB 0.088691f
C46 C1 VNB 0.139233f
C47 VPB VNB 0.781956f
C48 a_27_47# VNB 0.216317f
.ends

.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y a_27_47#
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.204706 pd=1.635294 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=6960,278
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.828235 as=0.143294 ps=1.144706 w=0.7 l=0.15
**devattr s=6960,278 d=7280,384
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=3510,184
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.611765 w=1 l=0.15
**devattr s=10400,504 d=4200,242
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=6760,364 d=4290,196
C0 A1 A2 0.098638f
C1 VPWR A2 0.10874f
C2 VGND A1 0.016299f
C3 VPWR VGND 0.038082f
C4 B1 A2 0.047196f
C5 A1 VPB 0.032652f
C6 VPWR VPB 0.056004f
C7 B1 VGND 0.016035f
C8 B1 VPB 0.074099f
C9 VGND A2 0.01829f
C10 Y VPWR 0.105149f
C11 a_27_47# A1 0.036956f
C12 VPB A2 0.030454f
C13 Y B1 0.081114f
C14 Y A2 0.123701f
C15 a_27_47# A2 0.038781f
C16 Y VGND 0.028878f
C17 a_27_47# VGND 0.142477f
C18 VPWR A1 0.049725f
C19 B1 VPWR 0.043328f
C20 Y a_27_47# 0.051702f
C21 VGND VNB 0.253652f
C22 Y VNB 0.054462f
C23 VPWR VNB 0.271009f
C24 B1 VNB 0.151859f
C25 A2 VNB 0.096175f
C26 A1 VNB 0.138363f
C27 VPB VNB 0.427572f
C28 a_27_47# VNB 0.031143f
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X a_27_413# a_207_413#
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111244 pd=0.929204 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=9116,348
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.264867 ps=2.212389 w=1 l=0.15
**devattr s=9116,348 d=10400,504
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2016,132
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13602 ps=1.457047 w=0.65 l=0.15
**devattr s=4052,198 d=6760,364
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.111244 ps=0.929204 w=0.42 l=0.15
**devattr s=2856,152 d=2436,142
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111244 pd=0.929204 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2856,152
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08789 pd=0.941476 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4052,198
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08789 ps=0.941476 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
C0 X VPWR 0.055194f
C1 B a_27_413# 0.092611f
C2 B VGND 0.01869f
C3 VPWR a_207_413# 0.111277f
C4 VPB X 0.012221f
C5 a_27_413# A_N 0.198147f
C6 VPB a_207_413# 0.047771f
C7 VGND A_N 0.047311f
C8 X a_207_413# 0.071579f
C9 a_27_413# VPWR 0.107953f
C10 VPWR VGND 0.056424f
C11 VPB a_27_413# 0.083441f
C12 B VPWR 0.086692f
C13 X VGND 0.065151f
C14 VPB B 0.111061f
C15 a_27_413# a_207_413# 0.185422f
C16 VPWR A_N 0.018219f
C17 X B 0.030307f
C18 VGND a_207_413# 0.114823f
C19 VPB A_N 0.080056f
C20 B a_207_413# 0.181991f
C21 a_27_413# VGND 0.086256f
C22 VPB VPWR 0.063352f
C23 VGND VNB 0.368472f
C24 X VNB 0.089221f
C25 VPWR VNB 0.291542f
C26 B VNB 0.132317f
C27 A_N VNB 0.201458f
C28 VPB VNB 0.604764f
C29 a_207_413# VNB 0.137402f
C30 a_27_413# VNB 0.196502f
.ends

.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X a_266_47# a_81_21#
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.117812 ps=1.0125 w=0.65 l=0.15
**devattr s=4745,203 d=2730,172
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169813 pd=1.1725 as=0.117812 ps=1.0125 w=0.65 l=0.15
**devattr s=4680,202 d=5460,214
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.23125 pd=1.4625 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=12500,325
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
**devattr s=2730,172 d=6760,364
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169813 pd=1.1725 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=8125,255
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.23125 ps=1.4625 w=1 l=0.15
**devattr s=12500,325 d=7200,272
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
**devattr s=7200,272 d=8400,284
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.117812 pd=1.0125 as=0.169813 ps=1.1725 w=0.65 l=0.15
**devattr s=5460,214 d=4745,203
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.117812 pd=1.0125 as=0.169813 ps=1.1725 w=0.65 l=0.15
**devattr s=8125,255 d=4680,202
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178333 pd=1.69 as=0.21 ps=1.42 w=1 l=0.15
**devattr s=8400,284 d=5500,255
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178333 pd=1.69 as=0.23125 ps=1.4625 w=1 l=0.15
**devattr s=6000,260 d=10400,504
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.23125 pd=1.4625 as=0.178333 ps=1.69 w=1 l=0.15
**devattr s=5500,255 d=6000,260
C0 a_81_21# A1 0.112746f
C1 VPB C1 0.038043f
C2 VGND A2 0.018378f
C3 X VPB 0.011438f
C4 a_368_297# A3 0.013389f
C5 B1 VPWR 0.016256f
C6 a_81_21# C1 0.118143f
C7 a_81_21# VPB 0.063191f
C8 X a_81_21# 0.08668f
C9 A2 VPWR 0.013141f
C10 VPB A3 0.03464f
C11 a_81_21# A3 0.08922f
C12 VGND VPWR 0.07715f
C13 B1 C1 0.058895f
C14 VPB B1 0.027915f
C15 A2 A1 0.076636f
C16 a_81_21# a_266_47# 0.043416f
C17 a_81_21# B1 0.092322f
C18 A2 VPB 0.031747f
C19 A3 a_266_47# 0.040304f
C20 VGND A1 0.045005f
C21 A3 B1 0.084907f
C22 a_81_21# A2 0.082341f
C23 a_81_21# a_266_297# 0.015752f
C24 X VGND 0.091215f
C25 B1 a_266_47# 0.03314f
C26 A2 A3 0.132989f
C27 a_81_21# VGND 0.136309f
C28 VPWR C1 0.02058f
C29 A2 a_266_47# 0.042515f
C30 VPB VPWR 0.074178f
C31 X VPWR 0.105139f
C32 VGND A3 0.01939f
C33 a_81_21# VPWR 0.487591f
C34 VGND a_266_47# 0.204958f
C35 VGND B1 0.016752f
C36 A3 VPWR 0.013837f
C37 VPB A1 0.031201f
C38 A2 a_266_297# 0.011011f
C39 a_368_297# a_81_21# 0.014848f
C40 VGND VNB 0.429376f
C41 VPWR VNB 0.361844f
C42 X VNB 0.093921f
C43 C1 VNB 0.144887f
C44 B1 VNB 0.092815f
C45 A3 VNB 0.09991f
C46 A2 VNB 0.092297f
C47 A1 VNB 0.09427f
C48 VPB VNB 0.781956f
C49 a_81_21# VNB 0.214691f
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X a_297_47# a_79_21#
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.943333 as=0.1525 ps=1.305 w=1 l=0.15
**devattr s=6100,261 d=10400,504
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.246667 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4030,192
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.246667 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.1235 ps=1.246667 w=0.65 l=0.15
**devattr s=4030,192 d=3510,184
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.943333 as=0.28 ps=2.56 w=1 l=0.15
**devattr s=11200,512 d=13100,331
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.305 ps=1.943333 w=1 l=0.15
**devattr s=13100,331 d=7800,278
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
**devattr s=7800,278 d=6100,261
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
C0 A2 a_79_21# 0.088854f
C1 A2 VPWR 0.083453f
C2 VPB X 0.011001f
C3 a_79_21# B1 0.13448f
C4 VGND a_297_47# 0.124631f
C5 VPWR B1 0.021269f
C6 A1 a_297_47# 0.049229f
C7 VGND a_79_21# 0.129186f
C8 A2 B1 0.06645f
C9 VGND VPWR 0.058833f
C10 A1 VPWR 0.044921f
C11 VGND A2 0.017086f
C12 VPB a_79_21# 0.048932f
C13 A2 A1 0.102437f
C14 VPB VPWR 0.062388f
C15 X a_79_21# 0.103737f
C16 X VPWR 0.095752f
C17 VGND B1 0.018231f
C18 VPB A2 0.033371f
C19 VPB B1 0.032789f
C20 VGND A1 0.015749f
C21 A2 a_382_297# 0.014523f
C22 a_79_21# a_297_47# 0.032587f
C23 A2 a_297_47# 0.048027f
C24 VPB A1 0.041226f
C25 a_79_21# VPWR 0.201029f
C26 VGND X 0.073624f
C27 VGND VNB 0.351611f
C28 VPWR VNB 0.304004f
C29 X VNB 0.09354f
C30 A1 VNB 0.152087f
C31 A2 VNB 0.098105f
C32 B1 VNB 0.101193f
C33 VPB VNB 0.604764f
C34 a_297_47# VNB 0.034813f
C35 a_79_21# VNB 0.158207f
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=10400,504
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=4200,242
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
C0 VPB Y 0.013918f
C1 A Y 0.047068f
C2 VGND Y 0.154448f
C3 VPB B 0.036697f
C4 VPWR Y 0.099513f
C5 A B 0.058413f
C6 VGND B 0.045088f
C7 a_109_297# Y 0.01129f
C8 VPWR B 0.014836f
C9 B Y 0.087653f
C10 VPB A 0.041461f
C11 VGND A 0.048556f
C12 VPB VPWR 0.044857f
C13 VPWR A 0.052823f
C14 VPWR VGND 0.031443f
C15 VGND VNB 0.263197f
C16 VPWR VNB 0.214143f
C17 Y VNB 0.060508f
C18 A VNB 0.14927f
C19 B VNB 0.143121f
C20 VPB VNB 0.338976f
.ends

.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X a_80_21# a_209_297#
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16875 pd=1.3375 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=6900,269
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.16875 ps=1.3375 w=1 l=0.15
**devattr s=6900,269 d=6400,264
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
**devattr s=4160,194 d=4290,196
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.144083 ps=1.31 w=0.65 l=0.15
**devattr s=4485,199 d=4160,194
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.144083 pd=1.31 as=0.17225 ps=1.83 w=0.65 l=0.15
**devattr s=6890,366 d=4485,199
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.144083 pd=1.31 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=8320,388
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=4290,196
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16875 pd=1.3375 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6400,264 d=6600,266
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6600,266 d=12800,528
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.16875 ps=1.3375 w=1 l=0.15
**devattr s=6600,266 d=6600,266
C0 A1 VGND 0.013522f
C1 A1 A2 0.104261f
C2 VPWR VPB 0.071542f
C3 A3 a_80_21# 0.116583f
C4 A2 a_209_297# 0.036649f
C5 X VPWR 0.117035f
C6 VGND VPWR 0.06622f
C7 a_80_21# VPB 0.050979f
C8 A2 VPWR 0.022678f
C9 B1 VPB 0.034195f
C10 A1 a_209_297# 0.037771f
C11 X a_80_21# 0.076532f
C12 A3 VPB 0.02968f
C13 a_80_21# VGND 0.216165f
C14 a_80_21# A2 0.035741f
C15 B1 VGND 0.017205f
C16 A1 VPWR 0.018013f
C17 a_80_21# a_303_47# 0.011458f
C18 A3 VGND 0.016898f
C19 a_209_297# VPWR 0.204727f
C20 A3 A2 0.108535f
C21 A1 a_80_21# 0.036671f
C22 A1 B1 0.101116f
C23 X VPB 0.010822f
C24 a_80_21# a_209_297# 0.062574f
C25 A2 VPB 0.028537f
C26 a_80_21# VPWR 0.09916f
C27 X VGND 0.057244f
C28 A3 a_209_297# 0.02681f
C29 B1 VPWR 0.01773f
C30 a_80_21# a_209_47# 0.010132f
C31 A2 VGND 0.014804f
C32 A1 VPB 0.028686f
C33 A3 VPWR 0.040256f
C34 a_80_21# B1 0.110759f
C35 VGND VNB 0.410332f
C36 VPWR VNB 0.331823f
C37 X VNB 0.08952f
C38 B1 VNB 0.11534f
C39 A1 VNB 0.089669f
C40 A2 VNB 0.089585f
C41 A3 VNB 0.089866f
C42 VPB VNB 0.69336f
C43 a_80_21# VNB 0.211154f
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X a_68_297#
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.087298 pd=0.938658 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.087298 ps=0.938658 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135104 ps=1.452685 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.086218 pd=0.789718 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.205282 ps=1.880282 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
C0 a_68_297# VPWR 0.088978f
C1 a_68_297# X 0.105343f
C2 a_68_297# A 0.157864f
C3 A B 0.07509f
C4 VPWR VPB 0.080528f
C5 X VPB 0.020902f
C6 a_68_297# B 0.098425f
C7 A VPB 0.030968f
C8 VGND VPWR 0.046447f
C9 VGND X 0.113947f
C10 a_68_297# VPB 0.061135f
C11 VPB B 0.046202f
C12 VGND A 0.034653f
C13 a_68_297# VGND 0.117961f
C14 VGND B 0.043653f
C15 VGND VPB 0.011204f
C16 X VPWR 0.128567f
C17 A X 0.013051f
C18 VGND VNB 0.320425f
C19 X VNB 0.100952f
C20 A VNB 0.110717f
C21 B VNB 0.182719f
C22 VPWR VNB 0.268565f
C23 VPB VNB 0.516168f
C24 a_68_297# VNB 0.153866f
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y a_113_297#
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=3835,189
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.181667 pd=1.696667 as=0.1475 ps=1.295 w=1 l=0.15
**devattr s=5900,259 d=10600,506
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
**devattr s=6890,366 d=3640,186
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.181667 ps=1.696667 w=1 l=0.15
**devattr s=5600,256 d=5900,259
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.181667 pd=1.696667 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
**devattr s=3835,189 d=6890,366
C0 VPWR Y 0.044654f
C1 B1 VPB 0.038865f
C2 A2 a_113_297# 0.047625f
C3 A2 VGND 0.049477f
C4 VPWR VPB 0.042396f
C5 B1 VPWR 0.01343f
C6 a_113_297# A1 0.050014f
C7 VGND A1 0.077964f
C8 A2 A1 0.091231f
C9 a_113_297# Y 0.09093f
C10 Y VGND 0.065351f
C11 a_113_297# VPB 0.010797f
C12 B1 VGND 0.043596f
C13 VPWR a_113_297# 0.1773f
C14 A2 VPB 0.037282f
C15 VPWR VGND 0.036961f
C16 Y A1 0.081255f
C17 VPWR A2 0.014703f
C18 A1 VPB 0.026387f
C19 B1 A1 0.051837f
C20 VPWR A1 0.015389f
C21 Y VPB 0.014642f
C22 B1 Y 0.112603f
C23 VGND VNB 0.285624f
C24 VPWR VNB 0.210674f
C25 Y VNB 0.054434f
C26 A2 VNB 0.143834f
C27 A1 VNB 0.098086f
C28 B1 VNB 0.161998f
C29 VPB VNB 0.427572f
C30 a_113_297# VNB 0.034004f
.ends

.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X a_240_47# a_51_297#
+ a_149_47#
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.114833 ps=1.22 w=0.65 l=0.15
**devattr s=3510,184 d=7280,372
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114833 pd=1.22 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.388333 pd=2.11 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=16500,365
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.122417 pd=1.243333 as=0.2015 ps=1.92 w=0.65 l=0.15
**devattr s=8060,384 d=3965,191
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.122417 ps=1.243333 w=0.65 l=0.15
**devattr s=3965,191 d=3510,184
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=6600,266
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=11200,512
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.122417 pd=1.243333 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=4200,242
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.388333 ps=2.11 w=1 l=0.15
**devattr s=13600,536 d=6600,266
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.388333 ps=2.11 w=1 l=0.15
**devattr s=16500,365 d=4200,242
C0 a_51_297# a_240_47# 0.03136f
C1 a_51_297# C1 0.10187f
C2 VPB A1 0.02547f
C3 VPWR A1 0.021536f
C4 VPWR VPB 0.087901f
C5 a_51_297# A1 0.12497f
C6 B2 a_240_47# 0.040822f
C7 a_51_297# VPB 0.063225f
C8 VPWR a_51_297# 0.414005f
C9 a_240_47# a_149_47# 0.068722f
C10 VPB B2 0.036569f
C11 VPWR B2 0.013541f
C12 A2 a_240_47# 0.056643f
C13 a_51_297# B2 0.077325f
C14 VGND X 0.143614f
C15 A2 A1 0.080079f
C16 B1 a_240_47# 0.011904f
C17 VPB A2 0.038559f
C18 B1 C1 0.051961f
C19 VPWR A2 0.015093f
C20 a_51_297# a_149_47# 0.024871f
C21 a_51_297# A2 0.088923f
C22 B1 VPB 0.025127f
C23 VGND a_240_47# 0.163798f
C24 VPWR B1 0.011497f
C25 VGND C1 0.014106f
C26 B2 A2 0.074588f
C27 a_51_297# B1 0.066861f
C28 VGND A1 0.027709f
C29 a_51_297# a_245_297# 0.012176f
C30 VPWR VGND 0.079939f
C31 B1 B2 0.079688f
C32 a_51_297# VGND 0.087412f
C33 B1 a_149_47# 0.017017f
C34 VPB X 0.026158f
C35 VPWR X 0.143364f
C36 VGND B2 0.010662f
C37 a_51_297# X 0.101431f
C38 VGND a_149_47# 0.122842f
C39 a_240_47# A1 0.023036f
C40 VGND A2 0.015861f
C41 VPB C1 0.05148f
C42 VPWR C1 0.020061f
C43 a_512_297# a_51_297# 0.011604f
C44 VGND VNB 0.493685f
C45 X VNB 0.106807f
C46 VPWR VNB 0.408842f
C47 A1 VNB 0.090821f
C48 A2 VNB 0.106876f
C49 B2 VNB 0.103396f
C50 B1 VNB 0.089709f
C51 C1 VNB 0.163785f
C52 VPB VNB 0.870552f
C53 a_240_47# VNB 0.013847f
C54 a_51_297# VNB 0.206675f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.102877 pd=0.95413 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.244946 ps=2.271739 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.087768 pd=0.816449 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.102877 ps=0.95413 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.135832 ps=1.263551 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
C0 VGND X 0.099328f
C1 VPWR VPB 0.072934f
C2 B a_59_75# 0.14331f
C3 VPWR VGND 0.046078f
C4 a_59_75# A 0.080877f
C5 B A 0.097088f
C6 a_59_75# X 0.10872f
C7 a_59_75# VPB 0.056305f
C8 VPWR a_59_75# 0.150282f
C9 VGND a_59_75# 0.115643f
C10 B VPB 0.06287f
C11 VPWR B 0.011747f
C12 VGND B 0.011461f
C13 A VPB 0.080573f
C14 VPWR A 0.036234f
C15 VGND A 0.014715f
C16 X VPB 0.012653f
C17 VPWR X 0.111215f
C18 VGND VNB 0.311398f
C19 X VNB 0.100184f
C20 B VNB 0.112872f
C21 A VNB 0.173792f
C22 VPWR VNB 0.273451f
C23 VPB VNB 0.516168f
C24 a_59_75# VNB 0.177062f
.ends

.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q a_891_413# a_193_47# a_381_47#
+ a_1062_300# a_475_413# a_634_183# a_27_47#
X0 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.199222 ps=1.797346 w=1 l=0.15
**devattr s=5700,257 d=5400,254
X1 a_1020_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0657 ps=0.725 w=0.36 l=0.15
**devattr s=2628,145 d=2640,149
X2 a_572_47# a_193_47# a_475_413# VNB sky130_fd_pr__nfet_01v8 ad=0.063415 pd=0.701538 as=0.0594 ps=0.69 w=0.36 l=0.15
**devattr s=2376,138 d=2748,152
X3 VPWR a_1062_300# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.083673 pd=0.754885 as=0.09135 ps=0.855 w=0.42 l=0.15
**devattr s=3654,171 d=4872,284
X4 a_634_183# a_475_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0.130634 ps=1.312053 w=0.64 l=0.15
**devattr s=5972,244 d=3956,199
X5 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.127502 pd=1.150302 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.083673 ps=0.754885 w=0.42 l=0.15
**devattr s=4368,272 d=2688,148
X7 a_475_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.060923 ps=0.687692 w=0.36 l=0.15
**devattr s=2640,149 d=2376,138
X8 VGND a_1062_300# a_1020_47# VNB sky130_fd_pr__nfet_01v8 ad=0.085728 pd=0.861035 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4788,282
X9 VPWR a_634_183# a_568_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.083673 pd=0.754885 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7155,252
X10 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.132675 ps=1.332554 w=0.65 l=0.15
**devattr s=3705,187 d=3510,184
X11 a_568_413# a_27_47# a_475_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2646,147 d=2772,150
X12 a_634_183# a_475_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0.149416 ps=1.34801 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X13 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3654,171
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.085728 ps=0.861035 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X15 a_891_413# a_27_47# a_634_183# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X16 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.132675 ps=1.332554 w=0.65 l=0.15
**devattr s=4225,195 d=3510,184
X17 VGND a_891_413# a_1062_300# VNB sky130_fd_pr__nfet_01v8 ad=0.132675 pd=1.332554 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4225,195
X18 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.199222 pd=1.797346 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5700,257
X19 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0.132675 pd=1.332554 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=7410,374
X20 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.199222 ps=1.797346 w=1 l=0.15
**devattr s=6500,265 d=5400,254
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.127502 ps=1.150302 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X22 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0.132675 pd=1.332554 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3705,187
X23 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.071077 pd=0.802308 as=0.085728 ps=0.861035 w=0.42 l=0.15
**devattr s=4368,272 d=2640,149
X24 VPWR a_891_413# a_1062_300# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.199222 pd=1.797346 as=0.28 ps=2.56 w=1 l=0.15
**devattr s=11200,512 d=6500,265
X25 a_891_413# a_193_47# a_634_183# VNB sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2628,145
X26 a_475_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
**devattr s=2688,148 d=2646,147
X27 VGND a_634_183# a_572_47# VNB sky130_fd_pr__nfet_01v8 ad=0.085728 pd=0.861035 as=0.073985 ps=0.818462 w=0.42 l=0.15
**devattr s=2748,152 d=5972,244
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.085728 pd=0.861035 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X29 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.199222 pd=1.797346 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=11200,512
C0 VPWR VGND 0.100633f
C1 a_27_47# a_1062_300# 0.048687f
C2 a_634_183# a_891_413# 0.035483f
C3 VGND a_193_47# 0.305428f
C4 D VPWR 0.027256f
C5 a_1062_300# a_891_413# 0.285494f
C6 VPB a_381_47# 0.013583f
C7 D a_193_47# 0.103962f
C8 VPB Q 0.013356f
C9 a_27_47# a_381_47# 0.03397f
C10 D VGND 0.026396f
C11 VPB a_27_47# 0.275432f
C12 a_634_183# a_475_413# 0.248641f
C13 VPWR CLK 0.019411f
C14 VPB a_891_413# 0.068757f
C15 a_27_47# a_891_413# 0.037767f
C16 VGND CLK 0.019463f
C17 a_634_183# VPWR 0.102093f
C18 a_381_47# a_475_413# 0.035644f
C19 VPB a_475_413# 0.075941f
C20 VPWR a_1062_300# 0.226048f
C21 a_634_183# a_193_47# 0.130991f
C22 a_193_47# a_1062_300# 0.030243f
C23 a_27_47# a_475_413# 0.178436f
C24 a_634_183# VGND 0.123913f
C25 VGND a_1062_300# 0.194826f
C26 a_381_47# VPWR 0.053383f
C27 VPB VPWR 0.198564f
C28 a_381_47# a_193_47# 0.16187f
C29 VPWR Q 0.335782f
C30 VPB a_193_47# 0.141384f
C31 a_27_47# VPWR 0.383097f
C32 a_381_47# VGND 0.044834f
C33 VPB VGND 0.014659f
C34 a_27_47# a_193_47# 0.723863f
C35 VPWR a_891_413# 0.113945f
C36 VGND Q 0.242058f
C37 D a_381_47# 0.076792f
C38 VPB D 0.09609f
C39 a_27_47# VGND 0.12468f
C40 a_193_47# a_891_413# 0.139283f
C41 a_27_47# D 0.096989f
C42 VGND a_891_413# 0.116731f
C43 VPWR a_475_413# 0.168224f
C44 VPB CLK 0.070057f
C45 a_193_47# a_475_413# 0.157543f
C46 VGND a_475_413# 0.09216f
C47 a_27_47# CLK 0.21376f
C48 VPB a_634_183# 0.073615f
C49 VPB a_1062_300# 0.24732f
C50 VPWR a_193_47# 0.106627f
C51 a_634_183# a_27_47# 0.166122f
C52 a_1062_300# Q 0.387919f
C53 Q VNB 0.060797f
C54 VGND VNB 0.988933f
C55 VPWR VNB 0.823111f
C56 D VNB 0.129726f
C57 CLK VNB 0.195983f
C58 VPB VNB 1.75651f
C59 a_381_47# VNB 0.016397f
C60 a_891_413# VNB 0.160892f
C61 a_1062_300# VNB 0.529662f
C62 a_475_413# VNB 0.137184f
C63 a_634_183# VNB 0.150209f
C64 a_193_47# VNB 0.271178f
C65 a_27_47# VNB 0.468295f
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X a_29_53#
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.208803 ps=1.887324 w=1 l=0.15
**devattr s=5930,268 d=11200,512
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.107931 ps=1.143456 w=0.65 l=0.15
**devattr s=4075,198 d=7280,372
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.087697 pd=0.792676 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.913333 as=0.06974 ps=0.738848 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.06974 pd=0.738848 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.06974 pd=0.738848 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
C0 VPB VPWR 0.064885f
C1 X VGND 0.035971f
C2 B a_29_53# 0.121149f
C3 VGND a_29_53# 0.216521f
C4 B VGND 0.0152f
C5 A a_29_53# 0.241867f
C6 VPB X 0.010881f
C7 C a_29_53# 0.085721f
C8 B A 0.07874f
C9 C B 0.080229f
C10 VPWR X 0.088535f
C11 VPB a_29_53# 0.049138f
C12 A VGND 0.018737f
C13 C VGND 0.016088f
C14 VPB B 0.096179f
C15 VPWR a_29_53# 0.08325f
C16 VPWR B 0.147145f
C17 C A 0.034282f
C18 VPWR VGND 0.045852f
C19 VPB A 0.037711f
C20 VPB C 0.039602f
C21 X a_29_53# 0.0991f
C22 VGND VNB 0.306355f
C23 X VNB 0.088191f
C24 A VNB 0.117495f
C25 C VNB 0.160014f
C26 B VNB 0.116674f
C27 VPWR VNB 0.252671f
C28 VPB VNB 0.516168f
C29 a_29_53# VNB 0.180006f
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X a_505_21# a_76_199#
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.084613 pd=0.797257 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.084613 ps=0.797257 w=0.42 l=0.15
**devattr s=2772,150 d=4704,280
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.084613 ps=0.797257 w=0.42 l=0.15
**devattr s=6334,279 d=3066,157
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.113356 pd=0.947749 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5796,222
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7728,268
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.113356 ps=0.947749 w=0.42 l=0.15
**devattr s=5796,222 d=4368,272
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
**devattr s=3990,179 d=2772,150
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
**devattr s=7728,268 d=1764,126
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=3990,179
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113356 ps=0.947749 w=0.42 l=0.15
**devattr s=4514,209 d=2772,150
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20146 pd=1.89823 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=6334,279
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.175432 pd=1.466754 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4514,209
C0 VPWR X 0.12783f
C1 A0 A1 0.266805f
C2 a_76_199# S 0.318161f
C3 VGND X 0.058643f
C4 VPB S 0.168493f
C5 VPWR VGND 0.080355f
C6 A1 S 0.087223f
C7 VPB a_505_21# 0.078063f
C8 a_76_199# X 0.077637f
C9 A0 S 0.034107f
C10 VPWR a_76_199# 0.054214f
C11 VPB X 0.012046f
C12 A1 a_505_21# 0.099273f
C13 VGND a_76_199# 0.160129f
C14 VPWR VPB 0.10994f
C15 VPB VGND 0.013448f
C16 A0 a_505_21# 0.038286f
C17 VPWR A1 0.011366f
C18 A1 VGND 0.075211f
C19 a_505_21# S 0.197515f
C20 VPB a_76_199# 0.048093f
C21 A0 VGND 0.043233f
C22 A1 a_76_199# 0.186672f
C23 VPWR S 0.392437f
C24 A1 VPB 0.072083f
C25 VGND S 0.032964f
C26 A0 a_76_199# 0.054443f
C27 VPWR a_505_21# 0.081832f
C28 A0 VPB 0.106597f
C29 a_505_21# VGND 0.123871f
C30 VGND VNB 0.498664f
C31 A1 VNB 0.140423f
C32 A0 VNB 0.13429f
C33 S VNB 0.268143f
C34 VPWR VNB 0.419248f
C35 X VNB 0.092356f
C36 VPB VNB 0.870552f
C37 a_505_21# VNB 0.246761f
C38 a_76_199# VNB 0.139466f
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.073937 pd=0.752655 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.073937 pd=0.752655 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103351 pd=0.894953 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.943333 as=0.073937 ps=0.752655 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.17604 ps=1.792035 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.159949 ps=1.385047 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
C0 VPB B 0.083634f
C1 X VGND 0.070777f
C2 X C 0.01492f
C3 VPWR VGND 0.047507f
C4 a_27_47# X 0.087038f
C5 A VPWR 0.018456f
C6 A VGND 0.015376f
C7 a_27_47# VPWR 0.145445f
C8 C VGND 0.07031f
C9 VPB X 0.012079f
C10 a_27_47# VGND 0.133608f
C11 B VPWR 0.128453f
C12 A a_27_47# 0.156874f
C13 B A 0.086925f
C14 a_27_47# C 0.1862f
C15 VPB VPWR 0.079461f
C16 B C 0.074622f
C17 VPB A 0.042605f
C18 B a_27_47# 0.062464f
C19 VPB C 0.034705f
C20 VPB a_27_47# 0.050077f
C21 X VPWR 0.076623f
C22 VGND VNB 0.300125f
C23 X VNB 0.092275f
C24 C VNB 0.120257f
C25 A VNB 0.174122f
C26 VPWR VNB 0.274246f
C27 B VNB 0.101788f
C28 VPB VNB 0.516168f
C29 a_27_47# VNB 0.177187f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.139399 ps=0.987313 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.331903 ps=2.350746 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.139399 ps=0.987313 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.139399 pd=0.987313 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.154085 pd=1.044112 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.139399 pd=0.987313 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.238465 ps=1.615888 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
C0 VPB B 0.064328f
C1 VPWR D 0.020729f
C2 VGND A 0.015122f
C3 VPWR B 0.023081f
C4 VPB a_27_47# 0.082046f
C5 a_27_47# D 0.106582f
C6 VPWR a_27_47# 0.326283f
C7 VPB C 0.060876f
C8 a_27_47# B 0.129725f
C9 VGND X 0.09025f
C10 C D 0.180159f
C11 A VPB 0.090662f
C12 VPWR C 0.021032f
C13 C B 0.160614f
C14 VPWR A 0.043995f
C15 A B 0.083909f
C16 a_27_47# C 0.051593f
C17 VGND D 0.089796f
C18 VPWR VGND 0.066176f
C19 A a_27_47# 0.15343f
C20 VGND B 0.045272f
C21 VPB X 0.011072f
C22 VPWR X 0.094506f
C23 VGND a_27_47# 0.13176f
C24 VPB D 0.078225f
C25 VGND C 0.040816f
C26 a_27_47# X 0.075371f
C27 VPWR VPB 0.076952f
C28 VGND VNB 0.39291f
C29 X VNB 0.093317f
C30 VPWR VNB 0.334542f
C31 D VNB 0.130267f
C32 C VNB 0.109828f
C33 B VNB 0.112123f
C34 A VNB 0.220977f
C35 VPB VNB 0.69336f
C36 a_27_47# VNB 0.174893f
.ends

.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X a_215_47# a_79_21#
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.256667 as=0.151667 ps=1.333333 w=0.65 l=0.15
**devattr s=6760,364 d=4225,195
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.151667 ps=1.333333 w=0.65 l=0.15
**devattr s=5720,218 d=4550,200
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.246667 pd=1.826667 as=0.2175 ps=1.935 w=1 l=0.15
**devattr s=7000,270 d=12000,520
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.935 as=0.246667 ps=1.826667 w=1 l=0.15
**devattr s=8800,288 d=7000,270
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.246667 pd=1.826667 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6500,265 d=8800,288
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.2175 ps=1.935 w=1 l=0.15
**devattr s=10400,504 d=6500,265
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
**devattr s=4550,200 d=7800,380
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.935 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.256667 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.151667 pd=1.333333 as=0.12675 ps=1.256667 w=0.65 l=0.15
**devattr s=4225,195 d=5720,218
C0 VGND a_215_47# 0.226322f
C1 VPB A1 0.032154f
C2 VPB A2 0.033967f
C3 X VPWR 0.128521f
C4 a_79_21# a_215_47# 0.045837f
C5 VGND a_79_21# 0.125897f
C6 VGND VPWR 0.073222f
C7 VGND B1 0.018554f
C8 a_79_21# VPWR 0.361146f
C9 B1 a_79_21# 0.064904f
C10 VGND C1 0.013287f
C11 B1 VPWR 0.018452f
C12 a_79_21# C1 0.096495f
C13 a_297_297# a_79_21# 0.017351f
C14 A1 a_215_47# 0.049321f
C15 C1 VPWR 0.020287f
C16 A2 a_215_47# 0.046109f
C17 VGND A1 0.017007f
C18 A2 VGND 0.015871f
C19 VPB X 0.01253f
C20 B1 C1 0.049531f
C21 a_297_297# VPWR 0.010695f
C22 A1 a_79_21# 0.084353f
C23 A2 a_79_21# 0.047445f
C24 A1 VPWR 0.018399f
C25 VPB VGND 0.010817f
C26 A2 VPWR 0.014254f
C27 A2 B1 0.061079f
C28 VPB a_79_21# 0.075544f
C29 VPB VPWR 0.094379f
C30 VPB B1 0.029836f
C31 VPB C1 0.055253f
C32 A2 A1 0.069292f
C33 VGND X 0.099278f
C34 X a_79_21# 0.049137f
C35 VGND VNB 0.449857f
C36 VPWR VNB 0.376877f
C37 X VNB 0.095064f
C38 C1 VNB 0.167477f
C39 B1 VNB 0.095044f
C40 A2 VNB 0.100735f
C41 A1 VNB 0.098893f
C42 VPB VNB 0.781956f
C43 a_215_47# VNB 0.01011f
C44 a_79_21# VNB 0.225128f
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X a_110_47#
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2310,139
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=4452,274
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5500,255
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=4452,274 d=2352,140
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2310,139 d=2352,140
C0 A VPWR 0.111641f
C1 VGND VPWR 0.187357f
C2 X VPWR 1.36494f
C3 A VPB 0.133397f
C4 VGND VPB 0.011388f
C5 X VPB 0.03148f
C6 a_110_47# A 0.306578f
C7 a_110_47# VGND 0.512392f
C8 VPB VPWR 0.183858f
C9 a_110_47# X 1.62234f
C10 a_110_47# VPWR 0.669976f
C11 a_110_47# VPB 0.527557f
C12 VGND A 0.115353f
C13 X VGND 0.976879f
C14 VGND VNB 1.01442f
C15 X VNB 0.110579f
C16 VPWR VNB 0.834786f
C17 A VNB 0.494734f
C18 VPB VNB 1.84511f
C19 a_110_47# VNB 1.73295f
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X a_81_21# a_299_297#
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.228583 ps=1.57 w=0.65 l=0.15
**devattr s=10270,288 d=3575,185
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.693333 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5500,255
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.693333 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.693333 as=0.18 ps=1.693333 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.228583 pd=1.57 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=10270,288
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.228583 pd=1.57 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=6890,366
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.693333 as=0.18 ps=1.693333 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
**devattr s=3575,185 d=3640,186
C0 B1 VGND 0.018138f
C1 X VGND 0.05115f
C2 A1 VPB 0.026428f
C3 A1 a_299_297# 0.058511f
C4 B1 VPB 0.038719f
C5 X VPB 0.010847f
C6 A1 VPWR 0.020947f
C7 VPWR VGND 0.057888f
C8 a_299_297# VPB 0.011077f
C9 A2 A1 0.092059f
C10 B1 VPWR 0.019602f
C11 a_81_21# A1 0.056842f
C12 VPWR X 0.084724f
C13 A2 VGND 0.049499f
C14 a_81_21# VGND 0.173386f
C15 a_81_21# B1 0.147666f
C16 VPWR VPB 0.068018f
C17 a_81_21# X 0.112205f
C18 a_299_297# VPWR 0.201825f
C19 A2 VPB 0.03733f
C20 a_81_21# VPB 0.05926f
C21 A2 a_299_297# 0.046825f
C22 a_81_21# a_299_297# 0.08213f
C23 A2 VPWR 0.020087f
C24 a_81_21# VPWR 0.145912f
C25 A1 VGND 0.078569f
C26 B1 A1 0.081725f
C27 VGND VNB 0.364132f
C28 VPWR VNB 0.285747f
C29 X VNB 0.094473f
C30 A2 VNB 0.144001f
C31 A1 VNB 0.099647f
C32 B1 VNB 0.108793f
C33 VPB VNB 0.604764f
C34 a_299_297# VNB 0.034794f
C35 a_81_21# VNB 0.147141f
.ends

.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X a_448_47# a_79_199#
+ a_222_93#
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066633 ps=0.67519 w=0.42 l=0.15
**devattr s=4010,197 d=4368,272
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.278216 pd=2.336257 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=11200,512
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.103122 pd=1.044937 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4010,197
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.116851 ps=0.981228 w=0.42 l=0.15
**devattr s=7430,283 d=4704,280
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103122 pd=1.044937 as=0.128917 ps=1.263333 w=0.65 l=0.15
**devattr s=4290,196 d=3510,184
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.128917 pd=1.263333 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4290,196
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.278216 ps=2.336257 w=1 l=0.15
**devattr s=12000,520 d=6600,266
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=4200,242
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.128917 pd=1.263333 as=0.103122 ps=1.044937 w=0.65 l=0.15
**devattr s=3510,184 d=6890,366
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.278216 pd=2.336257 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=7430,283
C0 A2 a_79_199# 0.060906f
C1 B1_N VPB 0.041907f
C2 VPWR VGND 0.074192f
C3 A1 VPWR 0.050783f
C4 a_79_199# VPB 0.067563f
C5 VGND B1_N 0.016051f
C6 X VPB 0.013182f
C7 VPWR a_222_93# 0.022446f
C8 A2 VPB 0.02588f
C9 a_79_199# VGND 0.083599f
C10 X VGND 0.060887f
C11 a_222_93# B1_N 0.106015f
C12 a_79_199# a_448_47# 0.046138f
C13 A2 VGND 0.015713f
C14 A2 A1 0.079314f
C15 a_79_199# a_222_93# 0.221119f
C16 VPWR a_544_297# 0.013205f
C17 A2 a_448_47# 0.058101f
C18 VGND VPB 0.011612f
C19 a_79_199# VPWR 0.263251f
C20 X VPWR 0.072913f
C21 A1 VPB 0.038356f
C22 A2 a_222_93# 0.056213f
C23 a_79_199# B1_N 0.083315f
C24 A2 VPWR 0.022715f
C25 a_222_93# VPB 0.063897f
C26 A1 VGND 0.017036f
C27 VGND a_448_47# 0.167957f
C28 X a_79_199# 0.109983f
C29 A1 a_448_47# 0.057384f
C30 VPWR VPB 0.109668f
C31 VGND a_222_93# 0.073067f
C32 VGND VNB 0.468282f
C33 B1_N VNB 0.105165f
C34 VPWR VNB 0.400387f
C35 X VNB 0.086477f
C36 A1 VNB 0.13607f
C37 A2 VNB 0.09044f
C38 VPB VNB 0.781956f
C39 a_448_47# VNB 0.032359f
C40 a_222_93# VNB 0.158855f
C41 a_79_199# VNB 0.148299f
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
C0 A VPWR 0.04444f
C1 VPB A 0.037877f
C2 Y VPWR 0.211407f
C3 A B 0.050963f
C4 Y B 0.048071f
C5 VPB VPWR 0.050862f
C6 B VPWR 0.047843f
C7 VPB B 0.039072f
C8 VGND Y 0.138901f
C9 VGND VPWR 0.032185f
C10 VGND B 0.054404f
C11 Y A 0.085479f
C12 VGND VNB 0.23167f
C13 Y VNB 0.055661f
C14 VPWR VNB 0.245114f
C15 A VNB 0.143376f
C16 B VNB 0.145827f
C17 VPB VNB 0.338976f
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X a_93_21# a_250_297#
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
**devattr s=5850,220 d=5720,218
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.193 ps=1.586 w=1 l=0.15
**devattr s=7400,274 d=5600,256
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
**devattr s=5720,218 d=2730,172
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.23375 pd=1.4675 as=0.33 ps=2.66 w=1 l=0.15
**devattr s=13200,532 d=9700,297
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.386667 as=0.06825 ps=0.86 w=0.65 l=0.15
**devattr s=2730,172 d=6890,366
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.169 ps=1.386667 w=0.65 l=0.15
**devattr s=6695,233 d=3900,190
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.586 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.386667 as=0.2145 ps=1.96 w=0.65 l=0.15
**devattr s=8580,392 d=6695,233
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.586 as=0.23375 ps=1.4675 w=1 l=0.15
**devattr s=9700,297 d=6600,266
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.23375 pd=1.4675 as=0.193 ps=1.586 w=1 l=0.15
**devattr s=6600,266 d=9000,290
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.586 as=0.23375 ps=1.4675 w=1 l=0.15
**devattr s=9000,290 d=7400,274
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
**devattr s=3900,190 d=5850,220
C0 a_93_21# a_250_297# 0.188241f
C1 B2 VPB 0.035517f
C2 a_93_21# A1 0.064134f
C3 X VPWR 0.084928f
C4 VGND VPWR 0.075955f
C5 A2 VPWR 0.013294f
C6 VGND B1 0.034397f
C7 A3 VPWR 0.015799f
C8 A1 VPB 0.029574f
C9 VGND B2 0.046938f
C10 a_93_21# VPB 0.048485f
C11 B1 VPWR 0.010035f
C12 a_250_297# A2 0.012898f
C13 A1 A2 0.09713f
C14 VGND A1 0.01333f
C15 B2 VPWR 0.010807f
C16 a_93_21# X 0.084123f
C17 B1 B2 0.082331f
C18 a_93_21# A2 0.074739f
C19 VGND a_93_21# 0.25085f
C20 a_250_297# VPWR 0.313499f
C21 a_93_21# A3 0.124344f
C22 A1 VPWR 0.015992f
C23 X VPB 0.010825f
C24 a_250_297# B1 0.012541f
C25 A1 B1 0.096524f
C26 A2 VPB 0.028677f
C27 a_93_21# a_256_47# 0.011416f
C28 a_93_21# VPWR 0.090657f
C29 a_250_297# B2 0.034435f
C30 A3 VPB 0.029118f
C31 a_93_21# B1 0.077421f
C32 VGND X 0.059994f
C33 VGND A2 0.011437f
C34 a_93_21# B2 0.014717f
C35 VPB VPWR 0.075576f
C36 A1 a_250_297# 0.012929f
C37 a_93_21# a_346_47# 0.011948f
C38 B1 VPB 0.027632f
C39 A3 A2 0.078809f
C40 VGND VNB 0.465075f
C41 VPWR VNB 0.364756f
C42 X VNB 0.093662f
C43 B2 VNB 0.140129f
C44 B1 VNB 0.100974f
C45 A1 VNB 0.095135f
C46 A2 VNB 0.092101f
C47 A3 VNB 0.092873f
C48 VPB VNB 0.781956f
C49 a_250_297# VNB 0.02777f
C50 a_93_21# VNB 0.150721f
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X a_80_21# a_217_297#
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.181667 pd=1.696667 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=10600,506
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
**devattr s=6200,262 d=10600,506
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.181667 pd=1.696667 as=0.181667 ps=1.696667 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.180375 pd=1.205 as=0.118083 ps=1.23 w=0.65 l=0.15
**devattr s=3640,186 d=4030,192
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.180375 pd=1.205 as=0.17225 ps=1.83 w=0.65 l=0.15
**devattr s=6890,366 d=10400,290
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.180375 ps=1.205 w=0.65 l=0.15
**devattr s=10400,290 d=3640,186
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.181667 pd=1.696667 as=0.181667 ps=1.696667 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.118083 pd=1.23 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=3640,186
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.181667 ps=1.696667 w=1 l=0.15
**devattr s=5600,256 d=6200,262
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118083 pd=1.23 as=0.180375 ps=1.205 w=0.65 l=0.15
**devattr s=4030,192 d=6890,366
C0 a_80_21# X 0.11763f
C1 A1 VGND 0.014726f
C2 B1 C1 0.084607f
C3 X VGND 0.065404f
C4 A2 VPB 0.038351f
C5 a_80_21# VPB 0.066072f
C6 a_80_21# a_472_297# 0.016359f
C7 A1 VPB 0.026604f
C8 X VPB 0.011762f
C9 a_80_21# VPWR 0.119311f
C10 A2 VPWR 0.016058f
C11 VPWR VGND 0.066493f
C12 C1 a_80_21# 0.079043f
C13 A1 VPWR 0.014884f
C14 a_217_297# a_80_21# 0.126609f
C15 A2 a_217_297# 0.013474f
C16 VPWR X 0.088406f
C17 C1 VGND 0.01758f
C18 a_217_297# A1 0.012424f
C19 VPWR VPB 0.075404f
C20 B1 a_80_21# 0.096355f
C21 B1 VGND 0.017479f
C22 C1 VPB 0.037912f
C23 B1 A1 0.083391f
C24 B1 VPB 0.026706f
C25 C1 VPWR 0.013731f
C26 a_217_297# VPWR 0.197242f
C27 A2 a_80_21# 0.127893f
C28 A2 VGND 0.019089f
C29 a_80_21# VGND 0.292585f
C30 B1 VPWR 0.01289f
C31 A2 A1 0.088064f
C32 A1 a_80_21# 0.111494f
C33 VGND VNB 0.38475f
C34 VPWR VNB 0.325154f
C35 X VNB 0.08992f
C36 C1 VNB 0.144368f
C37 B1 VNB 0.089926f
C38 A1 VNB 0.090508f
C39 A2 VNB 0.107869f
C40 VPB VNB 0.69336f
C41 a_80_21# VNB 0.209712f
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
C0 X VPWR 0.089678f
C1 VPB VPWR 0.035491f
C2 A VGND 0.018425f
C3 X VPB 0.012762f
C4 a_27_47# VGND 0.104759f
C5 A VPWR 0.021545f
C6 A VPB 0.052393f
C7 a_27_47# VPWR 0.135101f
C8 X a_27_47# 0.107446f
C9 a_27_47# VPB 0.059175f
C10 VGND VPWR 0.028968f
C11 X VGND 0.054627f
C12 a_27_47# A 0.181449f
C13 VGND VNB 0.207322f
C14 X VNB 0.094114f
C15 VPWR VNB 0.175402f
C16 A VNB 0.164055f
C17 VPB VNB 0.338976f
C18 a_27_47# VNB 0.207781f
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X a_489_413# a_226_47#
+ a_76_199#
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=4452,274
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.913333 as=0.083052 ps=0.789823 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.083052 ps=0.789823 w=0.42 l=0.15
**devattr s=6670,287 d=1764,126
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.083052 pd=0.789823 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.913333 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112949 ps=1.025665 w=0.42 l=0.15
**devattr s=5544,216 d=2268,138
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.112949 pd=1.025665 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.112949 pd=1.025665 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=5544,216
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112949 ps=1.025665 w=0.42 l=0.15
**devattr s=4804,217 d=2268,138
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.197743 pd=1.880531 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=6670,287
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.174803 pd=1.587339 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4804,217
C0 B1 a_489_413# 0.038152f
C1 a_76_199# a_226_47# 0.188181f
C2 A1_N VPB 0.033866f
C3 a_76_199# X 0.09953f
C4 A2_N VGND 0.017355f
C5 B1 VGND 0.047123f
C6 B2 a_489_413# 0.054108f
C7 B1 VPWR 0.018786f
C8 B2 VGND 0.033524f
C9 a_226_47# VPB 0.110695f
C10 A2_N A1_N 0.10971f
C11 X VPB 0.011346f
C12 B2 VPWR 0.016076f
C13 VPWR a_489_413# 0.142679f
C14 a_76_199# VPB 0.081664f
C15 a_226_47# A2_N 0.140761f
C16 VPWR VGND 0.074322f
C17 A1_N VGND 0.026061f
C18 B2 a_226_47# 0.097519f
C19 a_76_199# A2_N 0.012489f
C20 a_226_47# VGND 0.14876f
C21 a_76_199# B2 0.062591f
C22 X VGND 0.062661f
C23 A2_N VPB 0.032736f
C24 a_226_47# VPWR 0.018708f
C25 X VPWR 0.058912f
C26 a_76_199# a_489_413# 0.04732f
C27 B1 VPB 0.080343f
C28 a_76_199# VGND 0.108093f
C29 a_226_47# A1_N 0.020864f
C30 B2 VPB 0.064546f
C31 a_76_199# VPWR 0.199741f
C32 a_489_413# VPB 0.014986f
C33 a_76_199# A1_N 0.119207f
C34 VPB VGND 0.012835f
C35 X a_226_47# 0.010758f
C36 VPWR VPB 0.095098f
C37 B2 B1 0.181843f
C38 VGND VNB 0.461507f
C39 A2_N VNB 0.103283f
C40 A1_N VNB 0.111357f
C41 VPWR VNB 0.368878f
C42 X VNB 0.097534f
C43 B1 VNB 0.206073f
C44 B2 VNB 0.106213f
C45 VPB VNB 0.781956f
C46 a_489_413# VNB 0.025434f
C47 a_226_47# VNB 0.162324f
C48 a_76_199# VNB 0.140862f
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q a_543_47# a_193_47#
+ a_448_47# a_1283_21# a_761_289# a_1108_47# a_27_47#
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.061754 pd=0.692308 as=0.0711 ps=0.755 w=0.36 l=0.15
**devattr s=2844,151 d=2676,150
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.150877 ps=1.184615 w=0.42 l=0.15
**devattr s=5604,220 d=1764,126
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.179362 pd=1.667265 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.071928 ps=0.7092 w=0.36 l=0.15
**devattr s=3996,197 d=2844,151
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
**devattr s=2562,145 d=4368,272
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.1 as=0.07245 ps=0.765 w=0.42 l=0.15
**devattr s=2898,153 d=4620,194
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.222816 pd=2.269578 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115896 pd=1.077309 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5384,230
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.222816 ps=2.269578 w=1 l=0.15
**devattr s=12048,532 d=5400,254
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142602 pd=1.45253 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.093583 ps=0.953223 w=0.42 l=0.15
**devattr s=4368,272 d=2604,146
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127872 pd=1.2608 as=0.176603 ps=1.641614 w=0.64 l=0.15
**devattr s=5384,230 d=3996,197
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.115896 ps=1.077309 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0861 ps=0.79 w=0.42 l=0.15
**devattr s=5166,237 d=2352,140
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.060923 ps=0.687692 w=0.36 l=0.15
**devattr s=2640,149 d=2376,138
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.115896 ps=1.077309 w=0.42 l=0.15
**devattr s=4998,203 d=2562,145
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
**devattr s=2604,146 d=2898,153
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.071077 pd=0.802308 as=0.115896 ps=1.077309 w=0.42 l=0.15
**devattr s=8820,378 d=2640,149
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.093583 pd=0.953223 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3276,162
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.093583 pd=0.953223 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4536,276
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2268,138
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.142602 ps=1.45253 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.093583 ps=0.953223 w=0.42 l=0.15
**devattr s=3276,162 d=2268,138
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.093583 pd=0.953223 as=0.1134 ps=1.1 w=0.42 l=0.15
**devattr s=4620,194 d=2814,151
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.179362 ps=1.667265 w=0.65 l=0.15
**devattr s=8348,404 d=3510,184
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.129323 pd=1.015385 as=0.0594 ps=0.69 w=0.36 l=0.15
**devattr s=2376,138 d=5604,220
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115896 pd=1.077309 as=0.072046 ps=0.807692 w=0.42 l=0.15
**devattr s=2676,150 d=4998,203
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.1 as=0.093583 ps=0.953223 w=0.42 l=0.15
**devattr s=2814,151 d=4368,272
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115896 pd=1.077309 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1722 pd=1.58 as=0.187166 ps=1.906446 w=0.84 l=0.15
**devattr s=8736,440 d=5166,237
C0 RESET_B a_543_47# 0.153272f
C1 VPWR a_543_47# 0.100285f
C2 a_543_47# VPB 0.095793f
C3 a_1283_21# a_1108_47# 0.233657f
C4 a_27_47# a_1108_47# 0.102355f
C5 a_27_47# a_761_289# 0.07009f
C6 a_1283_21# Q 0.096297f
C7 a_193_47# RESET_B 0.026903f
C8 CLK VPWR 0.017406f
C9 RESET_B VGND 0.288034f
C10 a_193_47# VPWR 0.395957f
C11 CLK VPB 0.069345f
C12 VPWR VGND 0.071912f
C13 a_193_47# VPB 0.170907f
C14 a_448_47# a_543_47# 0.049827f
C15 a_27_47# a_543_47# 0.115353f
C16 VGND VPB 0.012153f
C17 a_651_413# a_761_289# 0.097745f
C18 a_651_413# a_543_47# 0.057222f
C19 a_761_289# a_1108_47# 0.051162f
C20 a_193_47# a_1283_21# 0.042509f
C21 CLK a_27_47# 0.233602f
C22 a_1283_21# VGND 0.259426f
C23 a_448_47# a_193_47# 0.064178f
C24 a_193_47# a_27_47# 0.906454f
C25 a_193_47# D 0.217945f
C26 a_27_47# VGND 0.253972f
C27 a_448_47# VGND 0.0661f
C28 D VGND 0.051614f
C29 RESET_B VPWR 0.065186f
C30 RESET_B VPB 0.138482f
C31 VPWR VPB 0.233696f
C32 a_193_47# a_651_413# 0.034619f
C33 a_761_289# a_543_47# 0.209641f
C34 RESET_B a_1283_21# 0.278919f
C35 a_27_47# RESET_B 0.296336f
C36 a_1283_21# VPWR 0.229753f
C37 a_193_47# a_1108_47# 0.125324f
C38 VGND a_1108_47# 0.148135f
C39 a_448_47# VPWR 0.068142f
C40 a_27_47# VPWR 0.152296f
C41 a_1283_21# VPB 0.168111f
C42 D VPWR 0.081188f
C43 a_193_47# a_761_289# 0.186387f
C44 a_27_47# VPB 0.261876f
C45 a_448_47# VPB 0.014137f
C46 D VPB 0.137565f
C47 a_761_289# VGND 0.073384f
C48 VGND Q 0.109665f
C49 a_651_413# RESET_B 0.012196f
C50 a_651_413# VPWR 0.12856f
C51 a_639_47# a_543_47# 0.013793f
C52 a_193_47# a_543_47# 0.229804f
C53 a_651_413# VPB 0.013543f
C54 VGND a_543_47# 0.122935f
C55 a_27_47# a_1283_21# 0.043587f
C56 a_448_47# a_27_47# 0.093133f
C57 RESET_B a_1108_47# 0.236601f
C58 a_448_47# D 0.155634f
C59 a_27_47# D 0.132849f
C60 VPWR a_1108_47# 0.173792f
C61 a_761_289# RESET_B 0.166114f
C62 VPB a_1108_47# 0.114634f
C63 a_761_289# VPWR 0.10497f
C64 CLK VGND 0.017208f
C65 a_193_47# VGND 0.063057f
C66 a_761_289# VPB 0.099418f
C67 VPWR Q 0.169355f
C68 Q VNB 0.029557f
C69 VGND VNB 1.09584f
C70 VPWR VNB 0.902284f
C71 RESET_B VNB 0.262848f
C72 D VNB 0.159894f
C73 CLK VNB 0.195254f
C74 VPB VNB 1.9337f
C75 a_448_47# VNB 0.013901f
C76 a_1108_47# VNB 0.13732f
C77 a_1283_21# VNB 0.389264f
C78 a_543_47# VNB 0.157869f
C79 a_761_289# VNB 0.120848f
C80 a_193_47# VNB 0.273213f
C81 a_27_47# VNB 0.495752f
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
R0A a_21_232# VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.0225
R0B a_21_232# HI sky130_fd_pr__res_generic_po w=0.48 l=0.0225
R1A a_159_232# LO sky130_fd_pr__res_generic_po w=0.48 l=0.0225
R1B a_159_232# VGND sky130_fd_pr__res_generic_po w=0.48 l=0.0225
C0 VPWR HI 0.072643f
C1 VGND LO 0.060475f
C2 VPB VPWR 0.157853f
C3 VGND HI 0.206798f
C4 HI LO 0.068275f
C5 VGND VPWR 0.031746f
C6 VPB LO 0.133883f
C7 VPWR LO 0.240897f
C8 VGND VNB 0.405957f
C9 LO VNB 0.165803f
C10 HI VNB 0.249567f
C11 VPWR VNB 0.297091f
C12 VPB VNB 0.338976f
.ends

.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X a_27_53# a_219_297#
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.114071 ps=0.949948 w=0.42 l=0.15
**devattr s=6300,234 d=2268,138
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.114071 pd=0.949948 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=6300,234
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.092605 pd=0.922174 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5930,268
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.176538 ps=1.470157 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.220489 ps=2.195652 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.092605 ps=0.922174 w=0.42 l=0.15
**devattr s=4368,272 d=4704,280
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0.114071 pd=0.949948 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
C0 a_219_297# VPB 0.047751f
C1 a_27_53# A 0.116384f
C2 VGND A 0.01651f
C3 VGND a_27_53# 0.144861f
C4 VPWR X 0.087835f
C5 VPB A 0.160525f
C6 a_27_53# VPB 0.045699f
C7 a_27_53# B_N 0.107716f
C8 VGND B_N 0.0173f
C9 VPB B_N 0.046613f
C10 a_219_297# VPWR 0.071899f
C11 VPWR A 0.194142f
C12 a_27_53# VPWR 0.037749f
C13 VGND VPWR 0.057039f
C14 VPWR VPB 0.097059f
C15 VPWR B_N 0.037442f
C16 a_219_297# X 0.094746f
C17 VGND X 0.035406f
C18 VPB X 0.010908f
C19 a_219_297# A 0.128105f
C20 a_219_297# a_27_53# 0.101254f
C21 VGND a_219_297# 0.134764f
C22 VGND VNB 0.353111f
C23 X VNB 0.08883f
C24 B_N VNB 0.169579f
C25 A VNB 0.135517f
C26 VPWR VNB 0.324987f
C27 VPB VNB 0.604764f
C28 a_27_53# VNB 0.175308f
C29 a_219_297# VNB 0.137194f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_285_297# a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.138125 ps=1.4 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.4 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.4 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.138125 ps=1.4 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
C0 a_35_297# VPB 0.069928f
C1 B A 0.221335f
C2 VPWR A 0.034845f
C3 B VPB 0.069694f
C4 VPWR VPB 0.068915f
C5 a_285_297# VPB 0.013272f
C6 VGND a_35_297# 0.176658f
C7 X VPB 0.015415f
C8 VPB A 0.051013f
C9 VGND B 0.030447f
C10 VPWR VGND 0.064265f
C11 VGND X 0.172898f
C12 B a_35_297# 0.203002f
C13 VPWR a_35_297# 0.096038f
C14 a_285_297# a_35_297# 0.025037f
C15 X a_35_297# 0.166001f
C16 VGND A 0.032545f
C17 VPWR B 0.070314f
C18 a_285_297# B 0.055317f
C19 VPWR a_285_297# 0.246305f
C20 a_35_297# A 0.063337f
C21 X B 0.014878f
C22 VPWR X 0.053654f
C23 X a_285_297# 0.071248f
C24 VGND VNB 0.434883f
C25 X VNB 0.064909f
C26 VPWR VNB 0.332777f
C27 A VNB 0.166719f
C28 B VNB 0.213371f
C29 VPB VNB 0.69336f
C30 a_35_297# VNB 0.254573f
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.723333 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=6500,265
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.723333 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.95 as=0.1113 ps=1.37 w=0.42 l=0.15
**devattr s=4452,274 d=2730,149
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.723333 w=1 l=0.15
**devattr s=6500,265 d=5400,254
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0819 ps=0.95 w=0.42 l=0.15
**devattr s=2730,149 d=2268,138
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.95 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
C0 a_27_47# VPWR 0.167265f
C1 VPB A 0.033457f
C2 VPWR VGND 0.038085f
C3 a_27_47# X 0.164973f
C4 X VGND 0.11464f
C5 a_27_47# A 0.208577f
C6 X VPWR 0.139126f
C7 A VGND 0.045291f
C8 a_27_47# VPB 0.068639f
C9 A VPWR 0.021971f
C10 VPB VPWR 0.043784f
C11 A X 0.012264f
C12 a_27_47# VGND 0.104722f
C13 VGND VNB 0.262974f
C14 X VNB 0.07314f
C15 VPWR VNB 0.220607f
C16 A VNB 0.147598f
C17 VPB VNB 0.427572f
C18 a_27_47# VNB 0.320141f
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X a_75_212#
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
C0 a_75_212# X 0.106512f
C1 VPB A 0.052491f
C2 X VGND 0.054484f
C3 a_75_212# VPWR 0.134042f
C4 VPWR VGND 0.028869f
C5 a_75_212# A 0.177899f
C6 VPWR X 0.089604f
C7 A VGND 0.018424f
C8 a_75_212# VPB 0.057101f
C9 VPB X 0.012788f
C10 A VPWR 0.021742f
C11 a_75_212# VGND 0.104971f
C12 VPB VPWR 0.035518f
C13 VGND VNB 0.20733f
C14 VPWR VNB 0.175531f
C15 X VNB 0.094159f
C16 A VNB 0.164205f
C17 VPB VNB 0.338976f
C18 a_75_212# VNB 0.210264f
.ends

.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X a_27_47#
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.206073 pd=1.674128 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=7800,380
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0.133155 pd=1.081744 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7006,253
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.305571 ps=2.383152 w=1 l=0.15
**devattr s=11198,323 d=6600,266
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
**devattr s=2478,143 d=3192,160
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.066675 pd=0.7375 as=0.12834 ps=1.000924 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305571 pd=2.383152 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=12000,520
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.066675 pd=0.7375 as=0.12834 ps=1.000924 w=0.42 l=0.15
**devattr s=4368,272 d=2982,155
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12834 pd=1.000924 as=0.066675 ps=0.7375 w=0.42 l=0.15
**devattr s=2352,140 d=11198,323
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.206073 ps=1.674128 w=0.65 l=0.15
**devattr s=7006,253 d=4290,196
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12834 pd=1.000924 as=0.066675 ps=0.7375 w=0.42 l=0.15
**devattr s=2982,155 d=3108,158
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2478,143
C0 VGND VPB 0.010944f
C1 VPB C 0.060875f
C2 a_27_47# VPWR 0.346707f
C3 VPWR B 0.023068f
C4 VPWR X 0.157615f
C5 VPWR A 0.040856f
C6 D VPWR 0.021477f
C7 a_27_47# VPB 0.113647f
C8 B VPB 0.064559f
C9 VPB A 0.090011f
C10 D VPB 0.079232f
C11 VGND C 0.037432f
C12 VPWR VPB 0.092393f
C13 a_27_47# VGND 0.153267f
C14 VGND B 0.041669f
C15 a_27_47# C 0.051213f
C16 X VGND 0.131519f
C17 B C 0.156914f
C18 VGND A 0.013622f
C19 D VGND 0.08079f
C20 D C 0.174741f
C21 a_27_47# B 0.126307f
C22 a_27_47# X 0.111239f
C23 VPWR VGND 0.086668f
C24 VPWR C 0.020869f
C25 a_27_47# A 0.154498f
C26 B A 0.082601f
C27 D a_27_47# 0.106425f
C28 VGND VNB 0.467438f
C29 X VNB 0.036881f
C30 VPWR VNB 0.397956f
C31 D VNB 0.12821f
C32 C VNB 0.109758f
C33 B VNB 0.112394f
C34 A VNB 0.219485f
C35 VPB VNB 0.781956f
C36 a_27_47# VNB 0.265166f
.ends

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X a_75_199# a_201_297#
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.256667 as=0.1235 ps=1.03 w=0.65 l=0.15
**devattr s=5395,213 d=6760,364
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.1235 ps=1.03 w=0.65 l=0.15
**devattr s=4485,199 d=5005,207
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125125 ps=1.035 w=0.65 l=0.15
**devattr s=5005,207 d=6760,234
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.12675 ps=1.256667 w=0.65 l=0.15
**devattr s=4225,195 d=5395,213
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.256667 as=0.169 ps=1.17 w=0.65 l=0.15
**devattr s=6760,234 d=4225,195
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2075 ps=1.415 w=1 l=0.15
**devattr s=8300,283 d=10400,504
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2075 pd=1.415 as=0.16375 ps=1.3275 w=1 l=0.15
**devattr s=6500,265 d=8300,283
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22375 pd=1.4475 as=0.285 ps=2.57 w=1 l=0.15
**devattr s=11400,514 d=5700,257
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16375 pd=1.3275 as=0.22375 ps=1.4475 w=1 l=0.15
**devattr s=5700,257 d=6600,266
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22375 pd=1.4475 as=0.16375 ps=1.3275 w=1 l=0.15
**devattr s=6600,266 d=12200,322
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16375 pd=1.3275 as=0.22375 ps=1.4475 w=1 l=0.15
**devattr s=12200,322 d=6500,265
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4485,199
C0 a_201_297# X 0.013143f
C1 A2 VGND 0.011854f
C2 VPWR C1 0.014612f
C3 A1 a_75_199# 0.069622f
C4 a_208_47# a_75_199# 0.015896f
C5 B1 C1 0.065975f
C6 VPB A3 0.026815f
C7 X a_75_199# 0.095935f
C8 VGND a_75_199# 0.362275f
C9 A1 VGND 0.011328f
C10 VPB C1 0.039357f
C11 B1 VPWR 0.012527f
C12 X VGND 0.060935f
C13 a_315_47# a_75_199# 0.020232f
C14 VPB VPWR 0.074935f
C15 A2 A3 0.074726f
C16 B1 VPB 0.029202f
C17 VPWR a_544_297# 0.010504f
C18 A3 a_75_199# 0.163342f
C19 C1 a_75_199# 0.062832f
C20 A3 VGND 0.01613f
C21 A2 VPWR 0.017412f
C22 VPWR a_201_297# 0.211447f
C23 C1 VGND 0.018145f
C24 VPWR a_75_199# 0.109364f
C25 B1 a_75_199# 0.102254f
C26 A1 VPWR 0.015144f
C27 B1 A1 0.071566f
C28 A2 VPB 0.037631f
C29 VPWR X 0.067555f
C30 VPWR VGND 0.07349f
C31 B1 VGND 0.017055f
C32 VPB a_75_199# 0.048628f
C33 a_544_297# a_75_199# 0.017594f
C34 A1 VPB 0.030611f
C35 VPB X 0.010651f
C36 A2 a_201_297# 0.011242f
C37 A2 a_75_199# 0.062124f
C38 a_201_297# a_75_199# 0.159564f
C39 VPWR A3 0.018105f
C40 A2 A1 0.068871f
C41 A1 a_201_297# 0.011032f
C42 VGND VNB 0.436573f
C43 VPWR VNB 0.365173f
C44 X VNB 0.090646f
C45 C1 VNB 0.14827f
C46 B1 VNB 0.094718f
C47 A1 VNB 0.101248f
C48 A2 VNB 0.110292f
C49 A3 VNB 0.090791f
C50 VPB VNB 0.781956f
C51 a_75_199# VNB 0.20459f
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X a_489_47# a_206_369#
+ a_76_199#
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.128382 ps=1.053134 w=0.42 l=0.15
**devattr s=5830,267 d=5160,236
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2646,147 d=4368,272
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06831 pd=0.73445 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
**devattr s=2688,148 d=1764,126
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.913333 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.913333 as=0.06831 ps=0.73445 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128382 pd=1.053134 as=0.129 ps=1.18 w=0.42 l=0.15
**devattr s=5160,236 d=8370,269
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.128382 ps=1.053134 w=0.42 l=0.15
**devattr s=8370,269 d=2688,148
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.06831 ps=0.73445 w=0.42 l=0.15
**devattr s=3945,196 d=2646,147
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305672 pd=2.507463 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5830,267
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128382 pd=1.053134 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=4368,272
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.105719 pd=1.136649 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3945,196
C0 a_76_199# a_489_47# 0.049785f
C1 a_206_369# VPWR 0.020722f
C2 B1 VPWR 0.048982f
C3 a_76_199# VPB 0.059746f
C4 A2_N VPB 0.053423f
C5 a_206_369# A1_N 0.029727f
C6 VPB VPWR 0.108864f
C7 a_76_199# VGND 0.066825f
C8 VPB A1_N 0.062218f
C9 VGND A2_N 0.064685f
C10 B1 a_489_47# 0.05284f
C11 a_206_369# VPB 0.097704f
C12 B1 VPB 0.06625f
C13 VGND VPWR 0.072388f
C14 VGND A1_N 0.027491f
C15 a_206_369# VGND 0.057063f
C16 B1 VGND 0.016305f
C17 VGND a_489_47# 0.136725f
C18 a_76_199# X 0.095561f
C19 X VPWR 0.061845f
C20 X VPB 0.010949f
C21 VGND X 0.086091f
C22 a_76_199# B2 0.122643f
C23 B2 VPWR 0.088044f
C24 a_206_369# B2 0.088505f
C25 B1 B2 0.162675f
C26 a_489_47# B2 0.063279f
C27 B2 VPB 0.055976f
C28 a_76_199# A2_N 0.01425f
C29 a_76_199# VPWR 0.195754f
C30 VGND B2 0.016247f
C31 a_76_199# A1_N 0.090301f
C32 A2_N A1_N 0.09394f
C33 a_76_199# a_206_369# 0.266837f
C34 a_206_369# A2_N 0.150178f
C35 VPWR A1_N 0.010805f
C36 VGND VNB 0.452597f
C37 B1 VNB 0.181469f
C38 B2 VNB 0.105231f
C39 A2_N VNB 0.125702f
C40 A1_N VNB 0.121561f
C41 VPWR VNB 0.391659f
C42 X VNB 0.094468f
C43 VPB VNB 0.781956f
C44 a_489_47# VNB 0.037211f
C45 a_206_369# VNB 0.153769f
C46 a_76_199# VNB 0.136541f
.ends

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X a_27_297# a_109_297#
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.187633 pd=1.713333 as=0.1475 ps=1.295 w=1 l=0.15
**devattr s=6400,264 d=6200,262
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
**devattr s=2990,176 d=6760,364
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.246667 as=0.11375 ps=1 w=0.65 l=0.15
**devattr s=4550,200 d=4030,192
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.187633 ps=1.713333 w=1 l=0.15
**devattr s=6200,262 d=10400,504
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.256425 pd=2.52 as=0.1475 ps=1.295 w=1 l=0.15
**devattr s=5400,254 d=10114,504
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.187633 ps=1.713333 w=1 l=0.15
**devattr s=10116,504 d=6400,264
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4550,200
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1235 ps=1.246667 w=0.65 l=0.15
**devattr s=4030,192 d=6760,364
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.256425 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.1235 ps=1.246667 w=0.65 l=0.15
**devattr s=6760,364 d=2990,176
C0 A1 VGND 0.013674f
C1 A2 a_27_297# 0.161036f
C2 B2 VGND 0.053784f
C3 VPWR X 0.09141f
C4 VGND a_27_297# 0.256693f
C5 A1 VPB 0.038674f
C6 A2 VGND 0.016221f
C7 VPB B2 0.029852f
C8 VPB a_27_297# 0.059098f
C9 A2 VPB 0.028389f
C10 A1 B1 0.065706f
C11 B2 B1 0.073857f
C12 B1 a_27_297# 0.083756f
C13 B1 a_109_297# 0.01063f
C14 X a_27_297# 0.108071f
C15 B1 VGND 0.026654f
C16 A1 VPWR 0.016808f
C17 X VGND 0.054267f
C18 VPB B1 0.03168f
C19 VPWR B2 0.012568f
C20 VPWR a_27_297# 0.129594f
C21 VPWR a_109_297# 0.187005f
C22 VPWR A2 0.017794f
C23 VPB X 0.011018f
C24 VPWR VGND 0.064099f
C25 a_373_47# a_27_297# 0.013377f
C26 VPWR VPB 0.07143f
C27 A1 a_27_297# 0.083856f
C28 B2 a_27_297# 0.056703f
C29 A1 a_109_297# 0.010516f
C30 VPWR B1 0.013891f
C31 A1 A2 0.073773f
C32 a_27_297# a_109_297# 0.171361f
C33 VGND VNB 0.421193f
C34 X VNB 0.091659f
C35 VPWR VNB 0.328062f
C36 A2 VNB 0.092694f
C37 A1 VNB 0.111912f
C38 B1 VNB 0.111541f
C39 B2 VNB 0.126407f
C40 VPB VNB 0.69336f
C41 a_27_297# VNB 0.190287f
.ends

.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X a_103_199# a_253_47#
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.0975 ps=0.95 w=0.65 l=0.15
**devattr s=4290,196 d=8060,384
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.245 pd=1.823333 as=0.36 ps=2.72 w=1 l=0.15
**devattr s=14400,544 d=7800,278
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=6600,266
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=8500,285
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.245 ps=1.823333 w=1 l=0.15
**devattr s=7800,278 d=5400,254
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.245 pd=1.823333 as=0.2125 ps=1.425 w=1 l=0.15
**devattr s=8500,285 d=13800,538
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.234 ps=2.02 w=0.65 l=0.15
**devattr s=9360,404 d=5070,208
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.117 ps=1.01 w=0.65 l=0.15
**devattr s=5070,208 d=3510,184
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.117 ps=1.01 w=0.65 l=0.15
**devattr s=4290,196 d=4290,196
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0975 ps=0.95 w=0.65 l=0.15
**devattr s=3510,184 d=4290,196
C0 X VPB 0.01546f
C1 A2 VPB 0.028397f
C2 VGND A3 0.013887f
C3 A2 A1 0.080246f
C4 VGND B1 0.015441f
C5 VPB A3 0.031009f
C6 a_103_199# VPWR 0.377206f
C7 VPB B1 0.034421f
C8 VGND A1 0.04324f
C9 VPB A1 0.027104f
C10 X a_103_199# 0.076224f
C11 a_253_297# a_103_199# 0.014832f
C12 A2 a_103_199# 0.085597f
C13 a_103_199# A3 0.085357f
C14 a_103_199# B1 0.102311f
C15 a_337_297# a_103_199# 0.01015f
C16 VGND a_103_199# 0.101569f
C17 a_103_199# VPB 0.049224f
C18 a_103_199# A1 0.123481f
C19 a_253_47# A2 0.030298f
C20 a_253_47# A3 0.030041f
C21 a_253_47# B1 0.013003f
C22 VGND a_253_47# 0.199693f
C23 X VPWR 0.120185f
C24 VPWR A3 0.011038f
C25 VPWR B1 0.018978f
C26 VGND VPWR 0.06508f
C27 VPB VPWR 0.072655f
C28 VPWR A1 0.011487f
C29 A2 A3 0.136697f
C30 a_253_47# a_103_199# 0.060607f
C31 VGND X 0.109334f
C32 A3 B1 0.073596f
C33 VGND A2 0.013332f
C34 VGND VNB 0.39103f
C35 VPWR VNB 0.349144f
C36 X VNB 0.097222f
C37 B1 VNB 0.121351f
C38 A3 VNB 0.089564f
C39 A2 VNB 0.08849f
C40 A1 VNB 0.090241f
C41 VPB VNB 0.69336f
C42 a_253_47# VNB 0.011031f
C43 a_103_199# VNB 0.196442f
.ends

.subckt r2r_dac_control clk data[0] data[1] data[2] data[3] data[4] data[5] data[6]
+ data[7] ext_data load_divider n_rst r2r_out[0] r2r_out[1] r2r_out[2] r2r_out[3]
+ r2r_out[4] r2r_out[5] r2r_out[6] r2r_out[7] VPWR VGND
X_294_ _046_ divider\[5\] divider\[4\] _041_ VGND VGND VPWR VPWR _047_ _294_/a_78_199#
+ _294_/a_215_47# sky130_fd_sc_hd__o22a_1
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_346_ clknet_2_0__leaf_clk _022_ VGND VGND VPWR VPWR counter\[5\] _346_/a_891_413#
+ _346_/a_466_413# _346_/a_1059_315# _346_/a_193_47# _346_/a_634_159# _346_/a_381_47#
+ _346_/a_27_47# sky130_fd_sc_hd__dfxtp_1
X_277_ counter\[10\] VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__inv_2
X_200_ _094_ _101_ _102_ _103_ _078_ VGND VGND VPWR VPWR _104_ _200_/a_227_47# _200_/a_77_199#
+ sky130_fd_sc_hd__o32a_1
X_329_ clknet_2_2__leaf_clk _005_ VGND VGND VPWR VPWR divider\[4\] _329_/a_891_413#
+ _329_/a_466_413# _329_/a_1059_315# _329_/a_193_47# _329_/a_634_159# _329_/a_381_47#
+ _329_/a_27_47# sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_293_ counter\[13\] VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_74 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_276_ net8 _148_ _158_ VGND VGND VPWR VPWR _008_ _276_/a_215_297# _276_/a_27_413#
+ _276_/a_298_297# sky130_fd_sc_hd__a21bo_1
X_345_ clknet_2_1__leaf_clk _021_ VGND VGND VPWR VPWR counter\[4\] _345_/a_891_413#
+ _345_/a_466_413# _345_/a_1059_315# _345_/a_193_47# _345_/a_634_159# _345_/a_381_47#
+ _345_/a_27_47# sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_259_ rst VGND VGND VPWR VPWR _149_ _259_/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_328_ clknet_2_2__leaf_clk _004_ VGND VGND VPWR VPWR divider\[3\] _328_/a_891_413#
+ _328_/a_466_413# _328_/a_1059_315# _328_/a_193_47# _328_/a_634_159# _328_/a_381_47#
+ _328_/a_27_47# sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_292_ _034_ _036_ _040_ _042_ _044_ VGND VGND VPWR VPWR _045_ _292_/a_516_297# _292_/a_85_193#
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_275_ net10 rst divider\[7\] VGND VGND VPWR VPWR _158_ _275_/a_215_53# _275_/a_109_93#
+ sky130_fd_sc_hd__or3b_1
X_344_ clknet_2_0__leaf_clk _020_ VGND VGND VPWR VPWR counter\[3\] _344_/a_891_413#
+ _344_/a_466_413# _344_/a_1059_315# _344_/a_193_47# _344_/a_634_159# _344_/a_381_47#
+ _344_/a_27_47# sky130_fd_sc_hd__dfxtp_1
X_327_ clknet_2_3__leaf_clk _003_ VGND VGND VPWR VPWR divider\[2\] _327_/a_891_413#
+ _327_/a_466_413# _327_/a_1059_315# _327_/a_193_47# _327_/a_634_159# _327_/a_381_47#
+ _327_/a_27_47# sky130_fd_sc_hd__dfxtp_1
X_258_ net10 VGND VGND VPWR VPWR _148_ _258_/a_27_47# sky130_fd_sc_hd__buf_2
X_189_ counter\[1\] counter\[0\] VGND VGND VPWR VPWR _095_ _189_/a_47_47# _189_/a_285_47#
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold10 r2r_out[7] VGND VGND VPWR VPWR net22 hold10/a_49_47# hold10/a_285_47# hold10/a_391_47#
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_291_ _041_ divider\[4\] divider\[3\] _035_ _043_ VGND VGND VPWR VPWR _044_ _291_/a_193_297#
+ _291_/a_109_297# _291_/a_27_47# sky130_fd_sc_hd__a221o_1
XFILLER_0_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_274_ _148_ net7 _157_ VGND VGND VPWR VPWR _007_ _274_/a_215_297# _274_/a_27_413#
+ _274_/a_298_297# sky130_fd_sc_hd__a21bo_1
X_343_ clknet_2_1__leaf_clk _019_ VGND VGND VPWR VPWR counter\[2\] _343_/a_891_413#
+ _343_/a_466_413# _343_/a_1059_315# _343_/a_193_47# _343_/a_634_159# _343_/a_381_47#
+ _343_/a_27_47# sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_257_ net11 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
X_326_ clknet_2_3__leaf_clk _002_ VGND VGND VPWR VPWR divider\[1\] _326_/a_891_413#
+ _326_/a_466_413# _326_/a_1059_315# _326_/a_193_47# _326_/a_634_159# _326_/a_381_47#
+ _326_/a_27_47# sky130_fd_sc_hd__dfxtp_1
X_188_ _052_ VGND VGND VPWR VPWR _094_ _188_/a_27_47# sky130_fd_sc_hd__buf_2
XFILLER_0_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_309_ _060_ _055_ r2r_out[1] VGND VGND VPWR VPWR _061_ _309_/a_27_47# sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_290_ counter\[13\] divider\[5\] VGND VGND VPWR VPWR _043_ _290_/a_27_413# _290_/a_207_413#
+ sky130_fd_sc_hd__and2b_1
X_273_ net10 rst divider\[6\] VGND VGND VPWR VPWR _157_ _273_/a_215_53# _273_/a_109_93#
+ sky130_fd_sc_hd__or3b_1
X_342_ clknet_2_1__leaf_clk _018_ VGND VGND VPWR VPWR counter\[1\] _342_/a_891_413#
+ _342_/a_466_413# _342_/a_1059_315# _342_/a_193_47# _342_/a_634_159# _342_/a_381_47#
+ _342_/a_27_47# sky130_fd_sc_hd__dfxtp_1
X_325_ clknet_2_2__leaf_clk _001_ VGND VGND VPWR VPWR divider\[0\] _325_/a_891_413#
+ _325_/a_466_413# _325_/a_1059_315# _325_/a_193_47# _325_/a_634_159# _325_/a_381_47#
+ _325_/a_27_47# sky130_fd_sc_hd__dfxtp_1
X_256_ _146_ _066_ _143_ _147_ _057_ VGND VGND VPWR VPWR _032_ _256_/a_266_47# _256_/a_81_21#
+ sky130_fd_sc_hd__o311a_1
X_187_ net19 _060_ _093_ VGND VGND VPWR VPWR _017_ _187_/a_297_47# _187_/a_79_21#
+ sky130_fd_sc_hd__o21a_1
X_239_ _065_ _134_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__nor2_1
X_308_ _059_ VGND VGND VPWR VPWR _060_ _308_/a_27_47# sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_272_ _148_ net6 _156_ VGND VGND VPWR VPWR _006_ _272_/a_215_297# _272_/a_27_413#
+ _272_/a_298_297# sky130_fd_sc_hd__a21bo_1
X_341_ clknet_2_1__leaf_clk _017_ VGND VGND VPWR VPWR counter\[0\] _341_/a_891_413#
+ _341_/a_466_413# _341_/a_1059_315# _341_/a_193_47# _341_/a_634_159# _341_/a_381_47#
+ _341_/a_27_47# sky130_fd_sc_hd__dfxtp_1
X_255_ counter\[14\] _060_ _141_ counter\[15\] VGND VGND VPWR VPWR _147_ _255_/a_80_21#
+ _255_/a_209_297# sky130_fd_sc_hd__a31o_1
X_324_ r2r_out[3] _069_ VGND VGND VPWR VPWR _074_ _324_/a_68_297# sky130_fd_sc_hd__or2_1
X_186_ _078_ counter\[0\] _149_ VGND VGND VPWR VPWR _093_ _186_/a_113_297# sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_169_ r2r_out[4] _076_ _079_ _060_ _057_ VGND VGND VPWR VPWR _013_ _169_/a_240_47#
+ _169_/a_51_297# _169_/a_149_47# sky130_fd_sc_hd__o221a_1
X_238_ _094_ _131_ _133_ _035_ _078_ VGND VGND VPWR VPWR _134_ _238_/a_227_47# _238_/a_77_199#
+ sky130_fd_sc_hd__o32a_1
X_307_ _045_ _051_ VGND VGND VPWR VPWR _059_ _307_/a_59_75# sky130_fd_sc_hd__and2_1
XFILLER_0_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_340_ clknet_2_3__leaf_clk _016_ VGND VGND VPWR VPWR r2r_out[7] _340_/a_891_413#
+ _340_/a_193_47# _340_/a_381_47# _340_/a_1062_300# _340_/a_475_413# _340_/a_634_183#
+ _340_/a_27_47# sky130_fd_sc_hd__dfxtp_4
X_271_ net10 _155_ _149_ VGND VGND VPWR VPWR _156_ _271_/a_29_53# sky130_fd_sc_hd__or3_1
X_185_ _090_ _092_ _065_ VGND VGND VPWR VPWR _016_ _185_/a_113_297# sky130_fd_sc_hd__a21oi_1
X_254_ net20 VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__inv_2
X_323_ _054_ _072_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_168_ net5 _077_ _078_ VGND VGND VPWR VPWR _079_ _168_/a_505_21# _168_/a_76_199#
+ sky130_fd_sc_hd__mux2_1
X_237_ counter\[7\] _112_ _132_ VGND VGND VPWR VPWR _133_ _237_/a_27_47# sky130_fd_sc_hd__and3_1
X_306_ _053_ _056_ _058_ VGND VGND VPWR VPWR _009_ _306_/a_113_297# sky130_fd_sc_hd__a21oi_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_270_ divider\[5\] VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__inv_2
X_322_ r2r_out[3] r2r_out[2] r2r_out[1] r2r_out[0] VGND VGND VPWR VPWR _072_ _322_/a_27_47#
+ sky130_fd_sc_hd__and4_1
X_184_ _060_ _091_ net22 VGND VGND VPWR VPWR _092_ _184_/a_27_47# sky130_fd_sc_hd__o21ai_1
X_253_ _066_ _143_ _145_ _057_ VGND VGND VPWR VPWR _031_ _253_/a_215_47# _253_/a_79_21#
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_167_ _048_ VGND VGND VPWR VPWR _078_ _167_/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_305_ _053_ _056_ _057_ VGND VGND VPWR VPWR _058_ _305_/a_27_47# sky130_fd_sc_hd__o21ai_1
X_236_ counter\[11\] counter\[10\] counter\[9\] counter\[8\] VGND VGND VPWR VPWR _132_
+ _236_/a_27_47# sky130_fd_sc_hd__and4_1
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_219_ _094_ _115_ _117_ _118_ _078_ VGND VGND VPWR VPWR _119_ _219_/a_227_47# _219_/a_77_199#
+ sky130_fd_sc_hd__o32a_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk clkbuf_0_clk/a_110_47# sky130_fd_sc_hd__clkbuf_16
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_183_ _078_ _084_ VGND VGND VPWR VPWR _091_ _183_/a_59_75# sky130_fd_sc_hd__and2_1
X_252_ _060_ _144_ counter\[14\] VGND VGND VPWR VPWR _145_ _252_/a_81_21# _252_/a_299_297#
+ sky130_fd_sc_hd__a21o_1
X_321_ net21 _053_ _071_ VGND VGND VPWR VPWR _011_ _321_/a_448_47# _321_/a_79_199#
+ _321_/a_222_93# sky130_fd_sc_hd__o21ba_1
X_304_ rst VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_235_ counter\[10\] _126_ counter\[11\] VGND VGND VPWR VPWR _131_ _235_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
X_166_ r2r_out[4] _072_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_218_ net18 VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk clkbuf_2_0__f_clk/a_110_47#
+ sky130_fd_sc_hd__clkbuf_16
X_182_ _053_ _089_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_251_ counter\[13\] counter\[12\] _136_ VGND VGND VPWR VPWR _144_ _251_/a_27_47#
+ sky130_fd_sc_hd__and3_1
X_320_ _053_ _067_ _070_ _149_ VGND VGND VPWR VPWR _071_ _320_/a_80_21# _320_/a_209_297#
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_165_ _060_ _073_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_303_ _054_ net1 _055_ VGND VGND VPWR VPWR _056_ _303_/a_113_297# sky130_fd_sc_hd__a21oi_1
X_234_ _128_ _130_ _149_ VGND VGND VPWR VPWR _027_ _234_/a_113_297# sky130_fd_sc_hd__a21oi_1
X_217_ counter\[7\] counter\[4\] _101_ _116_ VGND VGND VPWR VPWR _117_ _217_/a_27_47#
+ sky130_fd_sc_hd__and4_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_49 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_181_ r2r_out[6] _081_ _088_ net8 _054_ VGND VGND VPWR VPWR _089_ _181_/a_93_21#
+ _181_/a_250_297# sky130_fd_sc_hd__a32o_1
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_250_ counter\[14\] _141_ _053_ VGND VGND VPWR VPWR _143_ _250_/a_113_297# sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_164_ r2r_out[3] _053_ _075_ _057_ VGND VGND VPWR VPWR _012_ _164_/a_215_47# _164_/a_79_21#
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_302_ _054_ r2r_out[0] VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__nor2_1
X_233_ counter\[10\] _126_ _129_ _094_ VGND VGND VPWR VPWR _130_ _233_/a_80_21# _233_/a_217_297#
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_216_ counter\[6\] counter\[5\] VGND VGND VPWR VPWR _116_ _216_/a_59_75# sky130_fd_sc_hd__and2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_180_ net9 r2r_out[7] VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__nor2_1
X_301_ net9 VGND VGND VPWR VPWR _054_ _301_/a_27_47# sky130_fd_sc_hd__buf_2
X_163_ _066_ net4 _073_ _074_ _060_ VGND VGND VPWR VPWR _075_ _163_/a_193_297# _163_/a_109_297#
+ _163_/a_27_47# sky130_fd_sc_hd__a221o_1
X_232_ counter\[10\] _126_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_215_ counter\[7\] _112_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__nor2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_300_ _052_ VGND VGND VPWR VPWR _053_ _300_/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_231_ _066_ net15 VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__nand2_1
Xinput1 data[0] VGND VGND VPWR VPWR net1 input1/a_27_47# sky130_fd_sc_hd__buf_1
X_214_ _111_ _114_ _149_ VGND VGND VPWR VPWR _023_ _214_/a_113_297# sky130_fd_sc_hd__a21oi_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_230_ _065_ _127_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__nor2_1
Xinput2 data[1] VGND VGND VPWR VPWR net2 input2/a_27_47# sky130_fd_sc_hd__buf_1
X_213_ _112_ _052_ _113_ VGND VGND VPWR VPWR _114_ _213_/a_215_53# _213_/a_109_93#
+ sky130_fd_sc_hd__or3b_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput3 data[2] VGND VGND VPWR VPWR net3 input3/a_27_47# sky130_fd_sc_hd__buf_1
X_289_ divider\[4\] _041_ counter\[13\] _155_ VGND VGND VPWR VPWR _042_ _289_/a_489_413#
+ _289_/a_226_47# _289_/a_76_199# sky130_fd_sc_hd__a2bb2o_1
X_212_ counter\[5\] counter\[4\] _101_ counter\[6\] VGND VGND VPWR VPWR _113_ _212_/a_80_21#
+ _212_/a_209_297# sky130_fd_sc_hd__a31o_1
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 data[3] VGND VGND VPWR VPWR net4 input4/a_27_47# sky130_fd_sc_hd__buf_1
X_357_ clknet_2_3__leaf_clk net12 _000_ VGND VGND VPWR VPWR rst _357_/a_543_47# _357_/a_193_47#
+ _357_/a_448_47# _357_/a_1283_21# _357_/a_761_289# _357_/a_1108_47# _357_/a_27_47#
+ sky130_fd_sc_hd__dfrtp_2
X_288_ counter\[12\] VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__inv_2
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk clkbuf_2_1__f_clk/a_110_47#
+ sky130_fd_sc_hd__clkbuf_16
X_211_ counter\[6\] counter\[5\] counter\[4\] _101_ VGND VGND VPWR VPWR _112_ _211_/a_27_47#
+ sky130_fd_sc_hd__and4_1
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 data[4] VGND VGND VPWR VPWR net5 input5/a_27_47# sky130_fd_sc_hd__buf_1
XFILLER_0_23_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_356_ clknet_2_3__leaf_clk _032_ VGND VGND VPWR VPWR counter\[15\] _356_/a_891_413#
+ _356_/a_466_413# _356_/a_1059_315# _356_/a_193_47# _356_/a_634_159# _356_/a_381_47#
+ _356_/a_27_47# sky130_fd_sc_hd__dfxtp_1
X_287_ _037_ _038_ _039_ VGND VGND VPWR VPWR _040_ _287_/a_215_53# _287_/a_109_93#
+ sky130_fd_sc_hd__or3b_1
X_210_ _066_ net13 VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__nand2_1
X_339_ clknet_2_3__leaf_clk _015_ VGND VGND VPWR VPWR r2r_out[6] _339_/a_891_413#
+ _339_/a_193_47# _339_/a_381_47# _339_/a_1062_300# _339_/a_475_413# _339_/a_634_183#
+ _339_/a_27_47# sky130_fd_sc_hd__dfxtp_4
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_357__12 VGND VGND VPWR VPWR net12 _357__12/LO sky130_fd_sc_hd__conb_1
X_286_ divider\[6\] counter\[14\] VGND VGND VPWR VPWR _039_ _286_/a_27_53# _286_/a_219_297#
+ sky130_fd_sc_hd__or2b_1
X_355_ clknet_2_3__leaf_clk _031_ VGND VGND VPWR VPWR counter\[14\] _355_/a_891_413#
+ _355_/a_466_413# _355_/a_1059_315# _355_/a_193_47# _355_/a_634_159# _355_/a_381_47#
+ _355_/a_27_47# sky130_fd_sc_hd__dfxtp_1
Xinput6 data[5] VGND VGND VPWR VPWR net6 input6/a_27_47# sky130_fd_sc_hd__buf_1
XFILLER_0_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_269_ _148_ net5 _154_ VGND VGND VPWR VPWR _005_ _269_/a_215_297# _269_/a_27_413#
+ _269_/a_298_297# sky130_fd_sc_hd__a21bo_1
XFILLER_0_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_338_ clknet_2_3__leaf_clk _014_ VGND VGND VPWR VPWR r2r_out[5] _338_/a_891_413#
+ _338_/a_193_47# _338_/a_381_47# _338_/a_1062_300# _338_/a_475_413# _338_/a_634_183#
+ _338_/a_27_47# sky130_fd_sc_hd__dfxtp_4
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_285_ counter\[15\] divider\[7\] VGND VGND VPWR VPWR _038_ _285_/a_285_297# _285_/a_35_297#
+ sky130_fd_sc_hd__xor2_1
X_354_ clknet_2_2__leaf_clk _030_ VGND VGND VPWR VPWR counter\[13\] _354_/a_891_413#
+ _354_/a_466_413# _354_/a_1059_315# _354_/a_193_47# _354_/a_634_159# _354_/a_381_47#
+ _354_/a_27_47# sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput7 data[6] VGND VGND VPWR VPWR net7 input7/a_27_47# sky130_fd_sc_hd__buf_1
XFILLER_0_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_268_ net10 rst divider\[4\] VGND VGND VPWR VPWR _154_ _268_/a_215_53# _268_/a_109_93#
+ sky130_fd_sc_hd__or3b_1
X_337_ clknet_2_3__leaf_clk _013_ VGND VGND VPWR VPWR r2r_out[4] _337_/a_891_413#
+ _337_/a_193_47# _337_/a_381_47# _337_/a_1062_300# _337_/a_475_413# _337_/a_634_183#
+ _337_/a_27_47# sky130_fd_sc_hd__dfxtp_4
X_199_ net16 VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput10 load_divider VGND VGND VPWR VPWR net10 input10/a_27_47# sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_284_ counter\[14\] divider\[6\] VGND VGND VPWR VPWR _037_ _284_/a_27_413# _284_/a_207_413#
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_17_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_353_ clknet_2_1__leaf_clk _029_ VGND VGND VPWR VPWR counter\[12\] _353_/a_891_413#
+ _353_/a_466_413# _353_/a_1059_315# _353_/a_193_47# _353_/a_634_159# _353_/a_381_47#
+ _353_/a_27_47# sky130_fd_sc_hd__dfxtp_1
Xinput8 data[7] VGND VGND VPWR VPWR net8 input8/a_27_47# sky130_fd_sc_hd__buf_1
XFILLER_0_20_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_267_ _148_ net4 _153_ VGND VGND VPWR VPWR _004_ _267_/a_215_297# _267_/a_27_413#
+ _267_/a_298_297# sky130_fd_sc_hd__a21bo_1
X_336_ clknet_2_3__leaf_clk _012_ VGND VGND VPWR VPWR r2r_out[3] _336_/a_891_413#
+ _336_/a_193_47# _336_/a_381_47# _336_/a_1062_300# _336_/a_475_413# _336_/a_634_183#
+ _336_/a_27_47# sky130_fd_sc_hd__dfxtp_4
X_198_ counter\[3\] _097_ VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput11 n_rst VGND VGND VPWR VPWR net11 input11/a_75_212# sky130_fd_sc_hd__clkbuf_1
X_319_ net9 _068_ _069_ VGND VGND VPWR VPWR _070_ _319_/a_29_53# sky130_fd_sc_hd__or3_1
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 ext_data VGND VGND VPWR VPWR net9 input9/a_27_47# sky130_fd_sc_hd__clkbuf_2
X_283_ _035_ divider\[3\] divider\[2\] _159_ VGND VGND VPWR VPWR _036_ _283_/a_78_199#
+ _283_/a_215_47# sky130_fd_sc_hd__o22a_1
X_352_ clknet_2_2__leaf_clk _028_ VGND VGND VPWR VPWR counter\[11\] _352_/a_891_413#
+ _352_/a_466_413# _352_/a_1059_315# _352_/a_193_47# _352_/a_634_159# _352_/a_381_47#
+ _352_/a_27_47# sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_266_ net10 rst divider\[3\] VGND VGND VPWR VPWR _153_ _266_/a_215_53# _266_/a_109_93#
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_197_ counter\[3\] counter\[2\] counter\[1\] counter\[0\] VGND VGND VPWR VPWR _101_
+ _197_/a_27_47# sky130_fd_sc_hd__and4_2
X_335_ clknet_2_1__leaf_clk _011_ VGND VGND VPWR VPWR r2r_out[2] _335_/a_891_413#
+ _335_/a_193_47# _335_/a_381_47# _335_/a_1062_300# _335_/a_475_413# _335_/a_634_183#
+ _335_/a_27_47# sky130_fd_sc_hd__dfxtp_4
XFILLER_0_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_249_ _065_ _142_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_318_ r2r_out[2] r2r_out[1] r2r_out[0] VGND VGND VPWR VPWR _069_ _318_/a_27_47# sky130_fd_sc_hd__and3_1
Xhold1 counter\[6\] VGND VGND VPWR VPWR net13 hold1/a_49_47# hold1/a_285_47# hold1/a_391_47#
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_282_ counter\[11\] VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_351_ clknet_2_0__leaf_clk _027_ VGND VGND VPWR VPWR counter\[10\] _351_/a_891_413#
+ _351_/a_466_413# _351_/a_1059_315# _351_/a_193_47# _351_/a_634_159# _351_/a_381_47#
+ _351_/a_27_47# sky130_fd_sc_hd__dfxtp_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ clknet_2_1__leaf_clk _010_ VGND VGND VPWR VPWR r2r_out[1] _334_/a_891_413#
+ _334_/a_193_47# _334_/a_381_47# _334_/a_1062_300# _334_/a_475_413# _334_/a_634_183#
+ _334_/a_27_47# sky130_fd_sc_hd__dfxtp_4
X_265_ _148_ net3 _152_ VGND VGND VPWR VPWR _003_ _265_/a_215_297# _265_/a_27_413#
+ _265_/a_298_297# sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_196_ _065_ _100_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_179_ r2r_out[6] _053_ _087_ _057_ VGND VGND VPWR VPWR _015_ _179_/a_215_47# _179_/a_79_21#
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_248_ _094_ _140_ _141_ _046_ _078_ VGND VGND VPWR VPWR _142_ _248_/a_227_47# _248_/a_77_199#
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_317_ r2r_out[1] r2r_out[0] r2r_out[2] VGND VGND VPWR VPWR _068_ _317_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk clkbuf_2_2__f_clk/a_110_47#
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 counter\[4\] VGND VGND VPWR VPWR net14 hold2/a_49_47# hold2/a_285_47# hold2/a_391_47#
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_281_ _159_ divider\[2\] _160_ _161_ _033_ VGND VGND VPWR VPWR _034_ _281_/a_193_297#
+ _281_/a_109_297# _281_/a_27_47# sky130_fd_sc_hd__a221o_1
X_350_ clknet_2_0__leaf_clk _026_ VGND VGND VPWR VPWR counter\[9\] _350_/a_891_413#
+ _350_/a_466_413# _350_/a_1059_315# _350_/a_193_47# _350_/a_634_159# _350_/a_381_47#
+ _350_/a_27_47# sky130_fd_sc_hd__dfxtp_1
X_264_ net10 _149_ divider\[2\] VGND VGND VPWR VPWR _152_ _264_/a_215_53# _264_/a_109_93#
+ sky130_fd_sc_hd__or3b_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_195_ _094_ _097_ _098_ _099_ _078_ VGND VGND VPWR VPWR _100_ _195_/a_227_47# _195_/a_77_199#
+ sky130_fd_sc_hd__o32a_1
X_333_ clknet_2_1__leaf_clk _009_ VGND VGND VPWR VPWR r2r_out[0] _333_/a_891_413#
+ _333_/a_193_47# _333_/a_381_47# _333_/a_1062_300# _333_/a_475_413# _333_/a_634_183#
+ _333_/a_27_47# sky130_fd_sc_hd__dfxtp_4
XFILLER_0_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_316_ _066_ net3 VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__nand2_1
X_247_ counter\[13\] counter\[12\] _133_ VGND VGND VPWR VPWR _141_ _247_/a_27_47#
+ sky130_fd_sc_hd__and3_1
X_178_ _078_ _084_ _085_ _060_ _086_ VGND VGND VPWR VPWR _087_ _178_/a_75_199# _178_/a_201_297#
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3 counter\[10\] VGND VGND VPWR VPWR net15 hold3/a_49_47# hold3/a_285_47# hold3/a_391_47#
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_280_ counter\[9\] divider\[1\] VGND VGND VPWR VPWR _033_ _280_/a_27_413# _280_/a_207_413#
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_263_ _148_ net2 _151_ VGND VGND VPWR VPWR _002_ _263_/a_215_297# _263_/a_27_413#
+ _263_/a_298_297# sky130_fd_sc_hd__a21bo_1
X_332_ clknet_2_2__leaf_clk _008_ VGND VGND VPWR VPWR divider\[7\] _332_/a_891_413#
+ _332_/a_466_413# _332_/a_1059_315# _332_/a_193_47# _332_/a_634_159# _332_/a_381_47#
+ _332_/a_27_47# sky130_fd_sc_hd__dfxtp_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_194_ net17 VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_177_ _054_ net7 VGND VGND VPWR VPWR _086_ _177_/a_59_75# sky130_fd_sc_hd__and2_1
X_315_ net9 VGND VGND VPWR VPWR _066_ _315_/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_246_ counter\[12\] _133_ counter\[13\] VGND VGND VPWR VPWR _140_ _246_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_229_ _094_ _125_ _126_ _124_ _078_ VGND VGND VPWR VPWR _127_ _229_/a_227_47# _229_/a_77_199#
+ sky130_fd_sc_hd__o32a_1
Xhold4 counter\[3\] VGND VGND VPWR VPWR net16 hold4/a_49_47# hold4/a_285_47# hold4/a_391_47#
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ clknet_2_2__leaf_clk _007_ VGND VGND VPWR VPWR divider\[6\] _331_/a_891_413#
+ _331_/a_466_413# _331_/a_1059_315# _331_/a_193_47# _331_/a_634_159# _331_/a_381_47#
+ _331_/a_27_47# sky130_fd_sc_hd__dfxtp_1
X_262_ _148_ _149_ divider\[1\] VGND VGND VPWR VPWR _151_ _262_/a_215_53# _262_/a_109_93#
+ sky130_fd_sc_hd__or3b_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_193_ counter\[1\] counter\[0\] counter\[2\] VGND VGND VPWR VPWR _098_ _193_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_176_ r2r_out[6] _081_ VGND VGND VPWR VPWR _085_ _176_/a_68_297# sky130_fd_sc_hd__or2_1
XFILLER_0_3_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_314_ _061_ _064_ _065_ VGND VGND VPWR VPWR _010_ _314_/a_113_297# sky130_fd_sc_hd__a21oi_1
X_245_ _139_ VGND VGND VPWR VPWR _029_ _245_/a_75_212# sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_228_ counter\[9\] counter\[8\] _117_ VGND VGND VPWR VPWR _126_ _228_/a_27_47# sky130_fd_sc_hd__and3_1
Xhold5 counter\[2\] VGND VGND VPWR VPWR net17 hold5/a_49_47# hold5/a_285_47# hold5/a_391_47#
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_261_ _148_ net1 _150_ VGND VGND VPWR VPWR _001_ _261_/a_215_297# _261_/a_27_413#
+ _261_/a_298_297# sky130_fd_sc_hd__a21bo_1
X_330_ clknet_2_2__leaf_clk _006_ VGND VGND VPWR VPWR divider\[5\] _330_/a_891_413#
+ _330_/a_466_413# _330_/a_1059_315# _330_/a_193_47# _330_/a_634_159# _330_/a_381_47#
+ _330_/a_27_47# sky130_fd_sc_hd__dfxtp_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_192_ counter\[2\] counter\[1\] counter\[0\] VGND VGND VPWR VPWR _097_ _192_/a_27_47#
+ sky130_fd_sc_hd__and3_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_175_ r2r_out[6] _081_ VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__nand2_1
X_313_ _149_ VGND VGND VPWR VPWR _065_ _313_/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_244_ _057_ _138_ VGND VGND VPWR VPWR _139_ _244_/a_59_75# sky130_fd_sc_hd__and2_1
XFILLER_0_3_84 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_227_ _124_ _121_ VGND VGND VPWR VPWR _125_ _227_/a_59_75# sky130_fd_sc_hd__and2_1
XFILLER_0_20_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold6 counter\[7\] VGND VGND VPWR VPWR net18 hold6/a_49_47# hold6/a_285_47# hold6/a_391_47#
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_83 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_260_ _148_ _149_ divider\[0\] VGND VGND VPWR VPWR _150_ _260_/a_215_53# _260_/a_109_93#
+ sky130_fd_sc_hd__or3b_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_191_ _065_ _096_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_174_ r2r_out[5] _053_ _083_ _057_ VGND VGND VPWR VPWR _014_ _174_/a_215_47# _174_/a_79_21#
+ sky130_fd_sc_hd__o211a_1
X_312_ _053_ _063_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__nand2_1
X_243_ _059_ _135_ _137_ counter\[12\] _054_ VGND VGND VPWR VPWR _138_ _243_/a_93_21#
+ _243_/a_250_297# sky130_fd_sc_hd__a32o_1
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_226_ counter\[9\] VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__inv_2
Xhold7 counter\[0\] VGND VGND VPWR VPWR net19 hold7/a_49_47# hold7/a_285_47# hold7/a_391_47#
+ sky130_fd_sc_hd__dlygate4sd3_1
X_209_ _065_ _110_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_190_ _066_ counter\[1\] _094_ _095_ VGND VGND VPWR VPWR _096_ _190_/a_489_47# _190_/a_206_369#
+ _190_/a_76_199# sky130_fd_sc_hd__o2bb2a_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_173_ _066_ net6 _080_ _082_ _060_ VGND VGND VPWR VPWR _083_ _173_/a_193_297# _173_/a_109_297#
+ _173_/a_27_47# sky130_fd_sc_hd__a221o_1
X_242_ counter\[12\] _136_ VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__nand2_1
X_311_ _054_ net2 _062_ r2r_out[0] VGND VGND VPWR VPWR _063_ _311_/a_27_297# _311_/a_109_297#
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_225_ _123_ VGND VGND VPWR VPWR _025_ _225_/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xhold8 counter\[15\] VGND VGND VPWR VPWR net20 hold8/a_49_47# hold8/a_285_47# hold8/a_391_47#
+ sky130_fd_sc_hd__dlygate4sd3_1
X_208_ _066_ counter\[5\] _094_ _109_ VGND VGND VPWR VPWR _110_ _208_/a_489_47# _208_/a_206_369#
+ _208_/a_76_199# sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk clkbuf_2_3__f_clk/a_110_47#
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_310_ _054_ r2r_out[1] VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_172_ _054_ _081_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__nor2_1
X_241_ _117_ _132_ VGND VGND VPWR VPWR _136_ _241_/a_59_75# sky130_fd_sc_hd__and2_1
X_224_ _057_ _122_ VGND VGND VPWR VPWR _123_ _224_/a_59_75# sky130_fd_sc_hd__and2_1
Xhold9 r2r_out[2] VGND VGND VPWR VPWR net21 hold9/a_49_47# hold9/a_285_47# hold9/a_391_47#
+ sky130_fd_sc_hd__dlygate4sd3_1
X_207_ counter\[5\] _107_ VGND VGND VPWR VPWR _109_ _207_/a_285_297# _207_/a_35_297#
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_171_ r2r_out[5] r2r_out[4] _072_ VGND VGND VPWR VPWR _081_ _171_/a_27_47# sky130_fd_sc_hd__and3_1
X_240_ counter\[12\] _133_ VGND VGND VPWR VPWR _135_ _240_/a_68_297# sky130_fd_sc_hd__or2_1
X_223_ _059_ _120_ _121_ counter\[8\] _054_ VGND VGND VPWR VPWR _122_ _223_/a_93_21#
+ _223_/a_250_297# sky130_fd_sc_hd__a32o_1
XFILLER_0_20_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_206_ _105_ _108_ _149_ VGND VGND VPWR VPWR _021_ _206_/a_113_297# sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_170_ r2r_out[4] _072_ r2r_out[5] VGND VGND VPWR VPWR _080_ _170_/a_81_21# _170_/a_299_297#
+ sky130_fd_sc_hd__a21o_1
X_299_ _045_ _051_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__nand2_1
X_222_ counter\[8\] _117_ VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__nand2_1
X_205_ _106_ _094_ _107_ VGND VGND VPWR VPWR _108_ _205_/a_215_53# _205_/a_109_93#
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_298_ _040_ _047_ _043_ _050_ VGND VGND VPWR VPWR _051_ _298_/a_103_199# _298_/a_253_47#
+ sky130_fd_sc_hd__o31a_1
X_221_ counter\[8\] _117_ VGND VGND VPWR VPWR _120_ _221_/a_68_297# sky130_fd_sc_hd__or2_1
X_204_ counter\[4\] _101_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_297_ _038_ _039_ _048_ _049_ VGND VGND VPWR VPWR _050_ _297_/a_215_47# _297_/a_79_21#
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_220_ _065_ _119_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__nor2_1
X_349_ clknet_2_1__leaf_clk _025_ VGND VGND VPWR VPWR counter\[8\] _349_/a_891_413#
+ _349_/a_466_413# _349_/a_1059_315# _349_/a_193_47# _349_/a_634_159# _349_/a_381_47#
+ _349_/a_27_47# sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_203_ counter\[4\] _101_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_296_ divider\[7\] counter\[15\] VGND VGND VPWR VPWR _049_ _296_/a_27_53# _296_/a_219_297#
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_279_ counter\[8\] divider\[0\] VGND VGND VPWR VPWR _161_ _279_/a_27_413# _279_/a_207_413#
+ sky130_fd_sc_hd__and2b_1
X_348_ clknet_2_0__leaf_clk _024_ VGND VGND VPWR VPWR counter\[7\] _348_/a_891_413#
+ _348_/a_466_413# _348_/a_1059_315# _348_/a_193_47# _348_/a_634_159# _348_/a_381_47#
+ _348_/a_27_47# sky130_fd_sc_hd__dfxtp_1
X_202_ _066_ net14 VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_295_ net9 VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_278_ divider\[1\] counter\[9\] VGND VGND VPWR VPWR _160_ _278_/a_27_53# _278_/a_219_297#
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_347_ clknet_2_0__leaf_clk _023_ VGND VGND VPWR VPWR counter\[6\] _347_/a_891_413#
+ _347_/a_466_413# _347_/a_1059_315# _347_/a_193_47# _347_/a_634_159# _347_/a_381_47#
+ _347_/a_27_47# sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_201_ _065_ _104_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
C0 VGND _063_ 0.146062f
C1 VPWR _328_/a_891_413# 0.016847f
C2 VGND clk 4.037947f
C3 input6/a_27_47# VGND 0.055564f
C4 _326_/a_193_47# clknet_2_3__leaf_clk 0.076025f
C5 _097_ net16 0.024092f
C6 counter\[2\] _103_ 0.075823f
C7 _321_/a_79_199# _011_ 0.010436f
C8 _060_ _086_ 0.027901f
C9 clk _324_/a_68_297# 0.02138f
C10 _146_ counter\[15\] 0.011701f
C11 VGND clknet_2_0__leaf_clk 2.144026f
C12 _265_/a_27_413# rst 0.013943f
C13 _276_/a_27_413# _158_ 0.055787f
C14 _094_ _052_ 0.12104f
C15 _255_/a_209_297# _147_ 0.015261f
C16 _149_ _212_/a_209_297# 0.035149f
C17 counter\[14\] _252_/a_81_21# 0.059316f
C18 _200_/a_77_199# counter\[3\] 0.052994f
C19 _348_/a_27_47# _350_/a_193_47# 0.011595f
C20 counter\[10\] _131_ 0.017731f
C21 _290_/a_207_413# divider\[4\] 0.010223f
C22 divider\[4\] _005_ 0.024499f
C23 counter\[15\] _280_/a_207_413# 0.021114f
C24 _111_ _094_ 0.067078f
C25 _330_/a_891_413# _156_ 0.01252f
C26 _326_/a_891_413# _002_ 0.035426f
C27 _265_/a_215_297# _325_/a_27_47# 0.012332f
C28 _045_ net9 0.019611f
C29 _133_ counter\[11\] 0.06813f
C30 _112_ clknet_2_0__leaf_clk 0.015631f
C31 counter\[0\] hold7/a_49_47# 0.015863f
C32 _055_ _060_ 0.258446f
C33 VPWR _128_ 0.022934f
C34 VGND _130_ 0.053984f
C35 _339_/a_27_47# clknet_2_3__leaf_clk 0.02777f
C36 counter\[4\] hold2/a_285_47# 0.021182f
C37 _083_ _065_ 0.031953f
C38 r2r_out[1] _333_/a_634_183# 0.01755f
C39 _167_/a_27_47# _354_/a_1059_315# 0.01599f
C40 VPWR hold5/a_285_47# 0.010822f
C41 VGND hold5/a_391_47# -0.019265f
C42 _066_ _205_/a_215_53# 0.072574f
C43 _043_ _050_ 0.105707f
C44 VGND _033_ 0.169393f
C45 r2r_out[4] _170_/a_299_297# 0.05257f
C46 clknet_0_clk _159_ 0.022668f
C47 VPWR _059_ 0.21631f
C48 _057_ _338_/a_27_47# 0.040776f
C49 _253_/a_79_21# _145_ 0.129149f
C50 _060_ counter\[8\] 0.035506f
C51 _331_/a_27_47# rst 0.026911f
C52 _066_ _212_/a_80_21# 0.015662f
C53 _265_/a_27_413# VPWR 0.040236f
C54 _265_/a_215_297# VGND -0.01682f
C55 _060_ _143_ 0.050533f
C56 clknet_2_1__leaf_clk _095_ 0.013269f
C57 _060_ _141_ 0.13452f
C58 clknet_2_0__leaf_clk _052_ 0.428073f
C59 _066_ _094_ 1.580559f
C60 _065_ _344_/a_634_159# 0.035805f
C61 _016_ clknet_2_3__leaf_clk 0.270177f
C62 _149_ _153_ 0.178288f
C63 _097_ _102_ 0.13835f
C64 net8 _276_/a_298_297# 0.029765f
C65 _126_ _124_ 0.167996f
C66 counter\[15\] _033_ 0.14199f
C67 _306_/a_113_297# _009_ 0.04786f
C68 VPWR counter\[0\] 1.384349f
C69 VGND _097_ 0.828372f
C70 _251_/a_27_47# counter\[12\] 0.08015f
C71 _106_ _108_ 0.096698f
C72 _066_ _146_ 0.060354f
C73 _149_ _200_/a_77_199# 0.013978f
C74 _149_ counter\[6\] 1.205161f
C75 _340_/a_27_47# _340_/a_193_47# -0.035352f
C76 VPWR load_divider 0.220566f
C77 _326_/a_193_47# net2 0.034562f
C78 r2r_out[6] r2r_out[5] 0.018227f
C79 _004_ divider\[2\] 0.044694f
C80 data[4] data[3] 0.039867f
C81 counter\[4\] _216_/a_59_75# 0.028355f
C82 _057_ _349_/a_193_47# 0.021547f
C83 _081_ _091_ 0.291951f
C84 VGND _331_/a_193_47# 0.035545f
C85 VPWR _331_/a_27_47# -0.108132f
C86 _287_/a_215_53# _039_ 0.074271f
C87 divider\[6\] net7 0.030982f
C88 _149_ _054_ 0.160425f
C89 divider\[1\] _327_/a_27_47# 0.193197f
C90 _066_ clknet_2_0__leaf_clk 0.057953f
C91 _057_ _146_ 0.086548f
C92 _136_ counter\[8\] 0.050442f
C93 clknet_0_clk _349_/a_1059_315# 0.023482f
C94 VPWR _124_ 0.275662f
C95 _356_/a_891_413# counter\[15\] 0.045358f
C96 net22 clknet_2_3__leaf_clk 0.094001f
C97 VPWR counter\[1\] 0.85035f
C98 _066_ _130_ 0.266072f
C99 _035_ net9 0.016608f
C100 VGND _186_/a_113_297# 0.012842f
C101 _114_ _219_/a_227_47# 0.029606f
C102 _053_ _339_/a_475_413# 0.023967f
C103 _057_ clk 0.332578f
C104 counter\[6\] _065_ 0.042502f
C105 divider\[6\] _331_/a_466_413# 0.034189f
C106 _351_/a_27_47# _149_ 0.023944f
C107 clkbuf_0_clk/a_110_47# clk 0.011176f
C108 _185_/a_113_297# _088_ 0.019013f
C109 data[0] data[1] 0.04444f
C110 net4 net7 0.017397f
C111 net2 hold8/a_391_47# 0.017854f
C112 _353_/a_466_413# _029_ 0.031764f
C113 _347_/a_1059_315# _023_ 0.01848f
C114 _072_ r2r_out[5] 0.076733f
C115 _227_/a_59_75# _117_ 0.039951f
C116 net5 counter\[8\] 0.164759f
C117 data[5] _329_/a_1059_315# 0.011103f
C118 _054_ r2r_out[2] 0.015364f
C119 VGND divider\[4\] 1.986324f
C120 _154_ net5 0.282289f
C121 _053_ _015_ 0.074706f
C122 divider\[3\] divider\[4\] 0.640958f
C123 _173_/a_27_47# _082_ 0.012091f
C124 _065_ _054_ 0.036623f
C125 _148_ _005_ 0.106221f
C126 divider\[1\] _325_/a_27_47# 0.035013f
C127 divider\[6\] _007_ 0.028753f
C128 VGND _306_/a_113_297# 0.011664f
C129 _326_/a_891_413# VPWR 0.01622f
C130 _089_ _090_ 0.018477f
C131 VGND _131_ 0.015435f
C132 _328_/a_466_413# divider\[2\] 0.010348f
C133 _229_/a_77_199# _126_ 0.042123f
C134 _070_ VGND 0.059085f
C135 _072_ _077_ 0.074195f
C136 _336_/a_381_47# clk 0.014365f
C137 r2r_out[1] _064_ 0.01293f
C138 _354_/a_193_47# clknet_2_2__leaf_clk 0.061044f
C139 _078_ _317_/a_113_297# 0.017463f
C140 _149_ clknet_2_3__leaf_clk 0.073635f
C141 _072_ _163_/a_27_47# 0.010833f
C142 _336_/a_193_47# _336_/a_475_413# -0.01329f
C143 _150_ _260_/a_215_53# 0.028643f
C144 divider\[4\] counter\[15\] 0.022022f
C145 counter\[0\] _341_/a_466_413# 0.016781f
C146 _325_/a_193_47# _001_ 0.068156f
C147 net6 _082_ 0.086562f
C148 _353_/a_891_413# VPWR 0.026108f
C149 divider\[1\] VGND 0.390246f
C150 counter\[6\] hold1/a_391_47# 0.041796f
C151 _339_/a_1062_300# VPWR 0.086892f
C152 _339_/a_891_413# VGND 0.021634f
C153 _039_ _049_ 0.013717f
C154 rst net10 0.75068f
C155 VGND _327_/a_1059_315# -0.012212f
C156 _345_/a_891_413# _021_ 0.010793f
C157 _072_ net4 0.020169f
C158 _094_ counter\[9\] 0.0474f
C159 VPWR _229_/a_77_199# 0.045969f
C160 VPWR _357_/a_543_47# 0.03143f
C161 _154_ _156_ 0.010443f
C162 VPWR _354_/a_891_413# 0.011633f
C163 _352_/a_466_413# counter\[11\] 0.032536f
C164 VPWR _127_ 0.691097f
C165 VGND net20 0.368074f
C166 VPWR _001_ 0.69125f
C167 divider\[1\] counter\[15\] 0.19559f
C168 _244_/a_59_75# _138_ 0.046045f
C169 _281_/a_27_47# divider\[2\] 0.031499f
C170 r2r_out[4] _337_/a_27_47# 0.031184f
C171 VGND _352_/a_193_47# 0.022715f
C172 VPWR _352_/a_27_47# -0.154821f
C173 clknet_2_1__leaf_clk _019_ 0.074125f
C174 _149_ _067_ 0.160639f
C175 _332_/a_193_47# _158_ 0.081988f
C176 clknet_0_clk _115_ 0.021166f
C177 VPWR input9/a_27_47# 0.121733f
C178 _065_ clknet_2_3__leaf_clk 0.36436f
C179 _332_/a_27_47# clknet_2_2__leaf_clk 0.011922f
C180 _120_ _117_ 0.011156f
C181 _094_ _248_/a_77_199# 0.034794f
C182 VPWR net10 3.221557f
C183 VGND _158_ 0.541352f
C184 divider\[7\] _275_/a_215_53# 0.051707f
C185 _028_ counter\[11\] 0.11254f
C186 VPWR hold7/a_391_47# 0.014689f
C187 VPWR _272_/a_298_297# 0.011301f
C188 VPWR _029_ 0.143435f
C189 counter\[15\] net20 0.306059f
C190 input5/a_27_47# net10 0.013299f
C191 hold5/a_49_47# counter\[0\] 0.060404f
C192 _177_/a_59_75# _054_ 0.024705f
C193 VGND _091_ 0.240305f
C194 _149_ _261_/a_215_297# 0.035121f
C195 r2r_out[7] clknet_2_3__leaf_clk 0.111653f
C196 counter\[10\] _307_/a_59_75# 0.019268f
C197 _353_/a_1059_315# counter\[12\] 0.038541f
C198 net21 r2r_out[2] 0.165738f
C199 VPWR net18 0.13597f
C200 r2r_out[1] _056_ 0.091137f
C201 counter\[7\] _094_ 0.361295f
C202 net8 _272_/a_215_297# 0.029076f
C203 VPWR _325_/a_466_413# 0.033371f
C204 clkbuf_2_0__f_clk/a_110_47# _348_/a_1059_315# 0.011588f
C205 VGND hold2/a_49_47# 0.019244f
C206 _178_/a_75_199# net9 0.010803f
C207 _149_ net2 0.231368f
C208 _291_/a_193_297# divider\[3\] 0.060881f
C209 clknet_0_clk counter\[8\] 1.543968f
C210 _149_ net9 0.020068f
C211 _301_/a_27_47# net4 0.043481f
C212 r2r_out[3] clk 0.333198f
C213 _355_/a_1059_315# VGND -0.011715f
C214 clknet_0_clk _143_ 0.021772f
C215 _342_/a_634_159# clknet_2_1__leaf_clk 0.044335f
C216 _325_/a_634_159# net8 0.017414f
C217 clknet_0_clk _141_ 0.07864f
C218 counter\[15\] _158_ 0.02554f
C219 VPWR _332_/a_1059_315# 0.048113f
C220 VGND _332_/a_891_413# 0.024091f
C221 data[0] n_rst 0.041969f
C222 _333_/a_27_47# _058_ 0.031821f
C223 _160_ net4 0.161126f
C224 _348_/a_381_47# clknet_2_0__leaf_clk 0.028074f
C225 _298_/a_253_47# _043_ 0.012332f
C226 _355_/a_193_47# _031_ 0.219606f
C227 _146_ _147_ 0.062108f
C228 _045_ _133_ 0.07145f
C229 _051_ clkbuf_2_2__f_clk/a_110_47# 0.033617f
C230 counter\[2\] counter\[0\] 0.533085f
C231 VGND _020_ 0.023401f
C232 _010_ _053_ 0.061807f
C233 VGND _285_/a_35_297# 0.070791f
C234 _105_ VGND 0.732024f
C235 _273_/a_215_53# net9 0.042256f
C236 VGND _044_ 0.107102f
C237 data[4] VGND 0.066781f
C238 _136_ _308_/a_27_47# 0.022791f
C239 _031_ VPWR 0.256933f
C240 _284_/a_27_413# VPWR 0.041004f
C241 net6 _272_/a_215_297# 0.057489f
C242 _086_ _078_ 0.011061f
C243 input8/a_27_47# net10 0.036607f
C244 _148_ VGND 1.433401f
C245 counter\[1\] hold5/a_49_47# 0.030436f
C246 _330_/a_27_47# net10 0.041823f
C247 counter\[7\] clknet_2_0__leaf_clk 0.59486f
C248 counter\[10\] _132_ 0.019188f
C249 _123_ _117_ 0.023744f
C250 _139_ _245_/a_75_212# 0.119207f
C251 _149_ _260_/a_215_53# 0.031746f
C252 VPWR _223_/a_250_297# -0.023583f
C253 _008_ net8 0.064824f
C254 _325_/a_634_159# net6 0.045019f
C255 _285_/a_35_297# counter\[15\] 0.015171f
C256 _342_/a_193_47# _096_ 0.019131f
C257 _072_ r2r_out[4] 0.840807f
C258 _081_ _054_ 0.015093f
C259 counter\[10\] _054_ 0.021681f
C260 _334_/a_891_413# VGND 0.018037f
C261 _334_/a_1062_300# VPWR 0.078852f
C262 _096_ _018_ 0.038159f
C263 net9 _041_ 0.024115f
C264 _060_ net3 0.025781f
C265 VGND _211_/a_27_47# 0.035326f
C266 _339_/a_891_413# _057_ 0.015843f
C267 _112_ _213_/a_215_53# 0.029328f
C268 _101_ _021_ 0.014479f
C269 _048_ _038_ 0.09463f
C270 _053_ _068_ 0.031936f
C271 r2r_out[7] net9 0.04539f
C272 _053_ _333_/a_381_47# 0.017639f
C273 counter\[1\] counter\[2\] 0.129327f
C274 _094_ _126_ 0.70848f
C275 VPWR _338_/a_27_47# 0.109945f
C276 VGND _338_/a_193_47# -0.128825f
C277 _055_ _061_ 0.013341f
C278 VGND _083_ 0.812721f
C279 _296_/a_219_297# divider\[7\] 0.010497f
C280 VGND input2/a_27_47# 0.051016f
C281 _004_ net5 0.021601f
C282 data[7] VGND 0.068829f
C283 _078_ counter\[8\] 0.031515f
C284 VPWR _330_/a_634_159# 0.047289f
C285 VGND _140_ 0.070276f
C286 _057_ net20 0.03622f
C287 _356_/a_193_47# clknet_2_3__leaf_clk 0.012118f
C288 _351_/a_27_47# counter\[10\] 0.040928f
C289 _355_/a_381_47# net4 0.012458f
C290 _238_/a_77_199# _133_ 0.025075f
C291 _078_ _141_ 0.111576f
C292 _065_ _098_ 0.030936f
C293 VPWR _258_/a_27_47# 0.018409f
C294 VPWR _208_/a_206_369# 0.017932f
C295 _066_ hold2/a_49_47# 0.036705f
C296 _101_ _189_/a_47_47# 0.010835f
C297 net6 net8 1.404028f
C298 _031_ counter\[14\] 0.031399f
C299 _213_/a_215_53# _052_ 0.017168f
C300 _284_/a_27_413# counter\[14\] 0.052235f
C301 _338_/a_475_413# r2r_out[5] 0.035906f
C302 _124_ _228_/a_27_47# 0.12257f
C303 clknet_2_1__leaf_clk _056_ 0.186579f
C304 VGND _205_/a_109_93# -0.011421f
C305 _065_ clknet_2_2__leaf_clk 0.422051f
C306 _355_/a_1059_315# _066_ 0.054635f
C307 _247_/a_27_47# _141_ 0.014401f
C308 _101_ _115_ 0.171867f
C309 _104_ _344_/a_27_47# 0.075675f
C310 VGND _344_/a_634_159# -0.011934f
C311 VPWR _344_/a_193_47# 0.013919f
C312 _173_/a_27_47# net6 0.075446f
C313 hold6/a_49_47# _078_ 0.013981f
C314 hold6/a_285_47# _117_ 0.014989f
C315 VGND _006_ 0.137899f
C316 VPWR _252_/a_299_297# 0.038294f
C317 _066_ _170_/a_81_21# 0.014245f
C318 _264_/a_109_93# data[3] 0.046529f
C319 _094_ _107_ 0.085587f
C320 VPWR _212_/a_80_21# 0.050788f
C321 _343_/a_193_47# clknet_2_1__leaf_clk 0.012082f
C322 clk rst 0.029308f
C323 _035_ _133_ 0.032245f
C324 VPWR _349_/a_193_47# 0.053357f
C325 VGND _349_/a_634_159# 0.018238f
C326 VGND _328_/a_27_47# 0.043311f
C327 VPWR _094_ 5.55662f
C328 data[1] net1 0.098442f
C329 _105_ _066_ 0.087325f
C330 net14 _094_ 0.053885f
C331 _279_/a_27_413# _161_ 0.034503f
C332 _289_/a_76_199# _155_ 0.074181f
C333 _339_/a_27_47# r2r_out[6] 0.011509f
C334 _348_/a_193_47# _024_ 0.397559f
C335 _017_ clknet_2_1__leaf_clk 0.190512f
C336 VPWR _146_ 0.059768f
C337 VGND _307_/a_59_75# -0.013636f
C338 _329_/a_381_47# clknet_2_2__leaf_clk 0.015567f
C339 _355_/a_1059_315# clkbuf_0_clk/a_110_47# 0.010486f
C340 VPWR _347_/a_891_413# 0.018815f
C341 _330_/a_1059_315# _271_/a_29_53# 0.017378f
C342 _343_/a_891_413# counter\[2\] 0.045557f
C343 _326_/a_1059_315# _263_/a_215_297# 0.011113f
C344 _188_/a_27_47# _094_ 0.035825f
C345 net3 net1 0.530498f
C346 VPWR _063_ 0.39948f
C347 _142_ _078_ 0.04843f
C348 VPWR clk 1.272621f
C349 net5 net3 0.024335f
C350 input6/a_27_47# VPWR 0.117154f
C351 _326_/a_634_159# clknet_2_3__leaf_clk 0.042342f
C352 counter\[0\] _103_ 0.163285f
C353 VGND _345_/a_193_47# -0.093962f
C354 VPWR _345_/a_27_47# 0.106226f
C355 _142_ _051_ 0.022608f
C356 VGND _153_ 0.214394f
C357 _300_/a_27_47# _123_ 0.091967f
C358 _060_ _084_ 0.118091f
C359 _038_ net9 0.016247f
C360 VPWR clknet_2_0__leaf_clk 2.898062f
C361 _265_/a_215_297# rst 0.048947f
C362 _276_/a_215_297# _158_ 0.055569f
C363 _053_ counter\[0\] 0.365793f
C364 counter\[14\] _252_/a_299_297# 0.017811f
C365 _200_/a_77_199# _102_ 0.020827f
C366 _328_/a_891_413# net8 0.043914f
C367 _278_/a_219_297# counter\[8\] 0.014843f
C368 _094_ _116_ 0.059583f
C369 _114_ _094_ 0.021268f
C370 net17 _099_ 0.13486f
C371 VGND counter\[6\] 0.234437f
C372 divider\[1\] counter\[9\] 0.258728f
C373 _094_ counter\[13\] 0.081045f
C374 _149_ net15 0.010271f
C375 _326_/a_381_47# _002_ 0.012491f
C376 VGND _135_ 0.38272f
C377 _084_ _183_/a_59_75# 0.032398f
C378 _078_ _195_/a_77_199# 0.012911f
C379 _207_/a_35_297# counter\[4\] 0.064941f
C380 _229_/a_227_47# _078_ 0.014708f
C381 _052_ _307_/a_59_75# 0.039582f
C382 VGND _050_ 0.26142f
C383 VPWR _130_ 0.243716f
C384 r2r_out[1] r2r_out[2] 0.217401f
C385 _327_/a_27_47# clknet_2_3__leaf_clk 0.03716f
C386 r2r_out[1] _333_/a_475_413# 0.032848f
C387 VGND _132_ 0.371519f
C388 _149_ _266_/a_215_53# 0.074175f
C389 _167_/a_27_47# _354_/a_891_413# 0.01508f
C390 _192_/a_27_47# counter\[3\] 0.090961f
C391 _066_ _205_/a_109_93# 0.062403f
C392 _035_ divider\[5\] 0.396762f
C393 r2r_out[1] _065_ 0.549655f
C394 _115_ _217_/a_27_47# 0.022747f
C395 VPWR _033_ 0.418428f
C396 VGND _161_ 0.211945f
C397 _188_/a_27_47# clknet_2_0__leaf_clk 0.038687f
C398 _047_ clkbuf_2_2__f_clk/a_110_47# 0.011301f
C399 clknet_2_1__leaf_clk clkbuf_2_1__f_clk/a_110_47# 0.251474f
C400 _279_/a_27_413# clknet_2_3__leaf_clk 0.019731f
C401 _205_/a_215_53# _106_ 0.011896f
C402 VGND _054_ 3.209671f
C403 _057_ _338_/a_193_47# 0.034903f
C404 _114_ _347_/a_891_413# 0.01113f
C405 _155_ _035_ 0.113311f
C406 divider\[1\] _002_ 0.058176f
C407 clknet_2_3__leaf_clk _357_/a_27_47# 0.043672f
C408 VGND input11/a_75_212# 0.057444f
C409 _038_ clknet_2_2__leaf_clk 0.133756f
C410 _083_ _057_ 0.114038f
C411 _331_/a_193_47# rst 0.028116f
C412 _081_ net9 0.031176f
C413 _057_ _145_ 0.364824f
C414 _333_/a_27_47# _333_/a_193_47# -0.138648f
C415 net6 _328_/a_891_413# 0.049411f
C416 counter\[1\] _103_ 0.326659f
C417 _065_ _344_/a_466_413# 0.026552f
C418 _094_ _106_ 0.034493f
C419 _334_/a_27_47# clknet_2_1__leaf_clk 0.17825f
C420 _079_ _077_ 0.097999f
C421 VGND _225_/a_75_212# 0.030751f
C422 counter\[15\] _161_ 0.255821f
C423 _148_ _276_/a_215_297# 0.040917f
C424 VPWR _097_ 0.06687f
C425 _223_/a_93_21# _059_ 0.020844f
C426 counter\[15\] _054_ 0.386862f
C427 _111_ counter\[6\] 0.019439f
C428 _351_/a_27_47# VGND 0.047117f
C429 _065_ net15 0.184318f
C430 _052_ _132_ 0.76898f
C431 divider\[2\] net5 0.129092f
C432 VPWR _314_/a_113_297# 0.073257f
C433 _149_ clknet_2_1__leaf_clk 1.01968f
C434 _326_/a_193_47# _089_ 0.012561f
C435 _157_ divider\[6\] 0.244788f
C436 hold10/a_49_47# _340_/a_27_47# 0.010568f
C437 _069_ net9 0.183453f
C438 _325_/a_27_47# clknet_2_3__leaf_clk 0.037583f
C439 VGND _331_/a_634_159# 0.028627f
C440 data[0] net1 0.110148f
C441 _159_ _034_ 0.0898f
C442 _287_/a_109_93# _039_ 0.056863f
C443 _149_ _192_/a_27_47# 0.015537f
C444 hold6/a_49_47# _217_/a_27_47# 0.011328f
C445 clkbuf_2_0__f_clk/a_110_47# _065_ 0.010734f
C446 divider\[1\] _327_/a_193_47# 0.017241f
C447 _073_ _076_ 0.14138f
C448 input3/a_27_47# data[2] 0.042223f
C449 _048_ VGND 0.331322f
C450 net8 _331_/a_27_47# 0.030463f
C451 _084_ net5 0.073797f
C452 divider\[4\] _294_/a_215_47# 0.067693f
C453 counter\[12\] _059_ 0.420862f
C454 _005_ clknet_2_2__leaf_clk 0.070057f
C455 _071_ _060_ 0.039999f
C456 clknet_0_clk _349_/a_891_413# 0.013821f
C457 divider\[4\] rst 0.289305f
C458 VPWR _263_/a_298_297# -0.012723f
C459 r2r_out[6] _178_/a_75_199# 0.021549f
C460 counter\[6\] _066_ 0.386629f
C461 _356_/a_381_47# counter\[15\] 0.016707f
C462 _149_ net7 0.150753f
C463 r2r_out[6] _179_/a_215_47# 0.05007f
C464 _174_/a_79_21# r2r_out[5] 0.029276f
C465 VGND clknet_2_3__leaf_clk 3.185497f
C466 _043_ divider\[5\] 0.130559f
C467 VGND _243_/a_93_21# -0.010606f
C468 _075_ _054_ 0.06032f
C469 VPWR _186_/a_113_297# 0.028962f
C470 _066_ _132_ 0.084508f
C471 _148_ _269_/a_27_413# 0.059037f
C472 _010_ counter\[0\] 0.011514f
C473 divider\[6\] _331_/a_1059_315# 0.054629f
C474 VGND _164_/a_79_21# 0.031049f
C475 _347_/a_466_413# clknet_2_0__leaf_clk 0.010102f
C476 _066_ _054_ 0.252073f
C477 _040_ divider\[4\] 0.051467f
C478 clknet_2_1__leaf_clk _065_ 0.354056f
C479 _054_ r2r_out[0] 0.196846f
C480 _353_/a_1059_315# _029_ 0.022946f
C481 divider\[1\] rst 0.028984f
C482 _347_/a_891_413# _023_ 0.042121f
C483 counter\[15\] clknet_2_3__leaf_clk 0.098225f
C484 VPWR _264_/a_215_53# 0.010378f
C485 _289_/a_76_199# _159_ 0.017728f
C486 VPWR divider\[4\] 0.36245f
C487 _149_ _348_/a_27_47# 0.031757f
C488 divider\[1\] _259_/a_27_47# 0.011409f
C489 _060_ _183_/a_59_75# 0.02242f
C490 _062_ hold7/a_285_47# 0.012751f
C491 divider\[1\] _325_/a_193_47# 0.013677f
C492 VPWR _306_/a_113_297# 0.024355f
C493 _023_ clknet_2_0__leaf_clk 0.119329f
C494 VPWR _131_ 0.332294f
C495 _067_ VGND 0.10795f
C496 _357_/a_27_47# net12 0.089677f
C497 divider\[0\] _150_ 0.040677f
C498 _149_ divider\[5\] 0.206605f
C499 _057_ _054_ 0.064149f
C500 r2r_out[6] _065_ 0.150904f
C501 data[5] data[6] 0.038372f
C502 _149_ _155_ 0.089669f
C503 divider\[5\] _271_/a_29_53# 0.085347f
C504 counter\[0\] _341_/a_1059_315# 0.043378f
C505 _094_ _233_/a_80_21# 0.020387f
C506 VGND _261_/a_215_297# -0.014721f
C507 VPWR _261_/a_27_413# 0.014827f
C508 net4 counter\[8\] 0.338256f
C509 VGND _315_/a_27_47# 0.102808f
C510 divider\[4\] _294_/a_78_199# 0.040514f
C511 divider\[1\] VPWR 1.890574f
C512 input7/a_27_47# data[6] 0.018659f
C513 _339_/a_891_413# VPWR 0.022634f
C514 net4 _141_ 0.018341f
C515 _155_ _271_/a_29_53# 0.011095f
C516 VGND _327_/a_891_413# -0.012523f
C517 VPWR _327_/a_1059_315# 0.015904f
C518 _087_ clknet_2_3__leaf_clk 0.028503f
C519 _345_/a_381_47# _021_ 0.020213f
C520 VGND net2 0.850393f
C521 _075_ clknet_2_3__leaf_clk 0.026518f
C522 _322_/a_27_47# r2r_out[2] 0.026556f
C523 VGND net9 5.198038f
C524 VPWR _357_/a_1283_21# 0.051363f
C525 VGND _275_/a_215_53# 0.011567f
C526 _322_/a_27_47# _065_ 0.013882f
C527 _352_/a_1059_315# counter\[11\] 0.054539f
C528 _060_ _168_/a_76_199# 0.026582f
C529 VPWR net20 0.183421f
C530 _075_ _164_/a_79_21# 0.095463f
C531 _066_ clknet_2_3__leaf_clk 0.792184f
C532 r2r_out[4] _337_/a_193_47# 0.049609f
C533 VGND _352_/a_634_159# 0.011529f
C534 clknet_0_clk _123_ 0.090806f
C535 _297_/a_79_21# _038_ 0.101951f
C536 clknet_0_clk _117_ 0.032781f
C537 divider\[5\] _041_ 0.040199f
C538 _021_ counter\[4\] 0.202338f
C539 _001_ net8 0.025867f
C540 net2 counter\[15\] 0.020449f
C541 r2r_out[1] _069_ 0.057418f
C542 _053_ _031_ 0.085099f
C543 _072_ r2r_out[2] 0.026655f
C544 _013_ _054_ 0.062493f
C545 VGND _121_ 0.305333f
C546 _035_ _159_ 0.014795f
C547 counter\[15\] net9 0.033176f
C548 counter\[10\] net15 0.041251f
C549 _332_/a_193_47# clknet_2_2__leaf_clk 0.010618f
C550 _060_ net1 0.028158f
C551 _155_ _041_ 0.044531f
C552 VGND net12 0.193427f
C553 VPWR _158_ 0.359294f
C554 divider\[7\] _275_/a_109_93# 0.040613f
C555 counter\[15\] _275_/a_215_53# 0.042069f
C556 _072_ _065_ 1.140675f
C557 hold8/a_49_47# net5 0.019957f
C558 hold5/a_285_47# counter\[0\] 0.083586f
C559 VPWR _091_ 0.234927f
C560 _149_ _261_/a_298_297# 0.039513f
C561 VGND clknet_2_2__leaf_clk 1.437137f
C562 _149_ _313_/a_27_47# 0.01305f
C563 _107_ hold2/a_49_47# 0.040949f
C564 _011_ r2r_out[2] 0.10793f
C565 r2r_out[1] _009_ 0.02652f
C566 _057_ clknet_2_3__leaf_clk 0.071485f
C567 net8 net10 0.219289f
C568 net8 _272_/a_298_297# 0.03749f
C569 VPWR _325_/a_1059_315# 0.039655f
C570 VGND hold2/a_285_47# -0.019962f
C571 VPWR hold2/a_49_47# 0.0704f
C572 _148_ rst 0.717658f
C573 VPWR _291_/a_193_297# -0.012207f
C574 _152_ divider\[2\] 0.225472f
C575 _177_/a_59_75# net7 0.032883f
C576 r2r_out[6] _177_/a_59_75# 0.025634f
C577 _067_ _066_ 0.115731f
C578 _243_/a_93_21# clkbuf_0_clk/a_110_47# 0.011385f
C579 _355_/a_891_413# VGND -0.016129f
C580 _355_/a_1059_315# VPWR 0.041083f
C581 _057_ _164_/a_79_21# 0.045686f
C582 _342_/a_466_413# clknet_2_1__leaf_clk 0.038657f
C583 _325_/a_466_413# net8 0.034082f
C584 counter\[4\] _115_ 0.017123f
C585 _265_/a_215_297# _003_ 0.011577f
C586 VGND _332_/a_381_47# 0.019019f
C587 VPWR _332_/a_891_413# 0.024385f
C588 _107_ _109_ 0.011259f
C589 _027_ _234_/a_113_297# 0.019617f
C590 net6 _001_ 0.059531f
C591 _135_ counter\[9\] 0.025439f
C592 _053_ _338_/a_27_47# 0.035193f
C593 _040_ _044_ 0.045078f
C594 _057_ net21 0.024076f
C595 counter\[15\] clknet_2_2__leaf_clk 0.027563f
C596 VPWR _170_/a_81_21# 0.015739f
C597 VPWR _109_ 0.106522f
C598 counter\[2\] _097_ 0.112203f
C599 _105_ _107_ 0.568433f
C600 VGND _151_ 0.115633f
C601 _219_/a_77_199# _115_ 0.041099f
C602 _060_ _088_ 0.021898f
C603 _052_ _121_ 0.023286f
C604 VPWR _020_ 0.013304f
C605 VPWR _285_/a_35_297# 0.133504f
C606 counter\[9\] _132_ 0.280316f
C607 net14 _105_ 0.038009f
C608 _273_/a_109_93# net9 0.010163f
C609 _066_ _315_/a_27_47# 0.021171f
C610 _037_ clknet_2_2__leaf_clk 0.243044f
C611 data[4] VPWR 0.272521f
C612 input5/a_27_47# data[4] 0.021116f
C613 _149_ divider\[0\] 0.30791f
C614 _036_ _159_ 0.067957f
C615 _284_/a_207_413# VPWR 0.015082f
C616 net6 net10 0.054611f
C617 counter\[9\] _054_ 0.2161f
C618 _148_ VPWR 2.183699f
C619 net2 _066_ 0.032324f
C620 _330_/a_193_47# net10 0.01752f
C621 counter\[5\] _101_ 0.108779f
C622 counter\[1\] hold5/a_285_47# 0.031803f
C623 clkbuf_2_3__f_clk/a_110_47# _054_ 0.037071f
C624 _084_ _078_ 0.350756f
C625 _330_/a_634_159# _272_/a_215_297# 0.011552f
C626 _066_ net9 0.522709f
C627 net2 r2r_out[0] 0.227784f
C628 counter\[10\] _133_ 0.526751f
C629 _313_/a_27_47# _065_ 0.044294f
C630 _013_ clknet_2_3__leaf_clk 0.140756f
C631 _117_ _078_ 0.081225f
C632 _325_/a_466_413# net6 0.030431f
C633 _342_/a_27_47# _018_ 0.015636f
C634 VGND _216_/a_59_75# 0.024176f
C635 VGND _296_/a_219_297# 0.04662f
C636 _094_ _103_ 0.029611f
C637 _168_/a_76_199# net5 0.010901f
C638 _135_ _137_ 0.019501f
C639 _267_/a_215_297# _004_ 0.013142f
C640 _334_/a_891_413# VPWR 0.023035f
C641 _057_ _315_/a_27_47# 0.075011f
C642 _035_ _266_/a_109_93# 0.010538f
C643 VPWR _211_/a_27_47# -0.013054f
C644 _112_ _213_/a_109_93# 0.059298f
C645 _093_ clknet_2_1__leaf_clk 0.064943f
C646 counter\[7\] _132_ 0.148277f
C647 _081_ net7 0.015238f
C648 _081_ r2r_out[6] 0.783648f
C649 net2 _057_ 0.018343f
C650 counter\[1\] counter\[0\] 0.7063f
C651 VPWR _338_/a_193_47# 0.022056f
C652 VGND _338_/a_634_183# 0.015425f
C653 _328_/a_27_47# rst 0.015492f
C654 _057_ net9 1.226548f
C655 net5 net1 0.021943f
C656 VPWR _083_ 0.117462f
C657 net5 _268_/a_215_53# 0.011048f
C658 _296_/a_27_53# divider\[7\] 0.019049f
C659 _296_/a_219_297# counter\[15\] 0.018957f
C660 VPWR input2/a_27_47# 0.07875f
C661 net7 _005_ 0.019529f
C662 _073_ _074_ 0.042347f
C663 VPWR _145_ 0.028353f
C664 data[7] VPWR 0.226709f
C665 VPWR _330_/a_466_413# 0.037286f
C666 _338_/a_193_47# _014_ 0.060658f
C667 r2r_out[1] VGND 1.840297f
C668 VPWR _140_ 0.131749f
C669 _351_/a_193_47# counter\[10\] 0.168386f
C670 VGND _139_ 0.029831f
C671 _083_ _014_ 0.027094f
C672 _066_ hold2/a_285_47# 0.059139f
C673 clknet_0_clk _060_ 0.182593f
C674 _284_/a_207_413# counter\[14\] 0.072995f
C675 _045_ _141_ 0.023727f
C676 _338_/a_1062_300# r2r_out[5] 0.109691f
C677 _053_ _063_ 0.081998f
C678 _053_ clk 0.332027f
C679 clknet_2_1__leaf_clk _009_ 0.043562f
C680 _065_ _028_ 0.140168f
C681 _355_/a_891_413# _066_ 0.048006f
C682 r2r_out[7] _000_ 0.015401f
C683 _101_ _117_ 0.133394f
C684 _104_ _344_/a_193_47# 0.457464f
C685 VPWR _344_/a_634_159# 0.022027f
C686 _214_/a_113_297# _149_ 0.021266f
C687 _221_/a_68_297# _121_ 0.03246f
C688 hold6/a_49_47# _118_ 0.012537f
C689 hold6/a_285_47# _078_ 0.03811f
C690 VPWR _006_ 0.277461f
C691 VPWR _212_/a_209_297# -0.016209f
C692 _328_/a_891_413# net10 0.015289f
C693 VGND _349_/a_466_413# 0.019363f
C694 _094_ _104_ 0.183777f
C695 _116_ _211_/a_27_47# 0.073146f
C696 VGND _328_/a_193_47# -0.108159f
C697 VPWR _328_/a_27_47# -0.165587f
C698 _004_ net4 0.047622f
C699 _178_/a_75_199# _085_ 0.030343f
C700 _279_/a_207_413# _161_ 0.033315f
C701 clknet_2_1__leaf_clk net16 0.037187f
C702 VGND net15 0.365514f
C703 _060_ _076_ 0.256607f
C704 _105_ _106_ 0.010836f
C705 _289_/a_226_47# _155_ 0.030737f
C706 _163_/a_27_47# _073_ 0.042235f
C707 _348_/a_634_159# _024_ 0.045436f
C708 _290_/a_207_413# divider\[5\] 0.021484f
C709 r2r_out[3] _164_/a_79_21# 0.044248f
C710 VGND _266_/a_215_53# 0.026466f
C711 VPWR _307_/a_59_75# 0.019575f
C712 _002_ clknet_2_3__leaf_clk 0.718044f
C713 counter\[14\] _145_ 0.019889f
C714 _071_ _078_ 0.067766f
C715 _115_ _113_ 0.086182f
C716 input8/a_27_47# data[7] 0.013204f
C717 clknet_2_1__leaf_clk _195_/a_227_47# 0.011668f
C718 r2r_out[3] net21 0.171385f
C719 counter\[13\] _140_ 0.377101f
C720 _003_ divider\[1\] 0.147456f
C721 clknet_0_clk _136_ 0.362508f
C722 _055_ _056_ 0.142716f
C723 _343_/a_381_47# counter\[2\] 0.023071f
C724 _243_/a_93_21# _137_ 0.044675f
C725 _073_ net4 0.064013f
C726 _016_ _185_/a_113_297# 0.010455f
C727 _054_ rst 0.010967f
C728 _326_/a_466_413# clknet_2_3__leaf_clk 0.023464f
C729 VGND _297_/a_79_21# 0.036696f
C730 _159_ _041_ 0.120752f
C731 hold7/a_49_47# _054_ 0.012812f
C732 _097_ _103_ 0.18292f
C733 VPWR _345_/a_193_47# 0.050196f
C734 _321_/a_448_47# net21 0.017564f
C735 VPWR _153_ 0.134214f
C736 clknet_2_0__leaf_clk _104_ 0.165518f
C737 _276_/a_298_297# _158_ 0.01676f
C738 _241_/a_59_75# _132_ 0.03681f
C739 _063_ _303_/a_113_297# 0.012192f
C740 clknet_0_clk hold4/a_49_47# 0.020163f
C741 _330_/a_27_47# _006_ 0.060987f
C742 r2r_out[6] _176_/a_68_297# 0.042832f
C743 _328_/a_381_47# net8 0.016525f
C744 hold8/a_49_47# _078_ 0.027784f
C745 _348_/a_193_47# _350_/a_634_159# 0.010213f
C746 _021_ _206_/a_113_297# 0.010455f
C747 _060_ _078_ 0.412121f
C748 _032_ net1 0.021978f
C749 VPWR _200_/a_77_199# -0.010496f
C750 _040_ _050_ 0.138753f
C751 VPWR counter\[6\] 0.422092f
C752 divider\[1\] _263_/a_27_413# 0.031878f
C753 VPWR _135_ 0.078574f
C754 clkbuf_2_3__f_clk/a_110_47# _315_/a_27_47# 0.031894f
C755 _066_ _139_ 0.090311f
C756 r2r_out[1] r2r_out[0] 0.779843f
C757 _065_ _085_ 0.034753f
C758 _071_ _321_/a_79_199# 0.021399f
C759 _149_ input3/a_27_47# 0.028261f
C760 _208_/a_76_199# _094_ 0.010363f
C761 clknet_0_clk net1 0.024862f
C762 _060_ _061_ 0.054468f
C763 VPWR _050_ 0.133741f
C764 _344_/a_27_47# _344_/a_193_47# -0.012897f
C765 VGND clknet_2_1__leaf_clk 2.961549f
C766 _327_/a_193_47# clknet_2_3__leaf_clk 0.015585f
C767 r2r_out[1] _333_/a_1062_300# 0.036256f
C768 VGND _133_ 0.804776f
C769 VPWR _132_ 0.492004f
C770 _149_ _266_/a_109_93# 0.04863f
C771 counter\[9\] net9 0.017841f
C772 _035_ _141_ 0.030406f
C773 _192_/a_27_47# _102_ 0.044288f
C774 net2 clkbuf_2_3__f_clk/a_110_47# 0.012597f
C775 clkbuf_2_0__f_clk/a_110_47# _052_ 0.090304f
C776 net4 net3 0.083444f
C777 _117_ _217_/a_27_47# 0.065699f
C778 clkbuf_2_3__f_clk/a_110_47# net9 0.02401f
C779 VPWR _161_ 0.627149f
C780 VGND _192_/a_27_47# 0.020109f
C781 _094_ _344_/a_27_47# 0.431097f
C782 _279_/a_207_413# clknet_2_3__leaf_clk 0.013101f
C783 VPWR _054_ 2.439288f
C784 _205_/a_215_53# _108_ 0.050586f
C785 _057_ _338_/a_634_183# 0.023824f
C786 VPWR input11/a_75_212# 0.082894f
C787 _343_/a_891_413# counter\[1\] 0.011995f
C788 _331_/a_27_47# net10 0.0128f
C789 _112_ _133_ 0.173001f
C790 r2r_out[1] _057_ 0.075845f
C791 net6 _328_/a_381_47# 0.027609f
C792 data[1] data[2] 0.035937f
C793 input1/a_27_47# VPWR 0.058131f
C794 _089_ _081_ 0.027504f
C795 _057_ _139_ 0.015046f
C796 _065_ _344_/a_1059_315# 0.035727f
C797 _320_/a_80_21# _319_/a_29_53# 0.017174f
C798 VGND net7 1.191676f
C799 _066_ net15 0.015376f
C800 net2 _002_ 0.357281f
C801 counter\[9\] _121_ 0.017027f
C802 VGND r2r_out[6] 1.576122f
C803 _334_/a_193_47# clknet_2_1__leaf_clk 0.257015f
C804 _094_ _108_ 0.028852f
C805 _053_ _186_/a_113_297# 0.053871f
C806 _274_/a_215_297# _148_ 0.067621f
C807 VPWR _225_/a_75_212# 0.069601f
C808 _101_ _197_/a_27_47# 0.022208f
C809 _223_/a_250_297# _059_ 0.011116f
C810 _136_ _078_ 0.025891f
C811 counter\[6\] _116_ 0.150789f
C812 _351_/a_27_47# VPWR -0.091195f
C813 _351_/a_193_47# VGND -0.078904f
C814 rst clknet_2_3__leaf_clk 0.051745f
C815 _052_ _133_ 0.870678f
C816 clkbuf_2_0__f_clk/a_110_47# _066_ 0.011384f
C817 _149_ _021_ 0.139678f
C818 _046_ net9 0.053171f
C819 _325_/a_193_47# clknet_2_3__leaf_clk 0.038017f
C820 VGND _331_/a_466_413# 0.010513f
C821 net4 _281_/a_27_47# 0.018477f
C822 _040_ _048_ 0.029276f
C823 _152_ net5 0.162976f
C824 _322_/a_27_47# VGND 0.033724f
C825 _053_ _306_/a_113_297# 0.013238f
C826 _348_/a_27_47# VGND 0.094131f
C827 _355_/a_193_47# clknet_2_3__leaf_clk 0.010604f
C828 _073_ r2r_out[4] 0.018508f
C829 _053_ _070_ 0.13302f
C830 _048_ VPWR 0.27452f
C831 net8 _331_/a_193_47# 0.032963f
C832 _340_/a_27_47# _016_ 0.151506f
C833 _286_/a_219_297# VPWR 0.015104f
C834 _078_ net1 0.048695f
C835 _086_ _178_/a_75_199# 0.011822f
C836 _142_ _354_/a_193_47# 0.041693f
C837 _063_ _341_/a_1059_315# 0.030999f
C838 r2r_out[6] _178_/a_201_297# 0.045932f
C839 VGND divider\[5\] 0.54941f
C840 _078_ net5 0.225497f
C841 _149_ _189_/a_47_47# 0.011832f
C842 divider\[3\] divider\[5\] 0.029486f
C843 _092_ clknet_2_3__leaf_clk 0.229051f
C844 counter\[5\] _110_ 0.260286f
C845 VPWR clknet_2_3__leaf_clk 3.01035f
C846 VGND _012_ 0.220444f
C847 VGND _007_ 0.120806f
C848 net4 divider\[2\] 0.129852f
C849 _005_ _329_/a_27_47# 0.034356f
C850 _072_ VGND 0.625449f
C851 VGND _155_ 0.211684f
C852 divider\[3\] _155_ 0.626393f
C853 _014_ clknet_2_3__leaf_clk 0.069486f
C854 _235_/a_113_297# counter\[11\] 0.066054f
C855 _148_ _263_/a_27_413# 0.031696f
C856 _291_/a_27_47# divider\[4\] 0.047977f
C857 _066_ _133_ 0.024215f
C858 _148_ _269_/a_215_297# 0.054529f
C859 clknet_2_1__leaf_clk r2r_out[0] 0.288495f
C860 divider\[6\] _331_/a_891_413# 0.039957f
C861 _246_/a_113_297# _078_ 0.017375f
C862 VPWR _164_/a_79_21# 0.063775f
C863 net4 input4/a_27_47# 0.034296f
C864 _336_/a_27_47# _057_ 0.033351f
C865 r2r_out[6] _087_ 0.420811f
C866 _060_ net19 0.275716f
C867 divider\[2\] _283_/a_215_47# 0.012189f
C868 _080_ clknet_2_3__leaf_clk 0.0406f
C869 counter\[15\] divider\[5\] 0.025958f
C870 VPWR net21 0.040524f
C871 VGND _011_ 0.223353f
C872 _021_ _065_ 0.017227f
C873 _353_/a_891_413# _029_ 0.050984f
C874 _347_/a_381_47# _023_ 0.019683f
C875 _289_/a_226_47# _159_ 0.01071f
C876 counter\[15\] _155_ 0.022954f
C877 VGND _138_ 0.231101f
C878 _149_ _348_/a_193_47# 0.033306f
C879 net2 rst 0.026151f
C880 counter\[10\] _159_ 0.014939f
C881 _327_/a_193_47# clknet_2_2__leaf_clk 0.031969f
C882 rst net9 0.19174f
C883 _057_ clknet_2_1__leaf_clk 0.204903f
C884 _057_ _337_/a_27_47# 0.062969f
C885 _048_ counter\[14\] 0.026089f
C886 _067_ VPWR 0.014724f
C887 _094_ counter\[0\] 0.138159f
C888 _048_ counter\[13\] 0.2215f
C889 divider\[4\] net8 0.024747f
C890 _134_ _028_ 0.025891f
C891 net2 _259_/a_27_47# 0.024317f
C892 _122_ _054_ 0.030931f
C893 _354_/a_466_413# clknet_2_2__leaf_clk 0.011003f
C894 _081_ _085_ 0.222212f
C895 counter\[0\] _341_/a_891_413# 0.047848f
C896 net10 input9/a_27_47# 0.062696f
C897 r2r_out[1] r2r_out[3] 0.209547f
C898 VPWR _261_/a_215_297# 0.018537f
C899 VPWR _315_/a_27_47# 0.132032f
C900 _096_ _065_ 0.08344f
C901 _160_ VGND 0.207459f
C902 VGND _313_/a_27_47# 0.077187f
C903 _025_ _349_/a_381_47# 0.022668f
C904 _040_ net9 0.041737f
C905 _057_ r2r_out[6] 0.312869f
C906 _128_ _130_ 0.11988f
C907 _353_/a_27_47# net1 0.033382f
C908 _345_/a_1059_315# counter\[4\] 0.056512f
C909 counter\[13\] _248_/a_227_47# 0.087546f
C910 VPWR net2 0.888041f
C911 divider\[1\] net8 0.017618f
C912 _075_ _012_ 0.056474f
C913 counter\[5\] counter\[4\] 1.306232f
C914 _060_ _074_ 0.137673f
C915 rst clknet_2_2__leaf_clk 0.3064f
C916 VPWR net9 2.854717f
C917 _030_ clknet_2_2__leaf_clk 0.275593f
C918 counter\[0\] _063_ 0.266672f
C919 _072_ _075_ 0.090828f
C920 _094_ _124_ 0.252935f
C921 _089_ VGND 0.317702f
C922 VPWR _357_/a_1108_47# 0.030347f
C923 VGND _275_/a_109_93# 0.01083f
C924 _148_ _327_/a_634_159# 0.011722f
C925 net6 divider\[4\] 0.072318f
C926 _346_/a_27_47# _065_ 0.051335f
C927 _352_/a_891_413# counter\[11\] 0.039792f
C928 _160_ counter\[15\] 0.016374f
C929 _100_ _019_ 0.368409f
C930 _325_/a_193_47# clknet_2_2__leaf_clk 0.010626f
C931 r2r_out[4] _337_/a_634_183# 0.010685f
C932 _013_ _337_/a_27_47# 0.173165f
C933 VPWR _352_/a_634_159# 0.016833f
C934 _195_/a_77_199# clkbuf_2_1__f_clk/a_110_47# 0.012339f
C935 clknet_0_clk _025_ 0.03367f
C936 counter\[1\] _094_ 0.353925f
C937 _141_ _041_ 0.078521f
C938 _332_/a_466_413# _158_ 0.019512f
C939 clknet_0_clk _078_ 0.112528f
C940 _072_ r2r_out[0] 0.016355f
C941 VGND ext_data 0.062787f
C942 hold4/a_391_47# _195_/a_77_199# 0.014107f
C943 _240_/a_68_297# _078_ 0.013963f
C944 VPWR _121_ 0.049571f
C945 _305_/a_27_47# VGND -0.011925f
C946 _151_ rst 0.013013f
C947 divider\[0\] VGND 0.300981f
C948 VPWR _098_ 0.404837f
C949 _253_/a_79_21# _143_ 0.058642f
C950 net19 net1 0.225906f
C951 _253_/a_79_21# _141_ 0.072441f
C952 VPWR net12 0.029883f
C953 VGND _000_ 0.044426f
C954 clkbuf_2_0__f_clk/a_110_47# counter\[9\] 0.022427f
C955 _060_ _077_ 0.065631f
C956 _011_ r2r_out[0] 0.048821f
C957 hold5/a_391_47# counter\[0\] 0.061571f
C958 divider\[1\] net6 0.024332f
C959 divider\[2\] _034_ 0.033509f
C960 VPWR clknet_2_2__leaf_clk 2.385854f
C961 VGND _028_ 0.054821f
C962 VGND _207_/a_35_297# 0.024977f
C963 _107_ hold2/a_285_47# 0.064146f
C964 VGND _262_/a_215_53# -0.016219f
C965 _184_/a_27_47# _092_ 0.015191f
C966 net8 _158_ 0.092911f
C967 _060_ _163_/a_27_47# 0.018167f
C968 _008_ _158_ 0.142056f
C969 VPWR _325_/a_891_413# 0.019937f
C970 VGND hold2/a_391_47# -0.014687f
C971 VPWR hold2/a_285_47# 0.041442f
C972 _072_ _057_ 0.020614f
C973 _148_ _272_/a_215_297# 0.039755f
C974 VPWR _298_/a_253_47# 0.015682f
C975 VGND _329_/a_27_47# -0.022916f
C976 counter\[14\] net9 0.136213f
C977 _355_/a_891_413# VPWR 0.034771f
C978 input8/a_27_47# net9 0.026421f
C979 _330_/a_27_47# net9 0.034245f
C980 _342_/a_1059_315# clknet_2_1__leaf_clk 0.068959f
C981 _325_/a_1059_315# net8 0.078537f
C982 counter\[13\] net9 0.102927f
C983 counter\[4\] _117_ 0.299773f
C984 _336_/a_27_47# r2r_out[3] 0.012566f
C985 _053_ _338_/a_193_47# 0.044881f
C986 _094_ _238_/a_227_47# 0.059602f
C987 _355_/a_466_413# _031_ 0.024948f
C988 VPWR _170_/a_299_297# 0.055065f
C989 _053_ _083_ 0.223489f
C990 _066_ _301_/a_27_47# 0.029451f
C991 counter\[0\] _097_ 0.232546f
C992 VPWR _151_ 0.520282f
C993 _219_/a_77_199# _117_ 0.020598f
C994 _060_ net4 0.091814f
C995 _176_/a_68_297# _085_ 0.024772f
C996 _104_ _020_ 0.226537f
C997 _144_ counter\[8\] 0.01577f
C998 clkbuf_2_0__f_clk/a_110_47# counter\[7\] 0.078611f
C999 VGND _285_/a_285_297# 0.020572f
C1000 counter\[9\] _133_ 0.032834f
C1001 _057_ _138_ 0.188589f
C1002 _066_ _313_/a_27_47# 0.07307f
C1003 _144_ _141_ 0.050032f
C1004 _090_ _088_ 0.07156f
C1005 r2r_out[7] _340_/a_27_47# 0.014593f
C1006 _187_/a_297_47# _349_/a_27_47# 0.010749f
C1007 _142_ _065_ 0.160989f
C1008 counter\[1\] hold5/a_391_47# 0.028713f
C1009 _149_ _262_/a_109_93# 0.013563f
C1010 _094_ _229_/a_77_199# 0.05795f
C1011 net10 _258_/a_27_47# 0.080065f
C1012 counter\[14\] clknet_2_2__leaf_clk 0.457401f
C1013 _117_ _118_ 0.114512f
C1014 _330_/a_27_47# clknet_2_2__leaf_clk 0.020368f
C1015 counter\[13\] clknet_2_2__leaf_clk 0.03559f
C1016 VGND _159_ 1.328217f
C1017 _094_ _127_ 0.013468f
C1018 _325_/a_1059_315# net6 0.042035f
C1019 _285_/a_285_297# counter\[15\] 0.010514f
C1020 VGND _296_/a_27_53# 0.047657f
C1021 _148_ net8 0.984413f
C1022 _060_ _341_/a_27_47# 0.098154f
C1023 divider\[3\] _159_ 0.010192f
C1024 _072_ _013_ 0.036424f
C1025 net7 _269_/a_27_413# 0.016025f
C1026 _051_ _078_ 0.343841f
C1027 _148_ _008_ 0.065514f
C1028 _168_/a_76_199# _077_ 0.044018f
C1029 _267_/a_215_297# net5 0.018347f
C1030 _267_/a_298_297# _004_ 0.027908f
C1031 _136_ _244_/a_59_75# 0.017767f
C1032 counter\[7\] _133_ 0.205754f
C1033 _081_ _086_ 0.181621f
C1034 _339_/a_1062_300# clk 0.02184f
C1035 VGND _085_ 0.02768f
C1036 counter\[1\] _097_ 0.147741f
C1037 VGND _338_/a_475_413# 0.013544f
C1038 _328_/a_193_47# rst 0.033275f
C1039 _003_ clknet_2_3__leaf_clk 0.084356f
C1040 counter\[15\] _159_ 0.074374f
C1041 _062_ _063_ 0.158066f
C1042 _296_/a_27_53# counter\[15\] 0.081041f
C1043 _136_ net4 0.094145f
C1044 _133_ _046_ 0.014052f
C1045 net5 _268_/a_109_93# 0.012202f
C1046 clknet_2_0__leaf_clk _350_/a_381_47# 0.048522f
C1047 net5 _077_ 0.036f
C1048 VPWR _330_/a_1059_315# 0.033628f
C1049 r2r_out[1] VPWR 3.448886f
C1050 _351_/a_634_159# counter\[10\] 0.038143f
C1051 VPWR _139_ 0.025143f
C1052 _094_ net18 0.054697f
C1053 _167_/a_27_47# _048_ 0.055349f
C1054 _065_ _099_ 0.025351f
C1055 VGND _208_/a_489_47# 0.035397f
C1056 _066_ hold2/a_391_47# 0.056193f
C1057 VGND _335_/a_27_47# 0.069929f
C1058 _148_ net6 0.230392f
C1059 _149_ _004_ 0.233809f
C1060 VGND _283_/a_78_199# 0.022108f
C1061 _338_/a_891_413# r2r_out[5] 0.045479f
C1062 _060_ _169_/a_51_297# 0.126645f
C1063 clknet_2_0__leaf_clk _127_ 0.016455f
C1064 _322_/a_27_47# r2r_out[3] 0.079542f
C1065 VGND _317_/a_113_297# 0.019054f
C1066 _355_/a_381_47# _066_ 0.016461f
C1067 _122_ _121_ 0.03464f
C1068 _104_ _344_/a_634_159# 0.040727f
C1069 _020_ _344_/a_27_47# 0.07982f
C1070 VPWR _344_/a_466_413# 0.010693f
C1071 VGND _344_/a_1059_315# 0.01561f
C1072 hold6/a_391_47# _078_ 0.03077f
C1073 hold6/a_285_47# _118_ 0.015561f
C1074 _296_/a_219_297# counter\[14\] 0.026118f
C1075 _263_/a_27_413# clknet_2_3__leaf_clk 0.027342f
C1076 net4 net1 0.037954f
C1077 counter\[10\] counter\[8\] 0.028653f
C1078 VGND _349_/a_1059_315# -0.012628f
C1079 VGND _328_/a_634_159# 0.032367f
C1080 VPWR _328_/a_193_47# 0.015776f
C1081 _039_ _048_ 0.090972f
C1082 net4 net5 0.396065f
C1083 _286_/a_219_297# _039_ 0.022359f
C1084 _006_ net8 0.059995f
C1085 counter\[15\] _283_/a_78_199# 0.074949f
C1086 VPWR net15 0.149193f
C1087 _060_ r2r_out[4] 0.16145f
C1088 r2r_out[3] _072_ 0.07894f
C1089 _105_ _108_ 0.157912f
C1090 _289_/a_489_413# _155_ 0.02174f
C1091 VGND input3/a_27_47# 0.035875f
C1092 _163_/a_109_297# _073_ 0.010099f
C1093 net8 _328_/a_27_47# 0.440469f
C1094 _348_/a_466_413# _024_ 0.038894f
C1095 _154_ _005_ 0.060361f
C1096 _353_/a_27_47# _078_ 0.440373f
C1097 _149_ data[1] 0.046132f
C1098 divider\[3\] _266_/a_109_93# 0.011347f
C1099 _357__12/LO VGND 0.071433f
C1100 _355_/a_466_413# clk 0.010238f
C1101 _053_ _054_ 0.178605f
C1102 VGND _329_/a_634_159# -0.014316f
C1103 r2r_out[3] _011_ 0.027091f
C1104 clkbuf_2_0__f_clk/a_110_47# VPWR 0.176906f
C1105 hold5/a_49_47# _098_ 0.043757f
C1106 _085_ _087_ 0.302884f
C1107 data[5] VGND 0.138754f
C1108 divider\[5\] _046_ 0.101237f
C1109 _326_/a_1059_315# clknet_2_3__leaf_clk 0.042429f
C1110 VPWR _297_/a_79_21# 0.051703f
C1111 VPWR _345_/a_634_159# 0.025541f
C1112 _148_ _280_/a_27_413# 0.010337f
C1113 _053_ _225_/a_75_212# 0.072307f
C1114 _336_/a_27_47# VPWR 0.132183f
C1115 _336_/a_193_47# VGND -0.220206f
C1116 _298_/a_103_199# _050_ 0.034919f
C1117 _330_/a_193_47# _006_ 0.220091f
C1118 hold8/a_285_47# _078_ 0.026197f
C1119 VGND input7/a_27_47# 0.045711f
C1120 _348_/a_27_47# _350_/a_1059_315# 0.010996f
C1121 _149_ net3 2.046946f
C1122 net19 _078_ 0.026641f
C1123 net6 _328_/a_27_47# 0.070264f
C1124 _104_ _200_/a_77_199# 0.010553f
C1125 net7 rst 2.757994f
C1126 divider\[1\] _263_/a_215_297# 0.029913f
C1127 VGND _079_ 0.072941f
C1128 _036_ divider\[2\] 0.109625f
C1129 counter\[2\] _098_ 0.048235f
C1130 _207_/a_285_297# counter\[4\] 0.062504f
C1131 _137_ _138_ 0.078266f
C1132 _167_/a_27_47# net9 0.04304f
C1133 _073_ _065_ 0.025284f
C1134 net7 _259_/a_27_47# 0.033551f
C1135 VGND _021_ 0.238491f
C1136 VPWR clknet_2_1__leaf_clk 1.840151f
C1137 VPWR _337_/a_27_47# 0.081077f
C1138 VGND _337_/a_193_47# -0.185768f
C1139 r2r_out[1] _333_/a_891_413# 0.042932f
C1140 VPWR _133_ 1.226605f
C1141 _094_ _205_/a_215_53# 0.051547f
C1142 VPWR _192_/a_27_47# 0.016639f
C1143 _094_ _344_/a_193_47# 0.051125f
C1144 _057_ _338_/a_475_413# 0.015268f
C1145 _157_ VGND 0.228254f
C1146 _082_ net9 0.039472f
C1147 _333_/a_27_47# _333_/a_475_413# -0.015098f
C1148 net9 _255_/a_80_21# 0.05644f
C1149 _054_ _303_/a_113_297# 0.023125f
C1150 net8 _054_ 0.199454f
C1151 _015_ clknet_2_3__leaf_clk 0.070111f
C1152 VGND _189_/a_47_47# 0.0364f
C1153 _053_ clknet_2_3__leaf_clk 0.370766f
C1154 _039_ net9 0.099063f
C1155 _065_ _344_/a_891_413# 0.036618f
C1156 VGND _086_ 0.108313f
C1157 VPWR net7 0.588971f
C1158 _125_ counter\[8\] 0.217568f
C1159 VPWR r2r_out[6] 1.239582f
C1160 _149_ counter\[5\] 0.052158f
C1161 _078_ counter\[11\] 0.586294f
C1162 _057_ _335_/a_27_47# 0.031988f
C1163 _274_/a_298_297# _148_ 0.014239f
C1164 _265_/a_27_413# _148_ 0.058973f
C1165 _058_ _056_ 0.493265f
C1166 _051_ counter\[11\] 0.079755f
C1167 clknet_0_clk net4 0.495026f
C1168 _223_/a_93_21# _054_ 0.070709f
C1169 VGND _115_ 0.25614f
C1170 _053_ _164_/a_79_21# 0.020812f
C1171 VGND _096_ 0.498083f
C1172 _351_/a_193_47# VPWR 0.014752f
C1173 _351_/a_634_159# VGND 0.026228f
C1174 _007_ rst 0.322462f
C1175 _292_/a_85_193# _042_ 0.010805f
C1176 _053_ net21 0.016494f
C1177 _326_/a_1059_315# net2 0.082362f
C1178 _135_ counter\[12\] 0.32846f
C1179 VGND _055_ 0.110306f
C1180 _047_ _051_ 0.245991f
C1181 _078_ _168_/a_505_21# 0.064325f
C1182 _057_ _349_/a_1059_315# 0.076157f
C1183 clknet_2_0__leaf_clk _344_/a_193_47# 0.010618f
C1184 _112_ _115_ 0.616098f
C1185 VGND _331_/a_1059_315# 0.045365f
C1186 _101_ _217_/a_27_47# 0.012969f
C1187 counter\[13\] _133_ 0.202094f
C1188 _224_/a_59_75# _057_ 0.041785f
C1189 _149_ divider\[2\] 0.031709f
C1190 _322_/a_27_47# VPWR 0.013664f
C1191 _356_/a_27_47# net1 0.032914f
C1192 _346_/a_27_47# VGND 0.064467f
C1193 VGND _174_/a_79_21# 0.04142f
C1194 _348_/a_27_47# VPWR -0.223862f
C1195 _348_/a_193_47# VGND -0.071802f
C1196 net6 _054_ 0.041092f
C1197 _039_ clknet_2_2__leaf_clk 0.19553f
C1198 _040_ divider\[5\] 0.087597f
C1199 _094_ clknet_2_0__leaf_clk 1.42759f
C1200 _053_ _067_ 0.296656f
C1201 _060_ _056_ 0.036689f
C1202 VGND counter\[8\] 0.998034f
C1203 net8 _331_/a_634_159# 0.018622f
C1204 counter\[12\] _054_ 0.135282f
C1205 _340_/a_193_47# _016_ 0.061544f
C1206 _263_/a_27_413# _151_ 0.010072f
C1207 _264_/a_215_53# net10 0.042243f
C1208 _286_/a_27_53# VPWR 0.013588f
C1209 VGND _143_ 0.081149f
C1210 divider\[4\] net10 0.809765f
C1211 _149_ input4/a_27_47# 0.027963f
C1212 VGND _141_ 0.704197f
C1213 _063_ _341_/a_891_413# 0.021861f
C1214 _084_ _178_/a_75_199# 0.095792f
C1215 VGND _154_ 0.046588f
C1216 VPWR divider\[5\] 0.370525f
C1217 _078_ _077_ 0.045936f
C1218 r2r_out[6] _181_/a_93_21# 0.012269f
C1219 _066_ _079_ 0.111879f
C1220 _174_/a_215_47# r2r_out[5] 0.03027f
C1221 _052_ _115_ 0.51889f
C1222 VPWR _012_ 0.161028f
C1223 VPWR _007_ 0.153422f
C1224 divider\[1\] _001_ 0.115274f
C1225 _005_ _329_/a_193_47# 0.068196f
C1226 VPWR _155_ 0.577289f
C1227 _072_ VPWR 0.546773f
C1228 VPWR _243_/a_250_297# 0.021742f
C1229 _149_ _342_/a_27_47# 0.010123f
C1230 _066_ _021_ 0.088691f
C1231 _148_ _263_/a_215_297# 0.043997f
C1232 _072_ _171_/a_27_47# 0.011837f
C1233 _200_/a_227_47# hold4/a_49_47# 0.029857f
C1234 _148_ _269_/a_298_297# 0.038875f
C1235 r2r_out[1] counter\[2\] 0.015844f
C1236 divider\[6\] _331_/a_381_47# 0.028183f
C1237 _152_ net4 0.014394f
C1238 net8 clknet_2_3__leaf_clk 0.022766f
C1239 counter\[15\] counter\[8\] 0.021848f
C1240 _336_/a_193_47# _057_ 0.032677f
C1241 _246_/a_113_297# _045_ 0.011805f
C1242 _065_ _100_ 0.076425f
C1243 counter\[9\] _159_ 0.100765f
C1244 _053_ net2 0.034992f
C1245 _060_ _017_ 0.159045f
C1246 VPWR _011_ 0.153891f
C1247 _053_ net9 0.493554f
C1248 _353_/a_381_47# _029_ 0.022557f
C1249 _347_/a_1059_315# counter\[6\] 0.024899f
C1250 _294_/a_78_199# divider\[5\] 0.016259f
C1251 _057_ _079_ 0.070472f
C1252 net4 _078_ 0.023982f
C1253 VPWR _138_ 0.088396f
C1254 _052_ counter\[8\] 0.048154f
C1255 _149_ _348_/a_634_159# 0.019383f
C1256 divider\[0\] _279_/a_207_413# 0.014538f
C1257 _054_ _341_/a_1059_315# 0.010374f
C1258 _027_ _149_ 0.162184f
C1259 _048_ _049_ 0.01425f
C1260 _057_ _337_/a_193_47# 0.361296f
C1261 _089_ rst 0.067339f
C1262 _286_/a_219_297# _049_ 0.01548f
C1263 _094_ _097_ 0.073555f
C1264 VGND _340_/a_27_47# 0.023286f
C1265 _286_/a_27_53# counter\[14\] 0.014947f
C1266 _066_ _096_ 0.020217f
C1267 counter\[13\] divider\[5\] 0.051123f
C1268 net6 clknet_2_3__leaf_clk 0.038675f
C1269 _089_ _259_/a_27_47# 0.010238f
C1270 _169_/a_51_297# _076_ 0.04902f
C1271 VPWR _301_/a_27_47# 0.033679f
C1272 _052_ hold6/a_49_47# 0.01186f
C1273 VGND _142_ 0.257003f
C1274 _342_/a_27_47# _065_ 0.040889f
C1275 clknet_0_clk counter\[4\] 0.010248f
C1276 _078_ _341_/a_27_47# 0.015161f
C1277 _055_ r2r_out[0] 0.21422f
C1278 counter\[9\] _283_/a_78_199# 0.027362f
C1279 counter\[13\] _155_ 0.02223f
C1280 counter\[12\] _243_/a_93_21# 0.054196f
C1281 _160_ VPWR 0.094842f
C1282 VPWR _313_/a_27_47# 0.177746f
C1283 rst _000_ 0.048606f
C1284 _159_ _046_ 0.012273f
C1285 net22 _060_ 0.016879f
C1286 _353_/a_193_47# net1 0.039437f
C1287 _345_/a_891_413# counter\[4\] 0.030396f
C1288 r2r_out[1] _318_/a_27_47# 0.07306f
C1289 _356_/a_27_47# _032_ 0.064592f
C1290 _066_ counter\[8\] 0.526263f
C1291 _135_ _059_ 0.132607f
C1292 _262_/a_215_53# rst 0.047547f
C1293 _066_ _143_ 0.227512f
C1294 _287_/a_215_53# clknet_2_2__leaf_clk 0.023109f
C1295 _076_ r2r_out[4] 0.066024f
C1296 _066_ _141_ 0.073308f
C1297 _089_ VPWR 0.045946f
C1298 _352_/a_381_47# counter\[11\] 0.016472f
C1299 _236_/a_27_47# counter\[8\] 0.030694f
C1300 _346_/a_27_47# _022_ 0.027306f
C1301 _346_/a_193_47# _065_ 0.042399f
C1302 net2 net8 0.018862f
C1303 net8 net9 0.048697f
C1304 _013_ _337_/a_193_47# 0.069738f
C1305 VPWR _352_/a_466_413# 0.014699f
C1306 VGND _352_/a_1059_315# 0.058905f
C1307 _197_/a_27_47# hold4/a_391_47# 0.010423f
C1308 _149_ _350_/a_27_47# 0.033396f
C1309 _008_ _275_/a_215_53# 0.011774f
C1310 _150_ net1 0.03618f
C1311 _059_ _054_ 0.404997f
C1312 VPWR ext_data 0.229312f
C1313 _057_ _174_/a_79_21# 0.031754f
C1314 clknet_0_clk _045_ 0.022319f
C1315 _148_ _001_ 0.032697f
C1316 divider\[0\] VPWR 0.637067f
C1317 VGND _099_ 0.290034f
C1318 _057_ counter\[8\] 0.392309f
C1319 _042_ _041_ 0.374079f
C1320 counter\[2\] clknet_2_1__leaf_clk 0.076035f
C1321 VPWR _000_ 0.243631f
C1322 _274_/a_27_413# _157_ 0.051499f
C1323 _057_ _143_ 0.199099f
C1324 data[4] net10 0.03489f
C1325 _057_ _141_ 0.180779f
C1326 clkbuf_0_clk/a_110_47# counter\[8\] 0.019273f
C1327 _221_/a_68_297# counter\[8\] 0.067021f
C1328 VPWR _028_ 0.062621f
C1329 _060_ _178_/a_75_199# 0.048292f
C1330 VPWR _207_/a_35_297# 0.093029f
C1331 _107_ hold2/a_391_47# 0.056122f
C1332 _274_/a_215_297# net7 0.044773f
C1333 VPWR _260_/a_109_93# 0.010558f
C1334 VGND _262_/a_109_93# -0.011543f
C1335 _149_ _060_ 0.052055f
C1336 _148_ net10 0.161688f
C1337 net14 hold2/a_391_47# 0.02476f
C1338 _223_/a_93_21# _121_ 0.02306f
C1339 net6 net2 0.025537f
C1340 net8 clknet_2_2__leaf_clk 0.179344f
C1341 divider\[2\] data[3] 0.126734f
C1342 net6 net9 1.041093f
C1343 _094_ _131_ 0.041801f
C1344 _008_ clknet_2_2__leaf_clk 0.017307f
C1345 _089_ _181_/a_93_21# 0.0441f
C1346 VPWR _329_/a_27_47# -0.208981f
C1347 VGND _329_/a_193_47# -0.13731f
C1348 _330_/a_193_47# net9 0.035331f
C1349 _342_/a_891_413# clknet_2_1__leaf_clk 0.052862f
C1350 _325_/a_891_413# net8 0.078768f
C1351 hold4/a_49_47# counter\[3\] 0.023473f
C1352 _333_/a_193_47# _056_ 0.011462f
C1353 _333_/a_27_47# _009_ 0.102006f
C1354 _071_ r2r_out[2] 1.040702f
C1355 _190_/a_76_199# _095_ 0.031512f
C1356 _311_/a_27_297# r2r_out[0] 0.010353f
C1357 input4/a_27_47# data[3] 0.021651f
C1358 _003_ net7 0.026777f
C1359 _071_ _065_ 0.022844f
C1360 r2r_out[1] _053_ 0.121289f
C1361 _124_ _132_ 0.035834f
C1362 VGND _308_/a_27_47# 0.052607f
C1363 r2r_out[7] _340_/a_193_47# 0.015407f
C1364 r2r_out[3] _337_/a_193_47# 0.010263f
C1365 _004_ VGND 0.121642f
C1366 data[7] net10 0.118972f
C1367 _070_ clk 0.179885f
C1368 net6 clknet_2_2__leaf_clk 0.180586f
C1369 _060_ r2r_out[2] 0.030376f
C1370 _342_/a_193_47# _342_/a_634_159# -0.016573f
C1371 _078_ _118_ 0.206749f
C1372 _330_/a_193_47# clknet_2_2__leaf_clk 0.010899f
C1373 _243_/a_93_21# _059_ 0.047395f
C1374 _325_/a_891_413# net6 0.040501f
C1375 VPWR _159_ 0.428239f
C1376 _342_/a_1059_315# _096_ 0.023802f
C1377 _214_/a_113_297# VPWR 0.034018f
C1378 _060_ _065_ 0.044381f
C1379 _060_ _341_/a_193_47# 0.474799f
C1380 net7 _269_/a_215_297# 0.066547f
C1381 _045_ _078_ 0.564172f
C1382 _163_/a_27_47# _074_ 0.017077f
C1383 divider\[1\] _280_/a_207_413# 0.01287f
C1384 _051_ _045_ 0.202807f
C1385 _101_ _019_ 0.021118f
C1386 r2r_out[5] _077_ 0.348944f
C1387 _060_ r2r_out[7] 0.011813f
C1388 _101_ counter\[4\] 0.749119f
C1389 _078_ _129_ 0.012759f
C1390 _149_ _267_/a_27_413# 0.044686f
C1391 _146_ net20 0.010519f
C1392 _081_ _084_ 0.108963f
C1393 clknet_0_clk _035_ 0.020281f
C1394 VGND _227_/a_59_75# -0.016621f
C1395 VPWR _085_ 0.046875f
C1396 VGND _338_/a_1062_300# 0.065553f
C1397 _061_ _064_ 0.051336f
C1398 _328_/a_634_159# rst 0.01831f
C1399 _046_ clkbuf_2_2__f_clk/a_110_47# 0.025914f
C1400 VGND data[1] 0.036556f
C1401 net4 _074_ 0.08671f
C1402 VPWR _330_/a_891_413# 0.043846f
C1403 _351_/a_466_413# counter\[10\] 0.033957f
C1404 _149_ net1 1.471234f
C1405 _094_ hold2/a_49_47# 0.034305f
C1406 _267_/a_215_297# net4 0.038017f
C1407 VGND _335_/a_193_47# 0.034093f
C1408 VPWR _335_/a_27_47# 0.121391f
C1409 _149_ net5 0.044019f
C1410 counter\[9\] counter\[8\] 0.76518f
C1411 _338_/a_381_47# r2r_out[5] 0.013934f
C1412 VPWR _317_/a_113_297# 0.035925f
C1413 counter\[9\] _141_ 0.024421f
C1414 counter\[7\] _115_ 0.154535f
C1415 _053_ _336_/a_27_47# 0.339167f
C1416 _104_ _344_/a_466_413# 0.034099f
C1417 _269_/a_27_413# _154_ 0.026164f
C1418 VPWR _344_/a_1059_315# 0.043323f
C1419 _187_/a_79_21# clknet_2_1__leaf_clk 0.068498f
C1420 divider\[1\] _033_ 0.151663f
C1421 _214_/a_113_297# _114_ 0.055778f
C1422 hold6/a_391_47# _118_ 0.037571f
C1423 VGND _256_/a_81_21# 0.039292f
C1424 counter\[14\] _159_ 0.024664f
C1425 _343_/a_27_47# _019_ 0.055379f
C1426 counter\[13\] _159_ 1.142187f
C1427 _263_/a_215_297# clknet_2_3__leaf_clk 0.088368f
C1428 _094_ _109_ 0.140012f
C1429 _027_ counter\[10\] 0.266294f
C1430 VGND net3 1.191278f
C1431 _094_ _020_ 0.032792f
C1432 net16 _100_ 0.245063f
C1433 VPWR _328_/a_634_159# 0.013219f
C1434 VGND _328_/a_466_413# 0.025776f
C1435 _105_ _094_ 0.042748f
C1436 clknet_2_1__leaf_clk _103_ 0.024103f
C1437 _062_ _054_ 0.509312f
C1438 _238_/a_77_199# _078_ 0.044623f
C1439 _338_/a_27_47# _338_/a_193_47# -0.157669f
C1440 _053_ clknet_2_1__leaf_clk 0.245067f
C1441 VPWR input3/a_27_47# 0.047859f
C1442 _163_/a_193_297# _073_ 0.061668f
C1443 _163_/a_27_47# net4 0.115212f
C1444 _141_ _248_/a_77_199# 0.047276f
C1445 _053_ _337_/a_27_47# 0.04902f
C1446 _083_ _338_/a_27_47# 0.031196f
C1447 _238_/a_77_199# _051_ 0.012427f
C1448 net8 _328_/a_193_47# 0.067734f
C1449 _348_/a_1059_315# _024_ 0.078197f
C1450 _192_/a_27_47# _103_ 0.014178f
C1451 _213_/a_215_53# _212_/a_80_21# 0.011431f
C1452 _353_/a_193_47# _078_ 0.05026f
C1453 r2r_out[3] _164_/a_215_47# 0.034051f
C1454 _137_ counter\[8\] 0.028359f
C1455 _195_/a_227_47# _100_ 0.03142f
C1456 _101_ _200_/a_227_47# 0.010856f
C1457 _357__12/LO VPWR 0.13209f
C1458 hold9/a_391_47# net21 0.016651f
C1459 counter\[15\] net3 0.032153f
C1460 VPWR _329_/a_634_159# 0.01645f
C1461 _143_ _147_ 0.158435f
C1462 _141_ _147_ 0.027955f
C1463 hold5/a_285_47# _098_ 0.059802f
C1464 _035_ _078_ 0.07256f
C1465 _059_ _121_ 0.019142f
C1466 _057_ _308_/a_27_47# 0.019347f
C1467 _073_ _075_ 0.246233f
C1468 _141_ _046_ 0.218338f
C1469 counter\[4\] _217_/a_27_47# 0.047377f
C1470 VGND _120_ 0.35194f
C1471 data[5] VPWR 0.419928f
C1472 _015_ r2r_out[6] 0.110047f
C1473 _326_/a_891_413# clknet_2_3__leaf_clk 0.03857f
C1474 _053_ r2r_out[6] 0.100252f
C1475 VPWR _345_/a_466_413# 0.028701f
C1476 VGND _237_/a_27_47# 0.01976f
C1477 counter\[7\] hold6/a_49_47# 0.048557f
C1478 clknet_2_0__leaf_clk _020_ 0.09221f
C1479 VGND counter\[5\] 1.053721f
C1480 _336_/a_193_47# VPWR 0.037833f
C1481 hold8/a_391_47# _078_ 0.016217f
C1482 VGND _281_/a_27_47# 0.043137f
C1483 VPWR input7/a_27_47# 0.070233f
C1484 _066_ _073_ 0.12261f
C1485 _144_ _136_ 0.051661f
C1486 _017_ _078_ 0.03297f
C1487 rst _185_/a_113_297# 0.048097f
C1488 net6 _328_/a_193_47# 0.374925f
C1489 _265_/a_27_413# clknet_2_2__leaf_clk 0.014618f
C1490 divider\[1\] _263_/a_298_297# 0.039009f
C1491 _094_ _140_ 0.026491f
C1492 VPWR _079_ 0.245843f
C1493 _040_ clkbuf_2_2__f_clk/a_110_47# 0.010055f
C1494 counter\[0\] _098_ 0.444682f
C1495 _107_ _021_ 0.03411f
C1496 _112_ _237_/a_27_47# 0.043652f
C1497 VGND _100_ 0.414555f
C1498 _125_ _117_ 0.028498f
C1499 _344_/a_27_47# _344_/a_466_413# -0.013083f
C1500 _344_/a_193_47# _344_/a_634_159# -0.016573f
C1501 r2r_out[1] _068_ 0.051803f
C1502 VPWR _021_ 0.265207f
C1503 VPWR _337_/a_193_47# 0.060558f
C1504 net2 _263_/a_215_297# 0.012678f
C1505 r2r_out[1] _333_/a_381_47# 0.014456f
C1506 VPWR clkbuf_2_2__f_clk/a_110_47# 0.164143f
C1507 _094_ _205_/a_109_93# 0.018979f
C1508 r2r_out[1] _341_/a_1059_315# 0.027665f
C1509 _101_ _113_ 0.235815f
C1510 VGND divider\[2\] 0.949219f
C1511 counter\[15\] _281_/a_27_47# 0.037512f
C1512 r2r_out[7] _088_ 0.011706f
C1513 r2r_out[4] r2r_out[5] 0.27502f
C1514 _079_ _080_ 0.076829f
C1515 _094_ _344_/a_634_159# 0.016202f
C1516 _081_ _060_ 0.248956f
C1517 _057_ _338_/a_1062_300# 0.013791f
C1518 _149_ clknet_0_clk 0.055212f
C1519 _066_ _256_/a_81_21# 0.033285f
C1520 _057_ _073_ 0.028316f
C1521 VGND n_rst 0.060671f
C1522 _157_ VPWR 0.279697f
C1523 divider\[6\] data[6] 0.228236f
C1524 _071_ _069_ 0.016223f
C1525 _066_ net3 0.384107f
C1526 _001_ clknet_2_3__leaf_clk 0.139762f
C1527 _333_/a_193_47# _333_/a_475_413# -0.022086f
C1528 VGND input4/a_27_47# 0.041948f
C1529 _052_ _237_/a_27_47# 0.013054f
C1530 data[0] VGND 0.058096f
C1531 VPWR _189_/a_47_47# 0.042486f
C1532 _149_ _234_/a_113_297# 0.012686f
C1533 _331_/a_27_47# clknet_2_2__leaf_clk 0.018652f
C1534 _053_ _012_ 0.139176f
C1535 _065_ _344_/a_381_47# 0.019416f
C1536 VPWR _086_ 0.102801f
C1537 _124_ _121_ 0.124208f
C1538 VGND _084_ 0.62237f
C1539 _081_ _183_/a_59_75# 0.012183f
C1540 _069_ _319_/a_29_53# 0.010925f
C1541 _149_ hold1/a_49_47# 0.04734f
C1542 _053_ _072_ 0.054559f
C1543 _057_ _335_/a_193_47# 0.033834f
C1544 _334_/a_475_413# clknet_2_1__leaf_clk 0.02067f
C1545 _264_/a_215_53# _327_/a_1059_315# 0.011703f
C1546 _078_ counter\[3\] 0.014258f
C1547 r2r_out[4] _077_ 0.060567f
C1548 VGND _123_ 0.112054f
C1549 _265_/a_215_297# _148_ 0.034534f
C1550 counter\[15\] divider\[2\] 0.08228f
C1551 _058_ _009_ 0.02823f
C1552 _045_ counter\[11\] 0.050396f
C1553 VGND _342_/a_27_47# 0.011634f
C1554 _154_ rst 0.226313f
C1555 _223_/a_250_297# _054_ 0.024136f
C1556 VGND _117_ 1.245088f
C1557 _060_ _093_ 0.071585f
C1558 VPWR _115_ 0.352861f
C1559 net7 net8 0.023663f
C1560 _057_ _333_/a_27_47# 0.238139f
C1561 VPWR _096_ 0.470503f
C1562 r2r_out[6] net8 0.021389f
C1563 _351_/a_466_413# VGND 0.03451f
C1564 _351_/a_634_159# VPWR 0.010112f
C1565 counter\[1\] _098_ 0.052585f
C1566 _057_ _256_/a_81_21# 0.126722f
C1567 _053_ _011_ 0.07457f
C1568 _326_/a_891_413# net2 0.042747f
C1569 _078_ clkbuf_2_1__f_clk/a_110_47# 0.134725f
C1570 counter\[11\] _129_ 0.014041f
C1571 _060_ _069_ 0.068116f
C1572 _057_ net3 0.015794f
C1573 _057_ _349_/a_891_413# 0.039146f
C1574 _291_/a_27_47# divider\[5\] 0.04513f
C1575 hold10/a_285_47# _340_/a_634_183# 0.010905f
C1576 _112_ _117_ 0.659763f
C1577 _325_/a_466_413# clknet_2_3__leaf_clk 0.014643f
C1578 _010_ clknet_2_1__leaf_clk 0.231668f
C1579 _149_ net13 0.024087f
C1580 counter\[14\] clkbuf_2_2__f_clk/a_110_47# 0.274005f
C1581 VGND _331_/a_891_413# 0.044712f
C1582 VPWR _331_/a_1059_315# 0.01149f
C1583 counter\[13\] clkbuf_2_2__f_clk/a_110_47# 0.037955f
C1584 counter\[12\] _133_ 0.14742f
C1585 _224_/a_59_75# _122_ 0.035274f
C1586 _356_/a_193_47# net1 0.041242f
C1587 VPWR _174_/a_79_21# 0.085252f
C1588 _346_/a_27_47# VPWR 0.095997f
C1589 _346_/a_193_47# VGND -0.010809f
C1590 _348_/a_634_159# VGND 0.017456f
C1591 _348_/a_193_47# VPWR -0.023663f
C1592 _291_/a_27_47# _155_ 0.018159f
C1593 clknet_0_clk _041_ 0.031382f
C1594 _073_ _013_ 0.061148f
C1595 _066_ counter\[5\] 0.21562f
C1596 _027_ VGND 0.014115f
C1597 VPWR counter\[8\] 1.538669f
C1598 net8 _331_/a_466_413# 0.015908f
C1599 _350_/a_27_47# _026_ 0.032439f
C1600 counter\[6\] _212_/a_80_21# 0.032959f
C1601 _148_ _331_/a_193_47# 0.0108f
C1602 VPWR _143_ 0.719947f
C1603 VPWR _141_ 0.59329f
C1604 _094_ _200_/a_77_199# 0.109431f
C1605 VPWR _154_ 0.200293f
C1606 counter\[6\] _094_ 0.161706f
C1607 r2r_out[6] _181_/a_250_297# 0.014098f
C1608 net6 net7 0.055715f
C1609 _081_ _168_/a_76_199# 0.011563f
C1610 net6 r2r_out[6] 0.07786f
C1611 hold1/a_49_47# _065_ 0.021624f
C1612 _052_ _117_ 0.298022f
C1613 _101_ counter\[3\] 0.169195f
C1614 _078_ _178_/a_75_199# 0.021969f
C1615 _062_ net2 0.056647f
C1616 VGND _042_ 0.105919f
C1617 _349_/a_27_47# clknet_2_1__leaf_clk 0.021213f
C1618 _114_ _115_ 0.284248f
C1619 _149_ _078_ 0.237492f
C1620 _148_ _263_/a_298_297# 0.017686f
C1621 _057_ _120_ 0.067323f
C1622 _197_/a_27_47# net16 0.049134f
C1623 r2r_out[1] counter\[0\] 0.044331f
C1624 net15 _128_ 0.071126f
C1625 VPWR hold6/a_49_47# 0.027747f
C1626 net11 r2r_out[7] 0.012103f
C1627 _347_/a_381_47# clknet_2_0__leaf_clk 0.019083f
C1628 _076_ _065_ 0.017848f
C1629 _021_ _106_ 0.012844f
C1630 _336_/a_634_183# _057_ 0.019105f
C1631 _238_/a_77_199# counter\[11\] 0.087712f
C1632 _053_ _089_ 0.034882f
C1633 net17 _065_ 0.021646f
C1634 _072_ _173_/a_27_47# 0.013125f
C1635 _149_ _348_/a_466_413# 0.0138f
C1636 _005_ net5 0.0215f
C1637 _044_ divider\[4\] 0.171112f
C1638 _325_/a_1059_315# _261_/a_27_413# 0.010054f
C1639 net10 net9 1.543959f
C1640 VGND _058_ 0.013733f
C1641 _227_/a_59_75# counter\[9\] 0.03056f
C1642 _057_ _337_/a_634_183# 0.036791f
C1643 _229_/a_227_47# _126_ 0.100786f
C1644 _071_ VGND 0.094059f
C1645 _286_/a_27_53# _049_ 0.094224f
C1646 counter\[14\] counter\[8\] 0.309267f
C1647 VPWR _340_/a_27_47# 0.121223f
C1648 _275_/a_215_53# net10 0.027108f
C1649 VGND _350_/a_27_47# 0.076646f
C1650 counter\[14\] _143_ 0.02972f
C1651 _035_ counter\[11\] 0.16185f
C1652 _053_ _305_/a_27_47# 0.057003f
C1653 counter\[14\] _141_ 0.775887f
C1654 _148_ divider\[4\] 0.019657f
C1655 _338_/a_27_47# clknet_2_3__leaf_clk 0.019803f
C1656 counter\[13\] _141_ 0.162188f
C1657 VPWR _311_/a_27_297# 0.041437f
C1658 VGND _311_/a_109_297# 0.016684f
C1659 VGND _319_/a_29_53# 0.043498f
C1660 _169_/a_51_297# r2r_out[4] 0.012655f
C1661 _063_ _054_ 0.234255f
C1662 _072_ net6 0.011345f
C1663 _054_ clk 0.032928f
C1664 VPWR _142_ 1.100309f
C1665 _342_/a_193_47# _065_ 0.036149f
C1666 _081_ _088_ 0.031837f
C1667 _149_ _101_ 1.085865f
C1668 _065_ _078_ 0.012557f
C1669 _352_/a_27_47# clknet_2_2__leaf_clk 0.022372f
C1670 _149_ _024_ 0.068557f
C1671 counter\[12\] _243_/a_250_297# 0.023907f
C1672 _018_ _065_ 0.1926f
C1673 _065_ _051_ 0.03601f
C1674 _300_/a_27_47# VGND 0.046222f
C1675 _149_ _320_/a_80_21# 0.028196f
C1676 VGND hold8/a_49_47# 0.101136f
C1677 VGND _197_/a_27_47# 0.049976f
C1678 VGND _060_ 1.765908f
C1679 _065_ _061_ 0.077928f
C1680 _123_ _057_ 0.067084f
C1681 _356_/a_193_47# _032_ 0.057611f
C1682 _060_ _324_/a_68_297# 0.013456f
C1683 net10 clknet_2_2__leaf_clk 1.488459f
C1684 _148_ _261_/a_27_413# 0.026485f
C1685 _262_/a_109_93# rst 0.014322f
C1686 _148_ divider\[1\] 0.156185f
C1687 net13 hold1/a_391_47# 0.02476f
C1688 VPWR _195_/a_77_199# -0.021671f
C1689 _221_/a_68_297# _117_ 0.011559f
C1690 VPWR _229_/a_227_47# 0.02009f
C1691 clkbuf_2_3__f_clk/a_110_47# net3 0.029931f
C1692 _346_/a_193_47# _022_ 0.083484f
C1693 hold1/a_285_47# _219_/a_77_199# 0.013605f
C1694 VGND _183_/a_59_75# 0.032149f
C1695 counter\[12\] _138_ 0.030206f
C1696 _149_ _353_/a_27_47# 0.03822f
C1697 _059_ _133_ 0.137628f
C1698 _033_ _161_ 0.169718f
C1699 r2r_out[4] _337_/a_1062_300# 0.04735f
C1700 VGND _352_/a_891_413# 0.053043f
C1701 VPWR _352_/a_1059_315# 0.028134f
C1702 _351_/a_27_47# clknet_2_0__leaf_clk 0.227695f
C1703 _279_/a_27_413# net5 0.031879f
C1704 _321_/a_79_199# r2r_out[2] 0.024474f
C1705 hold8/a_49_47# counter\[15\] 0.035549f
C1706 _149_ _350_/a_193_47# 0.039754f
C1707 _060_ counter\[15\] 0.02904f
C1708 _002_ net3 0.031468f
C1709 VPWR _099_ 0.061577f
C1710 _122_ counter\[8\] 0.116863f
C1711 _253_/a_215_47# _141_ 0.036505f
C1712 counter\[0\] clknet_2_1__leaf_clk 0.148042f
C1713 _274_/a_215_297# _157_ 0.044126f
C1714 _101_ _065_ 0.194736f
C1715 _024_ _065_ 0.28514f
C1716 _300_/a_27_47# _052_ 0.03445f
C1717 counter\[13\] _142_ 0.142525f
C1718 divider\[0\] net8 0.040919f
C1719 _256_/a_81_21# _147_ 0.022696f
C1720 _192_/a_27_47# counter\[0\] 0.047789f
C1721 _265_/a_27_413# net7 0.016003f
C1722 _353_/a_891_413# _139_ 0.011429f
C1723 _149_ net19 0.104325f
C1724 _105_ hold2/a_49_47# 0.030825f
C1725 VGND _136_ 0.748591f
C1726 clk clknet_2_3__leaf_clk 0.101411f
C1727 counter\[9\] _281_/a_27_47# 0.0141f
C1728 r2r_out[1] _062_ 0.099562f
C1729 VPWR _329_/a_193_47# 0.010314f
C1730 _089_ net6 0.147879f
C1731 _071_ r2r_out[0] 0.062691f
C1732 _342_/a_381_47# clknet_2_1__leaf_clk 0.011331f
C1733 _325_/a_381_47# net8 0.0166f
C1734 _015_ _085_ 0.010761f
C1735 _148_ _325_/a_1059_315# 0.03192f
C1736 _053_ _338_/a_475_413# 0.018044f
C1737 _190_/a_206_369# _095_ 0.018155f
C1738 _355_/a_27_47# net1 0.037804f
C1739 _167_/a_27_47# clkbuf_2_2__f_clk/a_110_47# 0.020129f
C1740 _219_/a_77_199# _118_ 0.031357f
C1741 VPWR _308_/a_27_47# 0.012996f
C1742 hold4/a_285_47# clkbuf_2_1__f_clk/a_110_47# 0.010854f
C1743 _082_ _079_ 0.015319f
C1744 divider\[0\] net6 0.023492f
C1745 counter\[9\] divider\[2\] 0.071131f
C1746 _053_ _335_/a_27_47# 0.03842f
C1747 _343_/a_27_47# _065_ 0.017249f
C1748 VGND net1 2.176015f
C1749 counter\[1\] clknet_2_1__leaf_clk 0.129138f
C1750 _066_ _060_ 0.198374f
C1751 _065_ _354_/a_27_47# 0.048413f
C1752 VGND net5 3.03153f
C1753 _060_ r2r_out[0] 0.269513f
C1754 _004_ VPWR 0.432254f
C1755 counter\[7\] _237_/a_27_47# 0.117897f
C1756 hold10/a_49_47# r2r_out[7] 0.041157f
C1757 _067_ clk 0.123464f
C1758 _289_/a_489_413# divider\[2\] 0.023313f
C1759 _243_/a_250_297# _059_ 0.013984f
C1760 _325_/a_381_47# net6 0.020497f
C1761 _342_/a_891_413# _096_ 0.024645f
C1762 VGND _179_/a_79_21# 0.029742f
C1763 _060_ _341_/a_634_159# 0.041517f
C1764 _017_ _341_/a_27_47# 0.04768f
C1765 _258_/a_27_47# clknet_2_2__leaf_clk 0.076588f
C1766 net6 _329_/a_27_47# 0.016262f
C1767 divider\[6\] divider\[7\] 0.050602f
C1768 counter\[9\] _117_ 0.125371f
C1769 counter\[15\] net1 0.025435f
C1770 _090_ _065_ 0.012833f
C1771 _331_/a_27_47# _331_/a_466_413# -0.013083f
C1772 counter\[15\] net5 0.011089f
C1773 _149_ _267_/a_215_297# 0.075402f
C1774 _057_ _060_ 0.391538f
C1775 VPWR _227_/a_59_75# 0.017482f
C1776 rst net3 0.024638f
C1777 _090_ r2r_out[7] 0.076927f
C1778 VPWR _338_/a_1062_300# 0.072032f
C1779 VPWR _073_ 0.651361f
C1780 VGND _088_ 0.141838f
C1781 net2 clk 0.017469f
C1782 VPWR data[1] 0.246898f
C1783 counter\[10\] _078_ 0.076068f
C1784 clk net9 0.22012f
C1785 _351_/a_1059_315# counter\[10\] 0.047259f
C1786 counter\[10\] _051_ 0.03188f
C1787 VGND _156_ 0.130197f
C1788 _094_ hold2/a_285_47# 0.046383f
C1789 divider\[3\] _156_ 0.011793f
C1790 _331_/a_27_47# _007_ 0.074263f
C1791 _266_/a_215_53# net10 0.043892f
C1792 counter\[10\] _247_/a_27_47# 0.011996f
C1793 VGND _335_/a_634_183# 0.017109f
C1794 VPWR _335_/a_193_47# 0.032789f
C1795 _066_ _136_ 0.04125f
C1796 _105_ _205_/a_109_93# 0.011495f
C1797 _065_ counter\[11\] 0.096164f
C1798 _025_ _093_ 0.017418f
C1799 counter\[4\] _113_ 0.01057f
C1800 _065_ _190_/a_76_199# 0.025415f
C1801 VPWR _333_/a_27_47# -0.120547f
C1802 VGND _333_/a_193_47# -0.113847f
C1803 _024_ _119_ 0.03241f
C1804 counter\[7\] _117_ 0.068494f
C1805 _053_ _336_/a_193_47# 0.208649f
C1806 _104_ _344_/a_1059_315# 0.066941f
C1807 _269_/a_215_297# _154_ 0.029587f
C1808 VPWR _344_/a_891_413# 0.030278f
C1809 _278_/a_27_53# _034_ 0.032962f
C1810 VPWR _256_/a_81_21# 0.084455f
C1811 _343_/a_193_47# _019_ 0.051459f
C1812 counter\[12\] _159_ 0.415636f
C1813 divider\[2\] _327_/a_193_47# 0.106155f
C1814 divider\[6\] _273_/a_215_53# 0.035711f
C1815 _074_ _065_ 0.060677f
C1816 VPWR net3 1.249206f
C1817 clkbuf_2_0__f_clk/a_110_47# net18 0.027972f
C1818 _334_/a_1062_300# r2r_out[1] 0.029068f
C1819 _069_ _078_ 0.01173f
C1820 VPWR _328_/a_466_413# 0.012585f
C1821 _143_ _255_/a_80_21# 0.012142f
C1822 _141_ _255_/a_80_21# 0.010881f
C1823 divider\[3\] _328_/a_1059_315# 0.024009f
C1824 _060_ _013_ 0.087574f
C1825 _148_ _006_ 0.03346f
C1826 _136_ _057_ 0.584781f
C1827 _065_ r2r_out[5] 0.39218f
C1828 _087_ _179_/a_79_21# 0.078501f
C1829 _053_ _337_/a_193_47# 0.037576f
C1830 _066_ net1 0.071216f
C1831 _083_ _338_/a_193_47# 0.287371f
C1832 _065_ _095_ 0.173139f
C1833 net8 _328_/a_634_159# 0.017098f
C1834 _348_/a_891_413# _024_ 0.056589f
C1835 _149_ net4 0.104142f
C1836 _136_ clkbuf_0_clk/a_110_47# 0.035138f
C1837 _353_/a_634_159# _078_ 0.015872f
C1838 _054_ net20 0.18372f
C1839 VGND _032_ 0.259347f
C1840 VPWR _329_/a_466_413# 0.017339f
C1841 _094_ _216_/a_59_75# 0.015702f
C1842 clknet_0_clk VGND 2.314655f
C1843 hold5/a_49_47# _099_ 0.036459f
C1844 hold5/a_391_47# _098_ 0.056393f
C1845 _065_ _077_ 0.022174f
C1846 VGND _240_/a_68_297# 0.032491f
C1847 counter\[2\] _195_/a_77_199# 0.010093f
C1848 divider\[2\] rst 0.095016f
C1849 _053_ _185_/a_113_297# 0.064257f
C1850 _107_ _345_/a_1059_315# 0.011356f
C1851 _035_ _045_ 0.807475f
C1852 VPWR _120_ 0.033546f
C1853 counter\[5\] _107_ 0.198766f
C1854 _326_/a_381_47# clknet_2_3__leaf_clk 0.019078f
C1855 _163_/a_27_47# _065_ 0.020893f
C1856 VPWR _345_/a_1059_315# 0.020211f
C1857 _057_ net1 0.249252f
C1858 _167_/a_27_47# _142_ 0.043054f
C1859 _032_ counter\[15\] 0.056568f
C1860 counter\[7\] hold6/a_285_47# 0.010734f
C1861 VGND hold1/a_49_47# 0.029031f
C1862 VPWR counter\[5\] 0.407694f
C1863 net11 VGND 0.397134f
C1864 net14 counter\[5\] 0.025348f
C1865 _071_ r2r_out[3] 0.650161f
C1866 _112_ clknet_0_clk 0.03298f
C1867 clkbuf_0_clk/a_110_47# net1 0.013819f
C1868 _330_/a_466_413# _006_ 0.029008f
C1869 VPWR _281_/a_27_47# 0.055701f
C1870 counter\[4\] _206_/a_113_297# 0.052104f
C1871 _298_/a_103_199# clkbuf_2_2__f_clk/a_110_47# 0.012341f
C1872 net6 _328_/a_634_159# 0.046582f
C1873 clknet_0_clk counter\[15\] 0.316781f
C1874 net7 net10 0.359631f
C1875 VGND _076_ -0.013647f
C1876 _057_ _179_/a_79_21# 0.015932f
C1877 _036_ _034_ 0.272114f
C1878 _097_ _098_ 0.017499f
C1879 counter\[2\] _099_ 0.235282f
C1880 VPWR _100_ 0.225809f
C1881 _126_ _117_ 0.015879f
C1882 _125_ _078_ 0.037444f
C1883 _149_ data[2] 0.079745f
C1884 load_divider ext_data 0.044567f
C1885 divider\[1\] clknet_2_3__leaf_clk 0.350491f
C1886 _060_ counter\[9\] 0.129935f
C1887 net4 _065_ 0.020849f
C1888 VPWR _337_/a_634_183# 0.024113f
C1889 clkbuf_2_3__f_clk/a_110_47# _060_ 0.279501f
C1890 net13 VGND 0.043667f
C1891 VGND net17 0.052051f
C1892 _305_/a_27_47# _309_/a_27_47# 0.010693f
C1893 _053_ _174_/a_79_21# 0.028617f
C1894 clknet_0_clk _052_ 0.487457f
C1895 VPWR divider\[2\] 0.58607f
C1896 counter\[15\] _281_/a_109_297# 0.046654f
C1897 r2r_out[3] _060_ 0.26491f
C1898 _253_/a_79_21# net4 0.016807f
C1899 _094_ _344_/a_466_413# 0.033115f
C1900 _057_ _338_/a_891_413# 0.013944f
C1901 _241_/a_59_75# _117_ 0.024845f
C1902 _053_ _143_ 0.058331f
C1903 _070_ _067_ 0.026106f
C1904 VPWR n_rst 0.298149f
C1905 _173_/a_27_47# _079_ 0.125549f
C1906 _053_ _141_ 0.088866f
C1907 _152_ VGND 0.198692f
C1908 VPWR input4/a_27_47# 0.065274f
C1909 data[0] VPWR 0.271629f
C1910 counter\[6\] _211_/a_27_47# 0.013456f
C1911 r2r_out[1] _063_ 0.094459f
C1912 _101_ net16 0.046551f
C1913 _110_ _065_ 0.521225f
C1914 _326_/a_27_47# _357_/a_27_47# 0.081178f
C1915 VPWR _084_ 0.074022f
C1916 _149_ hold1/a_285_47# 0.043283f
C1917 counter\[5\] _116_ 0.037534f
C1918 _157_ net8 0.273055f
C1919 _057_ _335_/a_634_183# 0.020153f
C1920 _078_ _102_ 0.104441f
C1921 VGND _025_ 0.189791f
C1922 VPWR _123_ 0.215726f
C1923 _265_/a_298_297# _148_ 0.032742f
C1924 VGND _342_/a_193_47# -0.099556f
C1925 VPWR _342_/a_27_47# 0.028073f
C1926 divider\[5\] net10 0.058516f
C1927 VGND _078_ 2.3832f
C1928 VPWR _117_ 0.508444f
C1929 net19 _093_ 0.072539f
C1930 _238_/a_77_199# _035_ 0.011847f
C1931 _053_ _164_/a_215_47# 0.01267f
C1932 _066_ _032_ 0.054074f
C1933 _057_ _333_/a_193_47# 0.383626f
C1934 VGND _018_ 0.192756f
C1935 _060_ _147_ 0.101435f
C1936 _351_/a_466_413# VPWR 0.015481f
C1937 _351_/a_1059_315# VGND 0.023415f
C1938 VGND _051_ 0.536125f
C1939 net6 _079_ 0.024093f
C1940 _007_ net10 0.02763f
C1941 _155_ net10 0.193725f
C1942 _091_ clknet_2_3__leaf_clk 0.030623f
C1943 VGND _247_/a_27_47# 0.06338f
C1944 clknet_0_clk _066_ 0.078233f
C1945 _070_ net2 0.026435f
C1946 clkbuf_2_0__f_clk/a_110_47# _094_ 0.105697f
C1947 _070_ net9 0.020303f
C1948 _149_ counter\[4\] 0.512328f
C1949 _291_/a_109_297# divider\[5\] 0.020543f
C1950 _273_/a_215_53# data[6] 0.065536f
C1951 _111_ net13 0.038658f
C1952 divider\[6\] _038_ 0.235684f
C1953 counter\[10\] counter\[11\] 0.224267f
C1954 clkbuf_2_1__f_clk/a_110_47# _064_ 0.012513f
C1955 _356_/a_634_159# net1 0.01719f
C1956 _346_/a_193_47# VPWR 0.047299f
C1957 _346_/a_634_159# VGND 0.018872f
C1958 counter\[15\] _078_ 0.027225f
C1959 _348_/a_466_413# VGND 0.019797f
C1960 counter\[13\] divider\[2\] 0.107019f
C1961 _200_/a_227_47# counter\[3\] 0.07088f
C1962 _066_ hold1/a_49_47# 0.051272f
C1963 _027_ VPWR 0.045731f
C1964 _053_ _340_/a_27_47# 0.055418f
C1965 _188_/a_27_47# _117_ 0.010253f
C1966 _057_ _032_ 0.021817f
C1967 divider\[1\] net2 0.182145f
C1968 _350_/a_193_47# _026_ 0.021205f
C1969 _142_ _354_/a_1059_315# 0.05569f
C1970 _170_/a_81_21# clknet_2_3__leaf_clk 0.048163f
C1971 _040_ _042_ 0.161112f
C1972 net6 _086_ 0.034014f
C1973 _066_ _076_ 0.036646f
C1974 clknet_0_clk _057_ 0.642016f
C1975 hold1/a_285_47# _065_ 0.014378f
C1976 _052_ _078_ 0.076172f
C1977 divider\[4\] clknet_2_2__leaf_clk 1.126392f
C1978 _101_ _102_ 0.097055f
C1979 _290_/a_27_413# _043_ 0.034818f
C1980 _052_ _051_ 0.123583f
C1981 clknet_0_clk clkbuf_0_clk/a_110_47# 0.026363f
C1982 VGND _101_ 1.369751f
C1983 _024_ VGND 0.282323f
C1984 _117_ _116_ 0.072011f
C1985 _114_ _117_ 0.026137f
C1986 clkbuf_2_3__f_clk/a_110_47# net1 0.023667f
C1987 net7 _258_/a_27_47# 0.015404f
C1988 _136_ _137_ 0.090823f
C1989 _094_ _133_ 0.31982f
C1990 _122_ _120_ 0.21204f
C1991 _292_/a_85_193# _035_ 0.010334f
C1992 net15 _130_ 0.132202f
C1993 _223_/a_93_21# counter\[8\] 0.014117f
C1994 net13 _066_ 0.143786f
C1995 VPWR hold6/a_285_47# 0.028169f
C1996 VGND hold6/a_391_47# -0.010925f
C1997 clkbuf_2_3__f_clk/a_110_47# net5 0.010255f
C1998 clkbuf_2_0__f_clk/a_110_47# clknet_2_0__leaf_clk 0.218368f
C1999 r2r_out[4] _065_ 0.387397f
C2000 VPWR _235_/a_113_297# 0.064635f
C2001 _021_ _108_ 0.026376f
C2002 net4 data[3] 0.032881f
C2003 _148_ clknet_2_3__leaf_clk 0.216915f
C2004 _336_/a_475_413# _057_ 0.018609f
C2005 _065_ _019_ 0.012539f
C2006 _336_/a_27_47# clk 0.034212f
C2007 counter\[4\] _065_ 0.044965f
C2008 _112_ _101_ 0.267082f
C2009 _034_ _041_ 0.049798f
C2010 _057_ _076_ 0.050776f
C2011 _352_/a_27_47# _352_/a_466_413# -0.013083f
C2012 _353_/a_27_47# VGND 0.045785f
C2013 _327_/a_1059_315# clknet_2_2__leaf_clk 0.085985f
C2014 _278_/a_219_297# VGND 0.031042f
C2015 VPWR _058_ 0.30461f
C2016 _057_ _337_/a_475_413# 0.048881f
C2017 _071_ VPWR 0.29032f
C2018 _275_/a_109_93# net10 0.052671f
C2019 _275_/a_215_53# _158_ 0.033596f
C2020 VPWR _340_/a_193_47# 0.039496f
C2021 _066_ _078_ 0.147828f
C2022 counter\[12\] counter\[8\] 0.213259f
C2023 VPWR _350_/a_27_47# 0.026774f
C2024 _134_ counter\[11\] 0.205487f
C2025 net6 _154_ 0.019963f
C2026 net1 _147_ 0.030756f
C2027 _078_ r2r_out[0] 0.02173f
C2028 _345_/a_27_47# clknet_2_1__leaf_clk 0.011533f
C2029 _003_ net3 0.070159f
C2030 counter\[12\] _141_ 0.216135f
C2031 input9/a_27_47# ext_data 0.038634f
C2032 VPWR _319_/a_29_53# 0.042148f
C2033 _083_ clknet_2_3__leaf_clk 0.075402f
C2034 _354_/a_381_47# clknet_2_2__leaf_clk 0.028508f
C2035 VGND hold10/a_49_47# 0.034385f
C2036 _343_/a_27_47# VGND 0.050049f
C2037 VGND _354_/a_27_47# 0.053747f
C2038 _352_/a_27_47# _028_ 0.074898f
C2039 net10 ext_data 0.163083f
C2040 divider\[1\] _151_ 0.04539f
C2041 _339_/a_193_47# r2r_out[5] 0.01027f
C2042 _043_ _035_ 0.021661f
C2043 _045_ _041_ 0.103963f
C2044 data[2] data[3] 0.038059f
C2045 _300_/a_27_47# VPWR 0.172954f
C2046 net22 _016_ 0.258937f
C2047 _193_/a_113_297# _098_ 0.065426f
C2048 _334_/a_27_47# _056_ 0.010061f
C2049 _252_/a_81_21# counter\[8\] 0.016494f
C2050 VPWR hold8/a_49_47# 0.016746f
C2051 VGND hold8/a_285_47# 0.071952f
C2052 VPWR _197_/a_27_47# -0.010735f
C2053 VPWR _060_ 2.575911f
C2054 VGND net19 0.818158f
C2055 _025_ _057_ 0.021322f
C2056 _123_ _122_ 0.010572f
C2057 r2r_out[6] clk 0.294725f
C2058 _252_/a_81_21# _141_ 0.044428f
C2059 _057_ _078_ 0.045323f
C2060 _148_ _261_/a_215_297# 0.063155f
C2061 _135_ _054_ 0.051496f
C2062 counter\[10\] hold3/a_49_47# 0.018411f
C2063 _076_ _013_ 0.18235f
C2064 _090_ VGND 0.309149f
C2065 _289_/a_76_199# _041_ 0.017395f
C2066 _348_/a_1059_315# _065_ 0.010107f
C2067 VPWR _183_/a_59_75# 0.016374f
C2068 _149_ _353_/a_193_47# 0.014213f
C2069 _148_ net2 0.029463f
C2070 r2r_out[4] _337_/a_891_413# 0.017893f
C2071 _060_ _080_ 0.025392f
C2072 _329_/a_27_47# net10 0.450532f
C2073 _351_/a_193_47# clknet_2_0__leaf_clk 0.029907f
C2074 _279_/a_207_413# net5 0.04074f
C2075 _326_/a_1059_315# data[1] 0.013038f
C2076 _148_ net9 0.065963f
C2077 _321_/a_222_93# r2r_out[2] 0.031792f
C2078 VGND _217_/a_27_47# 0.018044f
C2079 _149_ _113_ 0.330924f
C2080 hold8/a_285_47# counter\[15\] 0.07513f
C2081 _066_ _101_ 0.08287f
C2082 _024_ _066_ 0.027354f
C2083 _149_ _350_/a_634_159# 0.018196f
C2084 _332_/a_381_47# _158_ 0.018127f
C2085 counter\[2\] _100_ 0.019334f
C2086 _097_ clknet_2_1__leaf_clk 0.072781f
C2087 clknet_0_clk counter\[9\] 0.028241f
C2088 _274_/a_298_297# _157_ 0.015487f
C2089 _112_ _217_/a_27_47# 0.015934f
C2090 _207_/a_285_297# _107_ 0.015469f
C2091 _348_/a_27_47# clknet_2_0__leaf_clk 0.509568f
C2092 _149_ _150_ 0.065806f
C2093 VGND counter\[11\] 0.434087f
C2094 VPWR _207_/a_285_297# -0.019355f
C2095 net4 _327_/a_27_47# 0.044421f
C2096 _192_/a_27_47# _097_ 0.067927f
C2097 _265_/a_215_297# net7 0.071394f
C2098 rst net1 0.022173f
C2099 hold7/a_49_47# net1 0.053155f
C2100 net5 rst 0.072628f
C2101 _105_ hold2/a_285_47# 0.032654f
C2102 VPWR _136_ 1.085966f
C2103 _060_ counter\[14\] 1.021455f
C2104 clk _012_ 0.02625f
C2105 VGND _074_ 0.158173f
C2106 net2 input2/a_27_47# 0.015886f
C2107 _072_ clk 0.022129f
C2108 _148_ clknet_2_2__leaf_clk 0.465029f
C2109 data[7] net9 0.031586f
C2110 _074_ _324_/a_68_297# 0.014786f
C2111 counter\[0\] _189_/a_47_47# 0.04434f
C2112 _148_ _260_/a_215_53# 0.04345f
C2113 _313_/a_27_47# _205_/a_215_53# 0.016989f
C2114 _148_ _325_/a_891_413# 0.02217f
C2115 VGND _168_/a_505_21# 0.073197f
C2116 _267_/a_215_297# VGND 0.010429f
C2117 _267_/a_27_413# VPWR 0.059387f
C2118 _003_ input4/a_27_47# 0.010042f
C2119 _048_ _050_ 0.181969f
C2120 _355_/a_381_47# _031_ 0.01624f
C2121 _065_ _056_ 0.447822f
C2122 VGND r2r_out[5] 0.972585f
C2123 _039_ _297_/a_215_47# 0.010447f
C2124 _355_/a_193_47# net1 0.034946f
C2125 VPWR hold4/a_49_47# 0.046838f
C2126 VGND _095_ 0.259421f
C2127 clknet_0_clk _137_ 0.025945f
C2128 _157_ _331_/a_27_47# 0.037443f
C2129 clknet_0_clk counter\[7\] 0.029443f
C2130 _135_ _243_/a_93_21# 0.040117f
C2131 clknet_0_clk _147_ 0.079924f
C2132 _094_ _313_/a_27_47# 0.057877f
C2133 hold4/a_391_47# clkbuf_2_1__f_clk/a_110_47# 0.010856f
C2134 _081_ r2r_out[4] 0.037659f
C2135 _035_ _041_ 0.047736f
C2136 _059_ counter\[8\] 0.456003f
C2137 _053_ _335_/a_193_47# 0.037909f
C2138 _343_/a_193_47# _065_ 0.042714f
C2139 rst _088_ 0.037963f
C2140 _006_ net9 0.11376f
C2141 divider\[6\] VGND 0.501179f
C2142 VPWR net1 2.02882f
C2143 _148_ _151_ 0.248815f
C2144 clknet_0_clk _046_ 0.047845f
C2145 _186_/a_113_297# clknet_2_1__leaf_clk 0.011595f
C2146 _052_ counter\[11\] 0.022687f
C2147 _065_ _354_/a_193_47# 0.036822f
C2148 VPWR net5 0.791234f
C2149 VGND _077_ 0.128138f
C2150 _161_ clknet_2_3__leaf_clk 0.214286f
C2151 _053_ _333_/a_27_47# 0.067463f
C2152 hold10/a_285_47# r2r_out[7] 0.029418f
C2153 _054_ clknet_2_3__leaf_clk 0.165366f
C2154 _149_ counter\[3\] 0.042609f
C2155 _325_/a_27_47# net4 0.012201f
C2156 _118_ _119_ 0.024761f
C2157 _309_/a_27_47# _055_ 0.010304f
C2158 _065_ _016_ 0.254354f
C2159 _156_ _272_/a_27_413# 0.013537f
C2160 VPWR _179_/a_79_21# 0.071766f
C2161 _004_ net8 0.031559f
C2162 _060_ _341_/a_466_413# 0.037715f
C2163 _017_ _341_/a_193_47# 0.010208f
C2164 _053_ net3 0.01852f
C2165 _117_ _228_/a_27_47# 0.03801f
C2166 VPWR _246_/a_113_297# 0.037151f
C2167 _136_ counter\[14\] 0.028459f
C2168 _355_/a_27_47# net4 0.076161f
C2169 VGND _244_/a_59_75# 0.024148f
C2170 net6 _329_/a_193_47# 0.039135f
C2171 r2r_out[7] _016_ 0.050387f
C2172 _292_/a_85_193# _041_ 0.089933f
C2173 counter\[9\] _078_ 0.287605f
C2174 divider\[6\] counter\[15\] 0.044284f
C2175 counter\[1\] _189_/a_47_47# 0.031392f
C2176 clkbuf_2_3__f_clk/a_110_47# _078_ 0.044f
C2177 _149_ _267_/a_298_297# 0.034814f
C2178 divider\[6\] _037_ 0.032619f
C2179 VPWR _338_/a_891_413# 0.023945f
C2180 _131_ _133_ 0.015417f
C2181 VGND net4 1.744029f
C2182 VPWR _088_ 0.080566f
C2183 counter\[1\] _096_ 0.056445f
C2184 _066_ counter\[11\] 0.015482f
C2185 _328_/a_27_47# clknet_2_2__leaf_clk 0.017569f
C2186 _094_ _207_/a_35_297# 0.022793f
C2187 _351_/a_891_413# counter\[10\] 0.045234f
C2188 _066_ _190_/a_76_199# 0.019236f
C2189 _067_ _054_ 0.033682f
C2190 _036_ _041_ 0.023293f
C2191 _078_ _248_/a_77_199# 0.022047f
C2192 VPWR _156_ 0.402725f
C2193 _094_ hold2/a_391_47# 0.0434f
C2194 _331_/a_193_47# _007_ 0.092164f
C2195 _266_/a_109_93# net10 0.023611f
C2196 VGND _335_/a_475_413# 0.020701f
C2197 _236_/a_27_47# counter\[11\] 0.012063f
C2198 divider\[4\] net7 0.015489f
C2199 _004_ net6 0.244449f
C2200 VGND _283_/a_215_47# 0.041027f
C2201 VGND hold3/a_49_47# 0.022916f
C2202 _124_ counter\[8\] 0.182173f
C2203 _066_ _074_ 0.090789f
C2204 counter\[10\] _129_ 0.271183f
C2205 _329_/a_634_159# net10 0.016209f
C2206 _065_ counter\[3\] 0.26601f
C2207 _137_ _078_ 0.027382f
C2208 _065_ _190_/a_206_369# 0.026522f
C2209 net4 counter\[15\] 0.201672f
C2210 VPWR _333_/a_193_47# 0.039504f
C2211 VGND _333_/a_634_183# 0.016697f
C2212 counter\[7\] _078_ 0.192146f
C2213 _104_ _344_/a_891_413# 0.046639f
C2214 net22 _065_ 0.115017f
C2215 _187_/a_297_47# clknet_2_1__leaf_clk 0.043861f
C2216 VGND _110_ 0.510186f
C2217 VGND _341_/a_27_47# 0.077991f
C2218 _315_/a_27_47# _054_ 0.0289f
C2219 _066_ r2r_out[5] 0.036802f
C2220 divider\[2\] _327_/a_634_159# 0.041092f
C2221 divider\[6\] _273_/a_109_93# 0.020508f
C2222 _078_ _046_ 0.06557f
C2223 VPWR _349_/a_381_47# 0.020498f
C2224 r2r_out[3] _321_/a_79_199# 0.079631f
C2225 net22 r2r_out[7] 0.054639f
C2226 net16 _019_ 0.038508f
C2227 VPWR _328_/a_1059_315# 0.033111f
C2228 _065_ clkbuf_2_1__f_clk/a_110_47# 0.017309f
C2229 _149_ _271_/a_29_53# 0.011768f
C2230 VGND _347_/a_27_47# 0.1029f
C2231 _051_ _046_ 0.040701f
C2232 net11 rst 0.037159f
C2233 net2 _054_ 2.532385f
C2234 _054_ net9 0.406577f
C2235 _338_/a_27_47# _338_/a_475_413# -0.013973f
C2236 divider\[1\] net7 0.085171f
C2237 _136_ _122_ 0.024602f
C2238 net10 input7/a_27_47# 0.018742f
C2239 net8 net3 0.025663f
C2240 _247_/a_27_47# _046_ 0.019296f
C2241 VGND data[2] 0.050693f
C2242 _181_/a_93_21# _088_ 0.033428f
C2243 _083_ _338_/a_634_183# 0.016097f
C2244 net8 _328_/a_466_413# 0.032988f
C2245 _348_/a_381_47# _024_ 0.018928f
C2246 _066_ _077_ 0.059513f
C2247 _353_/a_466_413# _078_ 0.032527f
C2248 VPWR _032_ 0.136244f
C2249 _334_/a_27_47# _065_ 0.04389f
C2250 _121_ _132_ 0.034088f
C2251 _066_ _163_/a_27_47# 0.049393f
C2252 counter\[2\] _197_/a_27_47# 0.036039f
C2253 VPWR _329_/a_1059_315# 0.051977f
C2254 _251_/a_27_47# _136_ 0.015169f
C2255 _057_ r2r_out[5] 0.033573f
C2256 divider\[4\] divider\[5\] 0.028611f
C2257 clknet_0_clk VPWR 1.576429f
C2258 hold5/a_285_47# _099_ 0.034088f
C2259 _278_/a_219_297# counter\[9\] 0.019037f
C2260 _326_/a_27_47# _002_ 0.024044f
C2261 _054_ _121_ 0.182124f
C2262 _066_ _244_/a_59_75# 0.04115f
C2263 counter\[0\] _195_/a_77_199# 0.082402f
C2264 divider\[4\] _155_ 0.196549f
C2265 VPWR _234_/a_113_297# 0.075251f
C2266 VPWR _345_/a_891_413# 0.016564f
C2267 _067_ clknet_2_3__leaf_clk 0.025454f
C2268 _149_ _065_ 0.696259f
C2269 VPWR hold1/a_49_47# 0.054549f
C2270 VGND hold1/a_285_47# -0.015926f
C2271 _053_ _123_ 0.241873f
C2272 _336_/a_1062_300# VGND -0.017147f
C2273 _157_ net10 0.03905f
C2274 net11 VPWR 0.152123f
C2275 _152_ rst 0.018119f
C2276 _332_/a_27_47# _276_/a_27_413# 0.012449f
C2277 _260_/a_215_53# _054_ 0.01176f
C2278 input1/a_27_47# net12 0.06673f
C2279 net6 net3 0.024384f
C2280 VGND data[6] 0.222751f
C2281 _066_ net4 1.04277f
C2282 _326_/a_193_47# _326_/a_634_159# -0.016573f
C2283 net6 _328_/a_466_413# 0.039639f
C2284 VGND r2r_out[4] 1.124468f
C2285 VPWR _076_ 0.090844f
C2286 counter\[0\] _099_ 0.368704f
C2287 _071_ _318_/a_27_47# 0.062359f
C2288 r2r_out[6] _091_ 0.022422f
C2289 _188_/a_27_47# clknet_0_clk 0.04217f
C2290 _223_/a_93_21# _120_ 0.039897f
C2291 VGND _019_ 0.096487f
C2292 _126_ _078_ 0.385136f
C2293 _048_ net9 1.128161f
C2294 _057_ _244_/a_59_75# 0.048452f
C2295 VGND counter\[4\] 1.338996f
C2296 VGND _337_/a_1062_300# 0.07466f
C2297 VPWR _337_/a_475_413# 0.023585f
C2298 net13 VPWR 0.095132f
C2299 VPWR net17 0.17467f
C2300 _335_/a_1062_300# r2r_out[2] 0.018246f
C2301 VGND _034_ 0.797782f
C2302 counter\[15\] _281_/a_193_297# 0.05613f
C2303 net2 clknet_2_3__leaf_clk 0.146565f
C2304 _094_ _344_/a_1059_315# 0.049095f
C2305 clknet_2_3__leaf_clk net9 0.569015f
C2306 _066_ _110_ 0.0263f
C2307 _082_ _060_ 0.234289f
C2308 counter\[6\] _216_/a_59_75# 0.067084f
C2309 _308_/a_27_47# _059_ 0.023154f
C2310 _057_ net4 0.249253f
C2311 _060_ _255_/a_80_21# 0.040468f
C2312 clknet_0_clk counter\[14\] 0.776419f
C2313 _173_/a_109_297# _079_ 0.022112f
C2314 clknet_0_clk counter\[13\] 0.017531f
C2315 _112_ counter\[4\] 0.039589f
C2316 _152_ VPWR 0.24881f
C2317 counter\[1\] _195_/a_77_199# 0.026605f
C2318 net8 divider\[2\] 0.023821f
C2319 _065_ r2r_out[2] 0.029617f
C2320 _328_/a_27_47# _328_/a_193_47# -0.015164f
C2321 _060_ _318_/a_27_47# 0.013042f
C2322 _356_/a_27_47# VGND 0.051452f
C2323 _110_ _022_ 0.0167f
C2324 _111_ hold1/a_285_47# 0.012522f
C2325 _149_ hold1/a_391_47# 0.056021f
C2326 _070_ _301_/a_27_47# 0.010433f
C2327 _353_/a_27_47# _353_/a_466_413# -0.013083f
C2328 _057_ _335_/a_475_413# 0.013013f
C2329 _040_ _051_ 0.035183f
C2330 VPWR _025_ 0.510222f
C2331 _056_ _009_ 0.052545f
C2332 VGND _342_/a_634_159# 0.01472f
C2333 VPWR _342_/a_193_47# 0.020179f
C2334 _048_ clknet_2_2__leaf_clk 0.075367f
C2335 _154_ net10 0.083116f
C2336 VGND _118_ 0.431394f
C2337 VPWR _078_ 6.048347f
C2338 _238_/a_77_199# _134_ 0.01025f
C2339 _339_/a_27_47# _339_/a_193_47# -0.01246f
C2340 r2r_out[7] _065_ 0.029904f
C2341 _057_ _333_/a_634_183# 0.037832f
C2342 _208_/a_76_199# counter\[5\] 0.033423f
C2343 VPWR _018_ 0.10571f
C2344 _351_/a_1059_315# VPWR 0.047689f
C2345 VGND _045_ 0.153505f
C2346 VPWR _051_ 0.579877f
C2347 clknet_2_3__leaf_clk net12 0.011907f
C2348 _148_ net7 1.264987f
C2349 counter\[9\] counter\[11\] 0.016412f
C2350 counter\[1\] _099_ 0.536652f
C2351 _292_/a_516_297# _042_ 0.011415f
C2352 VPWR _247_/a_27_47# 0.025038f
C2353 VGND _064_ 0.042171f
C2354 VPWR _061_ 0.150032f
C2355 _356_/a_27_47# counter\[15\] 0.428633f
C2356 _066_ _169_/a_51_297# 0.023977f
C2357 VGND _129_ 0.021987f
C2358 _112_ _118_ 0.0186f
C2359 _184_/a_27_47# clknet_2_3__leaf_clk 0.045794f
C2360 _273_/a_109_93# data[6] 0.039456f
C2361 _311_/a_27_297# _062_ 0.042737f
C2362 net6 divider\[2\] 0.031947f
C2363 VGND _289_/a_76_199# 0.028509f
C2364 _346_/a_634_159# VPWR 0.035817f
C2365 _346_/a_466_413# VGND 0.019314f
C2366 _053_ _058_ 0.026885f
C2367 _348_/a_1059_315# VGND 0.024438f
C2368 _111_ _219_/a_77_199# 0.029617f
C2369 _291_/a_193_297# _155_ 0.023265f
C2370 divider\[1\] _327_/a_381_47# 0.016521f
C2371 _200_/a_227_47# _102_ 0.010979f
C2372 r2r_out[3] _074_ 0.019298f
C2373 _066_ hold1/a_285_47# 0.069697f
C2374 _053_ _071_ 0.121695f
C2375 _053_ _340_/a_193_47# 0.045505f
C2376 r2r_out[1] _054_ 0.129711f
C2377 net2 _315_/a_27_47# 0.010498f
C2378 _315_/a_27_47# net9 0.034631f
C2379 _149_ data[3] 0.098917f
C2380 _142_ _354_/a_891_413# 0.04226f
C2381 _187_/a_79_21# _060_ 0.059746f
C2382 _053_ _319_/a_29_53# 0.06236f
C2383 VPWR _321_/a_79_199# 0.023531f
C2384 _151_ clknet_2_3__leaf_clk 0.078982f
C2385 _356_/a_193_47# _149_ 0.015445f
C2386 _066_ r2r_out[4] 0.487448f
C2387 net6 _084_ 0.160806f
C2388 _266_/a_215_53# _153_ 0.016576f
C2389 _031_ _143_ 0.36264f
C2390 _107_ _101_ 0.019925f
C2391 _031_ _141_ 0.151652f
C2392 _290_/a_207_413# _043_ 0.077037f
C2393 _057_ _169_/a_51_297# 0.056586f
C2394 net2 net9 0.024235f
C2395 _052_ _045_ 0.036862f
C2396 VPWR _101_ 2.146236f
C2397 _094_ _021_ 0.057733f
C2398 _066_ counter\[4\] 0.305976f
C2399 _024_ VPWR 0.600987f
C2400 _044_ _155_ 0.023715f
C2401 _269_/a_215_297# net5 0.019377f
C2402 _197_/a_27_47# _103_ 0.098113f
C2403 _223_/a_250_297# counter\[8\] 0.010701f
C2404 VPWR hold6/a_391_47# 0.013125f
C2405 counter\[13\] _078_ 0.452783f
C2406 hold10/a_49_47# rst 0.063033f
C2407 _326_/a_193_47# VGND -0.109622f
C2408 _326_/a_27_47# VPWR 0.035451f
C2409 counter\[14\] _051_ 0.026122f
C2410 _053_ _060_ 0.062484f
C2411 divider\[4\] _329_/a_27_47# 0.03226f
C2412 _281_/a_27_47# _280_/a_27_413# 0.011041f
C2413 _336_/a_1062_300# _057_ 0.01135f
C2414 _320_/a_80_21# VPWR 0.061152f
C2415 input6/a_27_47# data[5] 0.017763f
C2416 counter\[13\] _051_ 0.664224f
C2417 _148_ _007_ 0.096036f
C2418 divider\[0\] _261_/a_27_413# 0.039492f
C2419 _354_/a_27_47# _030_ 0.027484f
C2420 _345_/a_193_47# _345_/a_634_159# -0.016573f
C2421 _336_/a_193_47# clk 0.386797f
C2422 counter\[13\] _247_/a_27_47# 0.054929f
C2423 _031_ _250_/a_113_297# 0.136559f
C2424 _307_/a_59_75# _133_ 0.066491f
C2425 _057_ r2r_out[4] 0.113443f
C2426 _081_ _178_/a_75_199# 0.105656f
C2427 _353_/a_193_47# VGND -0.099938f
C2428 _353_/a_27_47# VPWR -0.131083f
C2429 _327_/a_891_413# clknet_2_2__leaf_clk 0.044932f
C2430 _278_/a_27_53# VGND 0.037374f
C2431 VGND _056_ 0.191218f
C2432 _227_/a_59_75# _124_ 0.048317f
C2433 _057_ _337_/a_1062_300# 0.012013f
C2434 _339_/a_27_47# VGND 0.02057f
C2435 _090_ rst 0.199156f
C2436 _357_/a_1283_21# _000_ 0.038095f
C2437 _094_ _115_ 0.03691f
C2438 VPWR _350_/a_193_47# 0.014167f
C2439 net9 clknet_2_2__leaf_clk 0.386419f
C2440 _345_/a_27_47# _021_ 0.059951f
C2441 _094_ _096_ 0.057011f
C2442 VPWR hold10/a_49_47# 0.054079f
C2443 VGND _035_ 0.864187f
C2444 _343_/a_193_47# VGND -0.099626f
C2445 _343_/a_27_47# VPWR 0.046554f
C2446 divider\[3\] _035_ 0.377584f
C2447 _169_/a_51_297# _013_ 0.028098f
C2448 _356_/a_1059_315# net3 0.028049f
C2449 _120_ _059_ 0.054157f
C2450 _236_/a_27_47# _045_ 0.012266f
C2451 divider\[4\] _159_ 0.058665f
C2452 _101_ _116_ 0.135898f
C2453 VPWR _354_/a_27_47# -0.03986f
C2454 _352_/a_193_47# _028_ 0.106315f
C2455 _065_ _119_ 0.119631f
C2456 _149_ _093_ 0.232976f
C2457 _112_ _113_ 0.080469f
C2458 _066_ _129_ 0.023661f
C2459 VGND _150_ 0.087021f
C2460 VGND _016_ 0.143169f
C2461 VPWR hold8/a_285_47# 0.02871f
C2462 VGND hold8/a_391_47# 0.014657f
C2463 VPWR net19 0.186885f
C2464 VGND _017_ 0.277207f
C2465 _126_ counter\[11\] 0.092342f
C2466 _148_ _261_/a_298_297# 0.013369f
C2467 counter\[15\] _035_ 0.131376f
C2468 _132_ _133_ 0.062757f
C2469 _090_ _092_ 0.07959f
C2470 r2r_out[4] _013_ 0.388803f
C2471 hold4/a_391_47# net16 0.011273f
C2472 _289_/a_226_47# _041_ 0.040709f
C2473 _346_/a_466_413# _022_ 0.010537f
C2474 VGND _245_/a_75_212# 0.013878f
C2475 clknet_2_1__leaf_clk _054_ 0.022245f
C2476 _052_ _113_ 0.029635f
C2477 _081_ _065_ 0.095749f
C2478 clknet_2_0__leaf_clk _115_ 0.017828f
C2479 _054_ _133_ 0.042228f
C2480 divider\[1\] _159_ 0.029846f
C2481 counter\[10\] _065_ 0.028437f
C2482 _329_/a_193_47# net10 0.057512f
C2483 VPWR _217_/a_27_47# 0.013235f
C2484 _111_ _113_ 0.042933f
C2485 hold8/a_391_47# counter\[15\] 0.072277f
C2486 _149_ _350_/a_466_413# 0.011263f
C2487 _146_ _143_ 0.032261f
C2488 _173_/a_27_47# _060_ 0.012787f
C2489 _280_/a_207_413# counter\[8\] 0.022446f
C2490 _053_ net1 0.025038f
C2491 _004_ _001_ 0.01259f
C2492 _101_ _106_ 0.028418f
C2493 counter\[0\] _100_ 0.048001f
C2494 VGND _036_ 0.269721f
C2495 VGND _332_/a_27_47# 0.060223f
C2496 counter\[3\] _102_ 0.428204f
C2497 net7 _054_ 0.076648f
C2498 _346_/a_27_47# clknet_2_0__leaf_clk 0.012547f
C2499 net17 counter\[2\] 0.058854f
C2500 _348_/a_193_47# clknet_2_0__leaf_clk 0.100673f
C2501 _048_ _297_/a_79_21# 0.02368f
C2502 _069_ r2r_out[2] 0.041031f
C2503 VPWR counter\[11\] 2.436851f
C2504 VGND counter\[3\] 0.452119f
C2505 net4 _327_/a_193_47# 0.040124f
C2506 _053_ _179_/a_79_21# 0.026977f
C2507 divider\[6\] rst 1.276404f
C2508 _148_ divider\[0\] 0.389362f
C2509 hold7/a_285_47# net1 0.091277f
C2510 _040_ _047_ 0.268036f
C2511 net22 VGND 0.91898f
C2512 net6 _060_ 0.073777f
C2513 _105_ hold2/a_391_47# 0.028675f
C2514 clknet_0_clk _255_/a_80_21# 0.103539f
C2515 VPWR _074_ 0.079008f
C2516 _056_ r2r_out[0] 0.434611f
C2517 _066_ _113_ 0.014163f
C2518 r2r_out[1] net2 0.021271f
C2519 VGND _043_ 0.607833f
C2520 VPWR _047_ 0.157518f
C2521 _036_ counter\[15\] 0.067291f
C2522 _336_/a_27_47# clknet_2_3__leaf_clk 0.018217f
C2523 _336_/a_1062_300# hold9/a_49_47# 0.019949f
C2524 _148_ _262_/a_215_53# 0.040395f
C2525 VGND clkbuf_2_1__f_clk/a_110_47# -0.017427f
C2526 _336_/a_1062_300# r2r_out[3] 0.033322f
C2527 VPWR _168_/a_505_21# 0.106701f
C2528 _267_/a_215_297# VPWR 0.012425f
C2529 _027_ _128_ 0.034185f
C2530 _071_ _068_ 0.171916f
C2531 _053_ _088_ 0.034081f
C2532 VPWR r2r_out[5] 1.404652f
C2533 VPWR hold4/a_285_47# 0.01042f
C2534 VGND hold4/a_391_47# -0.010796f
C2535 VPWR _095_ 0.057062f
C2536 divider\[4\] _329_/a_634_159# 0.020951f
C2537 _094_ _142_ 0.103397f
C2538 _171_/a_27_47# r2r_out[5] 0.011474f
C2539 _148_ _329_/a_27_47# 0.010534f
C2540 _157_ _331_/a_193_47# 0.034136f
C2541 VGND divider\[7\] 0.8958f
C2542 _136_ _223_/a_93_21# 0.020206f
C2543 _014_ r2r_out[5] 0.170142f
C2544 _033_ counter\[8\] 0.063879f
C2545 r2r_out[3] r2r_out[4] 0.178547f
C2546 data[7] ext_data 0.041759f
C2547 counter\[1\] _100_ 0.222454f
C2548 _337_/a_27_47# clknet_2_3__leaf_clk 0.017772f
C2549 counter\[9\] _034_ 0.207652f
C2550 _134_ _065_ 0.094591f
C2551 _343_/a_634_159# _065_ 0.012f
C2552 net4 rst 0.017836f
C2553 r2r_out[7] _340_/a_1062_300# 0.020769f
C2554 _060_ _349_/a_27_47# 0.011123f
C2555 divider\[6\] VPWR 1.403566f
C2556 _149_ _355_/a_27_47# 0.022657f
C2557 _091_ _085_ 0.029738f
C2558 _339_/a_27_47# _057_ 0.037793f
C2559 r2r_out[5] _080_ 0.033244f
C2560 _065_ _354_/a_634_159# 0.013241f
C2561 VPWR _077_ 0.469242f
C2562 _057_ _340_/a_475_413# 0.013618f
C2563 _053_ _333_/a_193_47# 0.272585f
C2564 hold10/a_391_47# r2r_out[7] 0.018835f
C2565 VGND _178_/a_75_199# 0.014741f
C2566 _094_ _195_/a_77_199# 0.031262f
C2567 _303_/a_113_297# net1 0.019125f
C2568 _149_ _102_ 0.20913f
C2569 net8 net1 0.02577f
C2570 _094_ _229_/a_227_47# 0.014251f
C2571 _072_ _054_ 0.187752f
C2572 VPWR _163_/a_27_47# 0.040039f
C2573 counter\[13\] counter\[11\] 0.02964f
C2574 _066_ _245_/a_75_212# 0.013757f
C2575 _223_/a_250_297# _308_/a_27_47# 0.044818f
C2576 divider\[7\] counter\[15\] 0.919434f
C2577 net8 net5 0.019903f
C2578 _149_ VGND 3.237053f
C2579 _133_ _248_/a_227_47# 0.012737f
C2580 _060_ _341_/a_1059_315# 0.068002f
C2581 _149_ divider\[3\] 0.237408f
C2582 _078_ _228_/a_27_47# 0.018741f
C2583 _065_ _176_/a_68_297# 0.010383f
C2584 _355_/a_193_47# net4 0.170904f
C2585 VPWR _244_/a_59_75# 0.010023f
C2586 net7 clknet_2_3__leaf_clk 0.026686f
C2587 _080_ _077_ 0.065015f
C2588 _136_ counter\[12\] 0.119511f
C2589 _334_/a_27_47# _334_/a_193_47# -0.078191f
C2590 _124_ _117_ 0.078325f
C2591 r2r_out[6] clknet_2_3__leaf_clk 0.029845f
C2592 VGND _271_/a_29_53# 0.037231f
C2593 _047_ counter\[13\] 0.035156f
C2594 net6 _168_/a_76_199# 0.06097f
C2595 _101_ counter\[2\] 0.044148f
C2596 VPWR net4 0.777394f
C2597 _149_ counter\[15\] 0.023022f
C2598 _297_/a_79_21# net9 0.016458f
C2599 _328_/a_193_47# clknet_2_2__leaf_clk 0.013799f
C2600 _351_/a_381_47# counter\[10\] 0.022282f
C2601 _053_ clknet_0_clk 0.042718f
C2602 net6 net1 0.024201f
C2603 divider\[6\] counter\[14\] 0.138406f
C2604 VGND _335_/a_1062_300# 0.074069f
C2605 net6 net5 0.284274f
C2606 _045_ _248_/a_77_199# 0.014154f
C2607 VGND hold3/a_285_47# 0.014532f
C2608 VPWR hold3/a_49_47# 0.035069f
C2609 _060_ _169_/a_240_47# 0.036574f
C2610 VGND r2r_out[2] 1.678056f
C2611 _329_/a_466_413# net10 0.033063f
C2612 _065_ _102_ 0.018045f
C2613 _301_/a_27_47# _054_ 0.031999f
C2614 net8 _156_ 0.069071f
C2615 VPWR _333_/a_634_183# 0.014792f
C2616 _053_ _336_/a_475_413# 0.042726f
C2617 _104_ _344_/a_381_47# 0.01471f
C2618 VGND _041_ 0.679179f
C2619 VPWR _110_ 0.15254f
C2620 VGND _065_ 6.477661f
C2621 _149_ _111_ 0.275087f
C2622 VPWR _341_/a_27_47# 0.065974f
C2623 VGND _341_/a_193_47# -0.080631f
C2624 divider\[3\] _041_ 0.029509f
C2625 divider\[2\] _327_/a_466_413# 0.024505f
C2626 r2r_out[3] _321_/a_222_93# 0.027155f
C2627 clknet_2_3__leaf_clk _012_ 0.059677f
C2628 VGND r2r_out[7] 1.247787f
C2629 _060_ _059_ 0.012503f
C2630 _253_/a_79_21# VGND -0.018679f
C2631 VGND _347_/a_193_47# -0.10118f
C2632 VPWR _347_/a_27_47# 0.086594f
C2633 _045_ _046_ 0.229664f
C2634 _072_ clknet_2_3__leaf_clk 0.735001f
C2635 _343_/a_27_47# counter\[2\] 0.052487f
C2636 _297_/a_79_21# clknet_2_2__leaf_clk 0.025965f
C2637 _338_/a_193_47# _338_/a_475_413# -0.01259f
C2638 rst data[6] 0.062323f
C2639 VPWR data[2] 0.260113f
C2640 _053_ _337_/a_475_413# 0.018897f
C2641 _083_ _338_/a_475_413# 0.028739f
C2642 net8 _328_/a_1059_315# 0.053842f
C2643 net6 _088_ 0.126862f
C2644 _353_/a_1059_315# _078_ 0.052631f
C2645 net4 counter\[14\] 0.149643f
C2646 _072_ _164_/a_79_21# 0.014728f
C2647 net2 net7 0.467853f
C2648 net7 net9 0.517376f
C2649 _121_ _133_ 0.035581f
C2650 counter\[0\] _197_/a_27_47# 0.047081f
C2651 VPWR _329_/a_891_413# 0.028599f
C2652 _066_ _163_/a_109_297# 0.033201f
C2653 clknet_2_1__leaf_clk _098_ 0.036863f
C2654 _060_ counter\[0\] 0.274401f
C2655 r2r_out[6] net9 0.018052f
C2656 _187_/a_79_21# _078_ 0.010272f
C2657 net6 _156_ 0.107962f
C2658 divider\[4\] _154_ 0.019148f
C2659 _149_ _066_ 0.455076f
C2660 hold5/a_391_47# _099_ 0.041195f
C2661 _278_/a_27_53# counter\[9\] 0.077837f
C2662 divider\[0\] _161_ 0.120642f
C2663 VPWR _169_/a_51_297# 0.043486f
C2664 _326_/a_193_47# _002_ 0.385725f
C2665 _097_ _195_/a_77_199# 0.010753f
C2666 divider\[2\] net10 0.028857f
C2667 divider\[0\] _054_ 0.118952f
C2668 _309_/a_27_47# _060_ 0.043251f
C2669 _021_ hold2/a_49_47# 0.014738f
C2670 data[4] data[5] 0.039497f
C2671 _078_ _103_ 0.011774f
C2672 _111_ _065_ 0.073197f
C2673 _051_ _354_/a_1059_315# 0.011201f
C2674 _053_ _025_ 0.152131f
C2675 VGND hold1/a_391_47# -0.012015f
C2676 VPWR hold1/a_285_47# 0.089225f
C2677 _336_/a_1062_300# VPWR 0.091239f
C2678 _336_/a_891_413# VGND -0.013271f
C2679 _053_ _078_ 0.114094f
C2680 _144_ VGND 0.106239f
C2681 _260_/a_109_93# _054_ 0.023217f
C2682 VPWR _281_/a_193_297# -0.018684f
C2683 VPWR data[6] 0.132476f
C2684 divider\[1\] counter\[8\] 0.738235f
C2685 net6 _328_/a_1059_315# 0.060323f
C2686 _301_/a_27_47# clknet_2_3__leaf_clk 0.037309f
C2687 _136_ _059_ 0.030508f
C2688 VPWR r2r_out[4] 1.176126f
C2689 _149_ _057_ 0.018413f
C2690 _053_ _061_ 0.049438f
C2691 _107_ counter\[4\] 0.412817f
C2692 VPWR _019_ 0.283407f
C2693 net7 clknet_2_2__leaf_clk 0.130827f
C2694 _171_/a_27_47# r2r_out[4] 0.029325f
C2695 _065_ _087_ 0.024607f
C2696 _294_/a_215_47# _045_ 0.041815f
C2697 VPWR counter\[4\] 1.635923f
C2698 VPWR _337_/a_1062_300# 0.080398f
C2699 VGND _337_/a_891_413# 0.021962f
C2700 _105_ _021_ 0.096998f
C2701 VGND _177_/a_59_75# 0.059752f
C2702 _035_ _248_/a_77_199# 0.01315f
C2703 divider\[5\] net9 0.034913f
C2704 _053_ _174_/a_215_47# 0.014675f
C2705 VPWR _034_ 0.057175f
C2706 counter\[1\] _197_/a_27_47# 0.049235f
C2707 r2r_out[2] r2r_out[0] 1.158713f
C2708 net6 _329_/a_1059_315# 0.014615f
C2709 _094_ _344_/a_891_413# 0.034485f
C2710 _066_ _065_ 1.982777f
C2711 _126_ _129_ 0.137684f
C2712 _060_ _255_/a_209_297# 0.04038f
C2713 _065_ r2r_out[0] 0.221974f
C2714 clknet_0_clk counter\[12\] 0.147528f
C2715 _338_/a_1062_300# clk 0.020674f
C2716 VGND input10/a_27_47# 0.035923f
C2717 _053_ _321_/a_79_199# 0.036f
C2718 VGND data[3] 0.049238f
C2719 net7 _151_ 0.01808f
C2720 _240_/a_68_297# counter\[12\] 0.01444f
C2721 VGND _038_ 0.273584f
C2722 _253_/a_79_21# _066_ 0.014955f
C2723 _356_/a_27_47# VPWR -0.143683f
C2724 _101_ _103_ 0.172096f
C2725 _065_ _022_ 0.236422f
C2726 _274_/a_215_297# divider\[6\] 0.011118f
C2727 _341_/a_193_47# _341_/a_634_159# -0.016573f
C2728 _035_ _046_ 0.452656f
C2729 _111_ hold1/a_391_47# 0.017494f
C2730 _067_ _301_/a_27_47# 0.029914f
C2731 _334_/a_381_47# clknet_2_1__leaf_clk 0.021289f
C2732 _256_/a_81_21# _146_ 0.057898f
C2733 _057_ _335_/a_1062_300# 0.012227f
C2734 _040_ _045_ 0.097967f
C2735 _036_ counter\[9\] 0.278979f
C2736 _265_/a_27_413# net5 0.02799f
C2737 _157_ _148_ 0.129093f
C2738 VPWR _342_/a_634_159# 0.018382f
C2739 VPWR _118_ 0.080267f
C2740 VGND _119_ 0.329242f
C2741 _057_ r2r_out[2] 0.031656f
C2742 divider\[0\] clknet_2_3__leaf_clk 0.050365f
C2743 _057_ _333_/a_475_413# 0.041684f
C2744 _208_/a_206_369# counter\[5\] 0.03388f
C2745 _053_ _320_/a_80_21# 0.025718f
C2746 _351_/a_891_413# VPWR 0.022899f
C2747 VPWR _045_ 0.470518f
C2748 _057_ _065_ 0.017519f
C2749 counter\[0\] net1 0.178239f
C2750 counter\[15\] _038_ 0.010603f
C2751 VPWR _064_ 0.151931f
C2752 _007_ clknet_2_2__leaf_clk 0.061966f
C2753 _356_/a_193_47# counter\[15\] 0.055036f
C2754 counter\[4\] _116_ 0.317377f
C2755 _347_/a_193_47# _347_/a_634_159# -0.016573f
C2756 _057_ r2r_out[7] 0.100652f
C2757 _253_/a_79_21# _057_ 0.074583f
C2758 _213_/a_215_53# _115_ 0.043458f
C2759 r2r_out[1] clknet_2_1__leaf_clk 0.061607f
C2760 _292_/a_85_193# _046_ 0.021525f
C2761 _037_ _038_ 0.070309f
C2762 VGND _289_/a_226_47# 0.032753f
C2763 counter\[5\] _212_/a_80_21# 0.01334f
C2764 _346_/a_466_413# VPWR 0.050477f
C2765 _346_/a_1059_315# VGND 0.029362f
C2766 _348_/a_891_413# VGND 0.01202f
C2767 _114_ _219_/a_77_199# 0.093497f
C2768 _200_/a_77_199# _344_/a_1059_315# 0.015723f
C2769 VGND _081_ 0.401976f
C2770 counter\[13\] _034_ 0.028825f
C2771 _301_/a_27_47# net9 0.024705f
C2772 _066_ hold1/a_391_47# 0.060044f
C2773 _094_ counter\[5\] 0.416318f
C2774 counter\[10\] VGND 2.340561f
C2775 _053_ _340_/a_634_183# 0.011828f
C2776 _343_/a_27_47# _103_ 0.011182f
C2777 VPWR _290_/a_27_413# 0.033118f
C2778 _187_/a_79_21# net19 0.011203f
C2779 VGND _005_ 0.062978f
C2780 _347_/a_27_47# _023_ 0.039936f
C2781 _072_ _170_/a_299_297# 0.012902f
C2782 _094_ _100_ 0.027813f
C2783 _263_/a_215_297# net1 0.023161f
C2784 net6 _078_ 0.055357f
C2785 VGND _093_ 0.011664f
C2786 _114_ _118_ 0.041687f
C2787 _111_ _119_ 0.179595f
C2788 _148_ _154_ 0.794131f
C2789 _089_ net9 0.095984f
C2790 counter\[12\] _078_ 0.304904f
C2791 _003_ net4 0.055821f
C2792 hold10/a_285_47# rst 0.09886f
C2793 _326_/a_634_159# VGND 0.024324f
C2794 _326_/a_193_47# VPWR 0.026253f
C2795 _013_ _065_ 0.096722f
C2796 counter\[14\] _045_ 0.0245f
C2797 divider\[4\] _329_/a_193_47# 0.01991f
C2798 _336_/a_891_413# _057_ 0.01015f
C2799 counter\[13\] _045_ 0.057411f
C2800 divider\[0\] _261_/a_215_297# 0.04939f
C2801 VGND _069_ 0.101172f
C2802 _354_/a_193_47# _030_ 0.079022f
C2803 _336_/a_634_183# clk 0.022114f
C2804 _265_/a_215_297# net3 0.016488f
C2805 _082_ _077_ 0.062315f
C2806 counter\[12\] _247_/a_27_47# 0.088036f
C2807 _149_ clkbuf_2_3__f_clk/a_110_47# 0.023462f
C2808 _010_ _061_ 0.010479f
C2809 _290_/a_27_413# _294_/a_78_199# 0.010632f
C2810 _053_ _090_ 0.061583f
C2811 _039_ divider\[6\] 0.075176f
C2812 VPWR _238_/a_77_199# 0.015666f
C2813 rst _016_ 0.091478f
C2814 _081_ _178_/a_201_297# 0.046678f
C2815 counter\[10\] _052_ 0.022884f
C2816 _083_ _174_/a_79_21# 0.014098f
C2817 divider\[1\] _262_/a_109_93# 0.014229f
C2818 r2r_out[1] _322_/a_27_47# 0.042373f
C2819 _353_/a_193_47# VPWR 0.047103f
C2820 VPWR _056_ 0.587274f
C2821 _057_ _337_/a_891_413# 0.011971f
C2822 _025_ _349_/a_27_47# 0.064056f
C2823 _339_/a_27_47# VPWR 0.114784f
C2824 VPWR _113_ 0.529459f
C2825 _040_ _035_ 0.024824f
C2826 _357_/a_448_47# net12 0.016786f
C2827 _357_/a_1108_47# _000_ 0.025775f
C2828 VGND _340_/a_1062_300# 0.077733f
C2829 VGND _327_/a_27_47# 0.052063f
C2830 _094_ _117_ 0.050063f
C2831 _145_ _143_ 0.049754f
C2832 _149_ _002_ 0.023317f
C2833 _085_ clknet_2_3__leaf_clk 0.026545f
C2834 clknet_0_clk _059_ 0.021474f
C2835 _345_/a_193_47# _021_ 0.362608f
C2836 _145_ _141_ 0.088122f
C2837 _140_ _141_ 0.010183f
C2838 _290_/a_27_413# counter\[13\] 0.010177f
C2839 _275_/a_109_93# clknet_2_2__leaf_clk 0.011481f
C2840 VPWR _035_ 0.454672f
C2841 _328_/a_381_47# divider\[2\] 0.012219f
C2842 VGND _134_ 0.11488f
C2843 _240_/a_68_297# _059_ 0.086118f
C2844 VPWR hold10/a_285_47# 0.01885f
C2845 _089_ _184_/a_27_47# 0.010496f
C2846 _081_ _087_ 0.112738f
C2847 _356_/a_891_413# net3 0.01106f
C2848 VGND _354_/a_634_159# 0.016987f
C2849 clk n_rst 0.042648f
C2850 VGND net16 0.244538f
C2851 VPWR _150_ 0.031318f
C2852 _281_/a_27_47# _033_ 0.011897f
C2853 hold9/a_49_47# _335_/a_1062_300# 0.021055f
C2854 _092_ _016_ 0.027133f
C2855 VPWR _016_ 0.445566f
C2856 VPWR hold8/a_391_47# 0.010225f
C2857 _346_/a_1059_315# _066_ 0.07382f
C2858 VGND _026_ 0.104318f
C2859 clknet_0_clk counter\[0\] 0.014994f
C2860 r2r_out[3] _335_/a_1062_300# 0.022277f
C2861 _040_ _292_/a_85_193# 0.060708f
C2862 counter\[9\] _065_ 0.039262f
C2863 VPWR _017_ 0.087392f
C2864 _053_ _074_ 0.087811f
C2865 hold9/a_49_47# r2r_out[2] 0.050442f
C2866 divider\[0\] _260_/a_215_53# 0.065341f
C2867 counter\[10\] _066_ 0.510682f
C2868 r2r_out[3] r2r_out[2] 1.147631f
C2869 VGND _195_/a_227_47# -0.020173f
C2870 VPWR _292_/a_85_193# -0.013455f
C2871 net22 rst 0.216235f
C2872 VGND _125_ -0.012092f
C2873 _342_/a_27_47# _345_/a_27_47# 0.042702f
C2874 counter\[10\] _236_/a_27_47# 0.045569f
C2875 r2r_out[3] _065_ 0.067372f
C2876 clknet_2_2__leaf_clk _028_ 0.106868f
C2877 VPWR _245_/a_75_212# 0.029854f
C2878 _053_ r2r_out[5] 0.063848f
C2879 clknet_2_0__leaf_clk _117_ 0.1094f
C2880 _139_ _138_ 0.0175f
C2881 _321_/a_448_47# r2r_out[2] 0.046172f
C2882 _149_ _350_/a_1059_315# 0.013154f
C2883 VGND _325_/a_27_47# 0.035732f
C2884 _329_/a_27_47# clknet_2_2__leaf_clk 0.085842f
C2885 _159_ net9 0.019662f
C2886 _101_ _108_ 0.013409f
C2887 _097_ _100_ 0.054484f
C2888 counter\[2\] _019_ 0.277771f
C2889 _355_/a_27_47# VGND 0.031596f
C2890 VPWR _036_ 0.345543f
C2891 _035_ counter\[14\] 0.020292f
C2892 VPWR _206_/a_113_297# 0.072857f
C2893 counter\[13\] _035_ 0.33509f
C2894 _069_ r2r_out[0] 0.017771f
C2895 counter\[7\] _065_ 0.032081f
C2896 VGND _332_/a_193_47# 0.015128f
C2897 VPWR _332_/a_27_47# 0.082255f
C2898 _115_ _132_ 0.013848f
C2899 _346_/a_193_47# clknet_2_0__leaf_clk 0.01084f
C2900 net17 counter\[0\] 0.139329f
C2901 _348_/a_634_159# clknet_2_0__leaf_clk 0.01894f
C2902 _298_/a_103_199# _047_ 0.028657f
C2903 VGND _102_ 0.076056f
C2904 VPWR counter\[3\] 0.29987f
C2905 _027_ clknet_2_0__leaf_clk 0.11807f
C2906 hold7/a_391_47# net1 0.069056f
C2907 net22 _092_ 0.098228f
C2908 _046_ _041_ 0.083315f
C2909 net1 _029_ 0.05269f
C2910 net10 _268_/a_215_53# 0.063277f
C2911 _040_ _043_ 0.074481f
C2912 net22 VPWR 0.254504f
C2913 _059_ _078_ 0.319121f
C2914 net5 net10 0.530572f
C2915 VGND divider\[3\] 0.183326f
C2916 _144_ counter\[9\] 0.207774f
C2917 r2r_out[6] net7 0.072947f
C2918 VPWR _043_ 0.183111f
C2919 _336_/a_193_47# clknet_2_3__leaf_clk 0.012641f
C2920 _135_ counter\[8\] 0.012093f
C2921 VPWR clkbuf_2_1__f_clk/a_110_47# 0.138727f
C2922 _149_ rst 0.071679f
C2923 _055_ _054_ 0.223497f
C2924 _267_/a_298_297# VPWR -0.015264f
C2925 _027_ _130_ 0.026554f
C2926 _112_ VGND 0.32836f
C2927 _053_ net4 0.02457f
C2928 VPWR hold4/a_391_47# -0.010683f
C2929 _048_ clkbuf_2_2__f_clk/a_110_47# 0.043015f
C2930 _132_ counter\[8\] 0.04734f
C2931 divider\[4\] _329_/a_466_413# 0.023332f
C2932 counter\[0\] _078_ 0.314145f
C2933 _219_/a_227_47# _078_ 0.014696f
C2934 _079_ clknet_2_3__leaf_clk 0.024741f
C2935 _149_ _259_/a_27_47# 0.014531f
C2936 _065_ _350_/a_1059_315# 0.018528f
C2937 _176_/a_68_297# _087_ 0.078411f
C2938 VGND counter\[15\] 1.158037f
C2939 VPWR divider\[7\] 1.02765f
C2940 divider\[1\] net3 0.106235f
C2941 _136_ _223_/a_250_297# 0.089695f
C2942 _161_ counter\[8\] 0.053097f
C2943 _356_/a_27_47# _356_/a_466_413# -0.013083f
C2944 divider\[3\] counter\[15\] 0.350004f
C2945 _334_/a_27_47# VPWR 0.110275f
C2946 _082_ r2r_out[4] 0.043817f
C2947 _054_ counter\[8\] 0.105471f
C2948 _273_/a_215_53# rst 0.011459f
C2949 _053_ _335_/a_475_413# 0.021961f
C2950 _057_ _009_ 0.123908f
C2951 counter\[0\] _061_ 0.061963f
C2952 _339_/a_193_47# _057_ 0.035735f
C2953 _065_ _354_/a_466_413# 0.022139f
C2954 _057_ _340_/a_1062_300# 0.040765f
C2955 _036_ counter\[13\] 0.278358f
C2956 counter\[1\] net17 0.041218f
C2957 _071_ clk 0.022091f
C2958 VGND _052_ 0.763969f
C2959 _031_ net1 0.081699f
C2960 VPWR _178_/a_75_199# 0.048948f
C2961 divider\[6\] net8 0.060209f
C2962 divider\[6\] _008_ 0.081079f
C2963 net3 net20 0.080157f
C2964 _342_/a_381_47# _018_ 0.023443f
C2965 _111_ VGND 0.324754f
C2966 _149_ VPWR 6.826027f
C2967 _060_ _341_/a_891_413# 0.048608f
C2968 clknet_2_0__leaf_clk _350_/a_27_47# 0.118473f
C2969 clk _319_/a_29_53# 0.06088f
C2970 _148_ _004_ 0.235648f
C2971 _294_/a_215_47# _041_ 0.032291f
C2972 _355_/a_634_159# net4 0.038837f
C2973 _233_/a_80_21# _129_ 0.090841f
C2974 net7 _007_ 0.041913f
C2975 _124_ _078_ 0.16126f
C2976 VPWR _271_/a_29_53# 0.041109f
C2977 _126_ _065_ 0.03553f
C2978 _112_ _052_ 0.092619f
C2979 _065_ rst 0.056768f
C2980 _043_ counter\[13\] 0.142403f
C2981 _065_ _030_ 0.136442f
C2982 hold7/a_49_47# _341_/a_193_47# 0.012378f
C2983 _173_/a_27_47# _077_ 0.079781f
C2984 VGND _087_ 0.018438f
C2985 _355_/a_27_47# _066_ 0.039234f
C2986 divider\[4\] divider\[2\] 0.053145f
C2987 _060_ _063_ 0.09748f
C2988 _101_ counter\[0\] 0.098814f
C2989 counter\[1\] _078_ 0.026778f
C2990 _060_ clk 0.024568f
C2991 _224_/a_59_75# _121_ 0.015235f
C2992 r2r_out[7] rst 0.336104f
C2993 VGND _075_ 0.093016f
C2994 divider\[1\] _281_/a_27_47# 0.015351f
C2995 divider\[7\] counter\[14\] 0.037029f
C2996 data[5] net9 0.034576f
C2997 net4 net8 0.01976f
C2998 divider\[6\] _049_ 0.134094f
C2999 VGND _066_ 3.263349f
C3000 _343_/a_193_47# hold5/a_49_47# 0.01236f
C3001 VPWR _335_/a_1062_300# 0.027719f
C3002 counter\[10\] counter\[9\] 0.419442f
C3003 net6 _077_ 0.195035f
C3004 VGND r2r_out[0] 3.560599f
C3005 input7/a_27_47# net9 0.046409f
C3006 _040_ _041_ 0.199323f
C3007 VPWR hold3/a_285_47# 0.029014f
C3008 VGND hold3/a_391_47# 0.019113f
C3009 _311_/a_27_297# _054_ 0.069673f
C3010 _356_/a_193_47# _147_ 0.010611f
C3011 _313_/a_27_47# clknet_2_1__leaf_clk 0.017542f
C3012 _111_ _052_ 0.011351f
C3013 _236_/a_27_47# VGND 0.037749f
C3014 VPWR r2r_out[2] 0.879402f
C3015 _329_/a_1059_315# net10 0.062272f
C3016 _079_ net9 0.016141f
C3017 VGND _333_/a_1062_300# 0.075479f
C3018 VPWR _333_/a_475_413# 0.01025f
C3019 clknet_2_3__leaf_clk counter\[8\] 0.033499f
C3020 VPWR _041_ 0.18175f
C3021 divider\[1\] divider\[2\] 0.02996f
C3022 VGND _022_ 0.224246f
C3023 VPWR _065_ 5.447734f
C3024 _149_ _114_ 0.022135f
C3025 VGND _341_/a_634_159# 0.034241f
C3026 _243_/a_93_21# counter\[8\] 0.011271f
C3027 _329_/a_634_159# clknet_2_2__leaf_clk 0.03905f
C3028 _171_/a_27_47# _065_ 0.018096f
C3029 divider\[2\] _327_/a_1059_315# 0.060288f
C3030 _094_ hold4/a_49_47# 0.079546f
C3031 clkbuf_2_2__f_clk/a_110_47# net9 0.097327f
C3032 _155_ divider\[5\] 0.086212f
C3033 _092_ r2r_out[7] 0.066225f
C3034 _103_ _019_ 0.076393f
C3035 _066_ counter\[15\] 0.040376f
C3036 _053_ r2r_out[4] 0.044737f
C3037 VPWR r2r_out[7] 0.990398f
C3038 _253_/a_79_21# VPWR 0.016017f
C3039 VGND _347_/a_634_159# 0.017434f
C3040 VPWR _347_/a_193_47# 0.045404f
C3041 _072_ _012_ 0.028148f
C3042 VGND _057_ 2.710989f
C3043 _343_/a_193_47# counter\[2\] 0.168759f
C3044 _141_ _248_/a_227_47# 0.017365f
C3045 counter\[1\] _101_ 0.070629f
C3046 VGND clkbuf_0_clk/a_110_47# 0.032312f
C3047 VGND _221_/a_68_297# 0.048607f
C3048 net6 net4 0.021737f
C3049 _148_ net3 0.284279f
C3050 _157_ net9 0.022444f
C3051 _345_/a_1059_315# hold2/a_49_47# 0.013516f
C3052 _353_/a_891_413# _078_ 0.038529f
C3053 _004_ _328_/a_27_47# 0.052335f
C3054 input2/a_27_47# data[1] 0.016927f
C3055 _294_/a_78_199# _041_ 0.015333f
C3056 _066_ _052_ 0.022861f
C3057 r2r_out[3] _069_ 0.014694f
C3058 _066_ _163_/a_193_297# 0.02868f
C3059 _097_ _197_/a_27_47# 0.010981f
C3060 _072_ _011_ 0.01613f
C3061 _089_ net7 0.027111f
C3062 net1 _341_/a_891_413# 0.011946f
C3063 _111_ _066_ 0.079117f
C3064 _146_ net1 0.044022f
C3065 _057_ counter\[15\] 0.227116f
C3066 _326_/a_634_159# _002_ 0.029611f
C3067 _149_ _106_ 0.061572f
C3068 divider\[4\] _042_ 0.028078f
C3069 clkbuf_2_2__f_clk/a_110_47# clknet_2_2__leaf_clk 0.021304f
C3070 counter\[5\] _109_ 0.085029f
C3071 r2r_out[1] _317_/a_113_297# 0.03239f
C3072 net5 _280_/a_207_413# 0.013028f
C3073 _114_ _065_ 0.023842f
C3074 _048_ _142_ 0.150153f
C3075 _340_/a_27_47# clknet_2_3__leaf_clk 0.030688f
C3076 VPWR hold1/a_391_47# 0.018268f
C3077 counter\[14\] _041_ 0.028831f
C3078 _336_/a_891_413# VPWR 0.022151f
C3079 _152_ net10 0.048917f
C3080 _105_ counter\[5\] 0.031614f
C3081 counter\[13\] _041_ 0.022625f
C3082 _063_ net1 0.037773f
C3083 _144_ VPWR 0.314935f
C3084 clk net1 0.036028f
C3085 _330_/a_381_47# _006_ 0.022668f
C3086 _348_/a_891_413# _350_/a_1059_315# 0.010655f
C3087 hold5/a_49_47# clkbuf_2_1__f_clk/a_110_47# 0.018665f
C3088 _253_/a_79_21# counter\[14\] 0.03261f
C3089 VGND _013_ 0.041176f
C3090 _274_/a_27_413# VGND 0.017822f
C3091 _053_ _064_ 0.222537f
C3092 VGND _276_/a_215_297# 0.046157f
C3093 VPWR _276_/a_27_413# 0.04515f
C3094 _084_ _091_ 0.041078f
C3095 net7 _262_/a_215_53# 0.052009f
C3096 net9 counter\[8\] 0.017802f
C3097 _078_ _029_ 0.031812f
C3098 VPWR _177_/a_59_75# 0.030642f
C3099 net9 _143_ 0.020043f
C3100 _141_ net9 0.195959f
C3101 counter\[2\] counter\[3\] 0.045702f
C3102 _236_/a_27_47# _066_ 0.070092f
C3103 _125_ counter\[9\] 0.09202f
C3104 net6 _329_/a_891_413# 0.016556f
C3105 _094_ _344_/a_381_47# 0.016837f
C3106 _057_ _087_ 0.016339f
C3107 _333_/a_1062_300# r2r_out[0] 0.036475f
C3108 _308_/a_27_47# _054_ 0.132611f
C3109 _149_ _023_ 0.172133f
C3110 counter\[5\] _211_/a_27_47# 0.034525f
C3111 _057_ _075_ 0.041446f
C3112 _070_ _071_ 0.225403f
C3113 _173_/a_27_47# r2r_out[4] 0.029345f
C3114 VPWR input10/a_27_47# 0.097799f
C3115 _065_ _106_ 0.030023f
C3116 _053_ _321_/a_222_93# 0.016855f
C3117 VPWR data[3] 0.228412f
C3118 _033_ net5 0.021308f
C3119 _121_ counter\[8\] 0.36872f
C3120 _328_/a_193_47# _328_/a_634_159# -0.016573f
C3121 _328_/a_27_47# _328_/a_466_413# -0.013083f
C3122 VPWR _038_ 0.613658f
C3123 _148_ divider\[2\] 0.040456f
C3124 _356_/a_634_159# VGND 0.017302f
C3125 counter\[10\] _126_ 0.47129f
C3126 _070_ _319_/a_29_53# 0.014929f
C3127 _159_ _133_ 0.02255f
C3128 _066_ _057_ 1.884603f
C3129 _097_ hold4/a_49_47# 0.029815f
C3130 counter\[0\] hold4/a_285_47# 0.048157f
C3131 _057_ _335_/a_891_413# 0.011419f
C3132 counter\[0\] _095_ 0.07247f
C3133 _057_ r2r_out[0] 0.061563f
C3134 _265_/a_215_297# net5 0.043167f
C3135 _066_ clkbuf_0_clk/a_110_47# 0.039172f
C3136 VPWR _342_/a_466_413# 0.026548f
C3137 VGND _342_/a_1059_315# 0.012059f
C3138 _144_ counter\[14\] 0.218533f
C3139 _005_ rst 0.020822f
C3140 VPWR _119_ 0.220112f
C3141 _291_/a_27_47# _289_/a_76_199# 0.017347f
C3142 _334_/a_27_47# counter\[2\] 0.010583f
C3143 _053_ _320_/a_209_297# 0.044855f
C3144 net6 r2r_out[4] 0.034103f
C3145 _154_ clknet_2_2__leaf_clk 0.086761f
C3146 _227_/a_59_75# _132_ 0.016226f
C3147 VGND counter\[9\] 1.504232f
C3148 clknet_0_clk _094_ 0.034953f
C3149 _356_/a_634_159# counter\[15\] 0.017132f
C3150 VGND clkbuf_2_3__f_clk/a_110_47# 0.159557f
C3151 _213_/a_215_53# _117_ 0.059235f
C3152 _213_/a_109_93# _115_ 0.041994f
C3153 VGND hold9/a_49_47# 0.034261f
C3154 counter\[1\] _190_/a_76_199# 0.029224f
C3155 _311_/a_27_297# net2 0.07279f
C3156 VPWR _289_/a_226_47# 0.011073f
C3157 r2r_out[3] VGND 1.251787f
C3158 _073_ _054_ 0.045268f
C3159 _346_/a_1059_315# VPWR 0.033781f
C3160 _346_/a_891_413# VGND 0.020233f
C3161 _348_/a_891_413# VPWR -0.010084f
C3162 _053_ _056_ 0.564449f
C3163 hold6/a_391_47# net18 0.024845f
C3164 _339_/a_27_47# _015_ 0.027735f
C3165 VPWR _081_ 0.744663f
C3166 _053_ _339_/a_27_47# 0.05025f
C3167 _335_/a_27_47# clknet_2_1__leaf_clk 0.02079f
C3168 _057_ clkbuf_0_clk/a_110_47# 0.020497f
C3169 _057_ _221_/a_68_297# 0.014589f
C3170 r2r_out[3] _324_/a_68_297# 0.013137f
C3171 counter\[10\] VPWR 0.552701f
C3172 _142_ net9 0.030994f
C3173 divider\[6\] _331_/a_27_47# 0.344645f
C3174 _053_ _340_/a_475_413# 0.023224f
C3175 _081_ _171_/a_27_47# 0.012211f
C3176 VGND _248_/a_77_199# 0.015267f
C3177 counter\[15\] counter\[9\] 0.262006f
C3178 r2r_out[6] _085_ 0.267581f
C3179 VGND _002_ 0.055685f
C3180 VPWR _005_ 0.260075f
C3181 _053_ hold10/a_285_47# 0.019812f
C3182 _353_/a_27_47# _029_ 0.033289f
C3183 _347_/a_193_47# _023_ 0.409771f
C3184 _066_ _013_ 0.063211f
C3185 counter\[1\] hold4/a_285_47# 0.029704f
C3186 counter\[1\] _095_ 0.202979f
C3187 VGND _137_ 0.123828f
C3188 counter\[7\] VGND 0.590636f
C3189 VPWR _093_ 0.251394f
C3190 _114_ _119_ 0.032603f
C3191 _044_ _042_ 0.455349f
C3192 VGND _147_ 0.020772f
C3193 clknet_0_clk clknet_2_0__leaf_clk 0.02222f
C3194 _053_ _016_ 0.071626f
C3195 hold10/a_391_47# rst 0.076093f
C3196 _052_ counter\[9\] 0.05447f
C3197 _326_/a_634_159# VPWR 0.021698f
C3198 _326_/a_466_413# VGND 0.018779f
C3199 counter\[4\] _108_ 0.131518f
C3200 _328_/a_27_47# divider\[2\] 0.039288f
C3201 counter\[12\] _045_ 0.019919f
C3202 _054_ net3 0.230388f
C3203 VGND _046_ 0.395257f
C3204 VPWR _069_ 0.260442f
C3205 _336_/a_475_413# clk 0.023736f
C3206 net11 clk 0.016847f
C3207 _265_/a_298_297# net3 0.013686f
C3208 _010_ _064_ 0.012162f
C3209 r2r_out[1] _055_ 0.165876f
C3210 _142_ clknet_2_2__leaf_clk 0.023349f
C3211 _112_ counter\[7\] 0.222008f
C3212 _336_/a_27_47# _336_/a_193_47# -0.10052f
C3213 _291_/a_27_47# _035_ 0.035489f
C3214 _057_ _013_ 0.073179f
C3215 _155_ _159_ 0.082982f
C3216 counter\[2\] _065_ 0.096136f
C3217 counter\[0\] _341_/a_27_47# 0.04829f
C3218 _251_/a_27_47# _144_ 0.041572f
C3219 _353_/a_634_159# VPWR 0.016978f
C3220 _060_ _091_ 0.207479f
C3221 VPWR _009_ 0.401003f
C3222 _195_/a_77_199# _098_ 0.0473f
C3223 counter\[6\] counter\[5\] 0.846831f
C3224 _057_ _337_/a_381_47# 0.014583f
C3225 _025_ _349_/a_193_47# 0.224369f
C3226 _339_/a_193_47# VPWR 0.043304f
C3227 _125_ _126_ 0.050148f
C3228 VPWR _327_/a_27_47# -0.02559f
C3229 VGND _327_/a_193_47# -0.079822f
C3230 VPWR _340_/a_1062_300# 0.052194f
C3231 VGND _340_/a_891_413# 0.022385f
C3232 VGND _350_/a_1059_315# 0.052346f
C3233 _094_ _078_ 0.898834f
C3234 VPWR _350_/a_466_413# 0.012181f
C3235 _234_/a_113_297# _130_ 0.018132f
C3236 divider\[4\] _268_/a_215_53# 0.061808f
C3237 divider\[4\] net5 0.042287f
C3238 _345_/a_634_159# _021_ 0.053148f
C3239 _094_ _051_ 0.493109f
C3240 _073_ clknet_2_3__leaf_clk 0.31493f
C3241 _183_/a_59_75# _091_ 0.012903f
C3242 counter\[7\] _052_ 0.202689f
C3243 _237_/a_27_47# _132_ 0.031342f
C3244 VPWR _279_/a_27_413# 0.053182f
C3245 VPWR _134_ 0.130426f
C3246 VPWR hold10/a_391_47# 0.012889f
C3247 _343_/a_466_413# VGND 0.010682f
C3248 r2r_out[3] _075_ 0.074045f
C3249 _066_ counter\[9\] 0.079839f
C3250 _103_ counter\[3\] 0.31045f
C3251 _120_ _054_ 0.055363f
C3252 VGND _357_/a_193_47# 0.026641f
C3253 VPWR _357_/a_27_47# 0.060119f
C3254 _153_ divider\[2\] 0.040488f
C3255 _352_/a_27_47# counter\[11\] 0.423881f
C3256 _281_/a_27_47# _161_ 0.034903f
C3257 _098_ _099_ 0.068565f
C3258 _236_/a_27_47# counter\[9\] 0.029834f
C3259 _053_ net22 0.052556f
C3260 _326_/a_1059_315# _149_ 0.012281f
C3261 _346_/a_891_413# _066_ 0.024665f
C3262 VPWR _026_ 0.340731f
C3263 clkbuf_2_0__f_clk/a_110_47# _115_ 0.023295f
C3264 r2r_out[3] r2r_out[0] 0.264457f
C3265 _261_/a_27_413# net1 0.026366f
C3266 hold9/a_285_47# r2r_out[2] 0.071113f
C3267 divider\[1\] net1 0.02421f
C3268 divider\[0\] _260_/a_109_93# 0.05359f
C3269 _337_/a_27_47# _337_/a_193_47# -0.036505f
C3270 VPWR _176_/a_68_297# 0.012972f
C3271 _053_ clkbuf_2_1__f_clk/a_110_47# 0.015175f
C3272 divider\[1\] net5 0.023597f
C3273 VGND _294_/a_215_47# -0.018669f
C3274 _063_ _078_ 0.015829f
C3275 _256_/a_81_21# clknet_2_3__leaf_clk 0.010667f
C3276 _078_ clk 0.080636f
C3277 VGND _126_ 0.606044f
C3278 VPWR _125_ 0.402364f
C3279 VGND rst 4.293119f
C3280 VGND _030_ 0.048136f
C3281 VGND hold7/a_49_47# 0.030587f
C3282 _346_/a_381_47# _065_ 0.015201f
C3283 divider\[3\] rst 0.018948f
C3284 _011_ _335_/a_27_47# 0.027735f
C3285 net3 clknet_2_3__leaf_clk 0.201254f
C3286 clknet_2_0__leaf_clk _078_ 0.0584f
C3287 _160_ _159_ 0.027089f
C3288 _101_ _212_/a_80_21# 0.081633f
C3289 _318_/a_27_47# r2r_out[2] 0.033089f
C3290 _063_ _061_ 0.063495f
C3291 _010_ _056_ 0.097581f
C3292 VGND _259_/a_27_47# 0.031582f
C3293 _094_ _101_ 0.139418f
C3294 counter\[7\] _066_ 0.023505f
C3295 _149_ _350_/a_891_413# 0.017158f
C3296 VPWR _325_/a_27_47# -0.127956f
C3297 VGND _325_/a_193_47# -0.115211f
C3298 net20 net1 0.014245f
C3299 _149_ _187_/a_79_21# 0.01701f
C3300 r2r_out[3] _057_ 0.263612f
C3301 _329_/a_193_47# clknet_2_2__leaf_clk 0.255965f
C3302 _094_ hold6/a_391_47# 0.01808f
C3303 VGND _241_/a_59_75# 0.07969f
C3304 counter\[0\] _019_ 0.040199f
C3305 r2r_out[1] _311_/a_27_297# 0.029982f
C3306 input11/a_75_212# n_rst 0.020948f
C3307 _355_/a_193_47# VGND -0.121544f
C3308 _355_/a_27_47# VPWR 0.099331f
C3309 _291_/a_27_47# _043_ 0.11786f
C3310 counter\[15\] rst 0.182766f
C3311 VPWR _332_/a_193_47# 0.032803f
C3312 _117_ _132_ 0.121349f
C3313 _115_ _133_ 0.023419f
C3314 _040_ VGND 0.174084f
C3315 _096_ clknet_2_1__leaf_clk 0.037565f
C3316 _348_/a_466_413# clknet_2_0__leaf_clk 0.039904f
C3317 _048_ _297_/a_215_47# 0.049945f
C3318 _104_ counter\[3\] 0.304222f
C3319 VPWR _102_ 0.124891f
C3320 VGND _107_ 0.252189f
C3321 net4 _327_/a_466_413# 0.016673f
C3322 _053_ _149_ 0.198582f
C3323 divider\[6\] net10 0.323889f
C3324 input1/a_27_47# data[0] 0.0509f
C3325 _053_ _179_/a_215_47# 0.011125f
C3326 net10 _268_/a_109_93# 0.013389f
C3327 divider\[4\] _328_/a_1059_315# 0.021487f
C3328 _092_ VGND 0.220709f
C3329 VGND VPWR 20.264658f
C3330 net14 VGND 0.038652f
C3331 _332_/a_27_47# _008_ 0.079133f
C3332 VPWR divider\[3\] 0.727567f
C3333 _057_ _137_ 0.024352f
C3334 input5/a_27_47# VGND 0.060285f
C3335 clkbuf_2_0__f_clk/a_110_47# hold6/a_49_47# 0.017057f
C3336 VGND _171_/a_27_47# 0.064617f
C3337 VPWR _324_/a_68_297# 0.033721f
C3338 r2r_out[6] _086_ 0.096516f
C3339 VGND _014_ 0.239186f
C3340 _057_ _147_ 0.162595f
C3341 _004_ clknet_2_2__leaf_clk 0.211486f
C3342 _336_/a_193_47# _012_ 0.060567f
C3343 _336_/a_891_413# hold9/a_285_47# 0.014357f
C3344 _024_ clknet_2_0__leaf_clk 0.153085f
C3345 _112_ VPWR 0.459019f
C3346 _320_/a_80_21# clk 0.072207f
C3347 VGND _080_ 0.048767f
C3348 _133_ counter\[8\] 0.06714f
C3349 divider\[4\] _329_/a_1059_315# 0.024545f
C3350 _097_ _078_ 0.018275f
C3351 _219_/a_227_47# _118_ 0.075193f
C3352 _227_/a_59_75# _121_ 0.066981f
C3353 VPWR counter\[15\] 4.440105f
C3354 _157_ _331_/a_466_413# 0.018883f
C3355 _133_ _141_ 0.022331f
C3356 _334_/a_193_47# VPWR 0.037698f
C3357 _188_/a_27_47# VGND 0.076307f
C3358 _343_/a_1059_315# _065_ 0.016274f
C3359 _037_ VPWR 0.268888f
C3360 _339_/a_634_183# _057_ 0.018086f
C3361 net2 net3 0.029262f
C3362 _057_ _340_/a_891_413# 0.012739f
C3363 net3 net9 0.017623f
C3364 _053_ r2r_out[2] 0.114278f
C3365 _053_ _333_/a_475_413# 0.037695f
C3366 VPWR _052_ 0.473837f
C3367 _284_/a_27_413# divider\[6\] 0.010358f
C3368 VPWR _178_/a_201_297# -0.017899f
C3369 _053_ _065_ 0.212103f
C3370 _066_ _126_ 0.026148f
C3371 _314_/a_113_297# _061_ 0.021844f
C3372 VPWR _163_/a_193_297# -0.013693f
C3373 _148_ net1 0.555669f
C3374 VGND _116_ 0.479218f
C3375 _111_ VPWR 0.527024f
C3376 _114_ VGND 0.036805f
C3377 _060_ _341_/a_381_47# 0.017894f
C3378 clknet_2_0__leaf_clk _350_/a_193_47# 0.177359f
C3379 net7 _154_ 0.033172f
C3380 VGND counter\[14\] 1.510656f
C3381 _148_ net5 0.94963f
C3382 input8/a_27_47# VGND 0.058673f
C3383 VGND _330_/a_27_47# 0.050677f
C3384 VGND counter\[13\] 1.288893f
C3385 _351_/a_27_47# _027_ 0.107209f
C3386 _053_ r2r_out[7] 0.079688f
C3387 _355_/a_466_413# net4 0.017723f
C3388 _292_/a_516_297# _041_ 0.02293f
C3389 counter\[1\] _189_/a_285_47# 0.03219f
C3390 _149_ net8 0.026088f
C3391 hold7/a_285_47# _341_/a_193_47# 0.011561f
C3392 hold7/a_391_47# _341_/a_27_47# 0.011338f
C3393 _173_/a_109_297# _077_ 0.011215f
C3394 _338_/a_27_47# r2r_out[5] 0.483418f
C3395 divider\[2\] _264_/a_109_93# 0.013226f
C3396 _039_ _038_ 0.131938f
C3397 _112_ _116_ 0.155106f
C3398 counter\[10\] _233_/a_80_21# 0.11794f
C3399 VPWR _087_ 0.356621f
C3400 _355_/a_193_47# _066_ 0.02281f
C3401 _101_ _097_ 0.150649f
C3402 VPWR _075_ 0.404691f
C3403 _186_/a_113_297# _078_ 0.012045f
C3404 _348_/a_27_47# _348_/a_193_47# -0.012897f
C3405 _188_/a_27_47# _052_ 0.030073f
C3406 clknet_0_clk net20 0.025851f
C3407 _291_/a_27_47# _041_ 0.04558f
C3408 _057_ rst 0.014411f
C3409 counter\[15\] counter\[14\] 0.35758f
C3410 _260_/a_215_53# net3 0.021752f
C3411 _094_ counter\[11\] 0.047882f
C3412 _066_ _107_ 0.360637f
C3413 _031_ net4 0.196077f
C3414 _094_ _190_/a_76_199# 0.09095f
C3415 _308_/a_27_47# _139_ 0.010501f
C3416 _334_/a_27_47# _010_ 0.087146f
C3417 VPWR _066_ 5.55827f
C3418 _343_/a_193_47# hold5/a_285_47# 0.011479f
C3419 input2/a_27_47# net1 0.041167f
C3420 net14 _066_ 0.089224f
C3421 _037_ counter\[14\] 0.10395f
C3422 VPWR r2r_out[0] 2.531981f
C3423 net11 _357_/a_1283_21# 0.103018f
C3424 r2r_out[3] hold9/a_49_47# 0.068265f
C3425 VPWR hold3/a_391_47# 0.015471f
C3426 VGND _106_ 0.143612f
C3427 _114_ _052_ 0.014389f
C3428 net6 _178_/a_75_199# 0.010326f
C3429 _329_/a_891_413# net10 0.039071f
C3430 _036_ _280_/a_27_413# 0.057329f
C3431 _065_ _190_/a_489_47# 0.045409f
C3432 VGND _333_/a_891_413# 0.022519f
C3433 VPWR _333_/a_1062_300# 0.075233f
C3434 _065_ _104_ 0.314801f
C3435 VPWR _022_ 0.093647f
C3436 _149_ net6 0.024592f
C3437 VGND _341_/a_466_413# 0.041184f
C3438 _111_ _114_ 0.187821f
C3439 _120_ _121_ 0.474522f
C3440 _081_ _082_ 0.093031f
C3441 _329_/a_466_413# clknet_2_2__leaf_clk 0.021921f
C3442 _151_ net3 0.201677f
C3443 _066_ _080_ 0.244024f
C3444 divider\[2\] _327_/a_891_413# 0.047071f
C3445 _094_ hold4/a_285_47# 0.094453f
C3446 _131_ _078_ 0.016318f
C3447 _355_/a_193_47# clkbuf_0_clk/a_110_47# 0.013208f
C3448 _070_ _078_ 0.031969f
C3449 _094_ _095_ 0.106922f
C3450 clknet_2_1__leaf_clk _195_/a_77_199# 0.015751f
C3451 counter\[7\] counter\[9\] 0.111655f
C3452 hold8/a_49_47# _054_ 0.040396f
C3453 _131_ _051_ 0.156165f
C3454 _060_ _054_ 0.560197f
C3455 _253_/a_215_47# VGND -0.017416f
C3456 VGND _347_/a_466_413# 0.020077f
C3457 VPWR _347_/a_634_159# 0.018065f
C3458 hold5/a_49_47# _195_/a_227_47# 0.029857f
C3459 _159_ _283_/a_78_199# 0.020927f
C3460 _003_ _327_/a_27_47# 0.028922f
C3461 _152_ _327_/a_1059_315# 0.022348f
C3462 VPWR _057_ 3.414756f
C3463 VGND _122_ 0.200719f
C3464 _343_/a_634_159# counter\[2\] 0.038223f
C3465 clkbuf_2_3__f_clk/a_110_47# _147_ 0.02408f
C3466 net10 data[6] 0.300281f
C3467 VPWR clkbuf_0_clk/a_110_47# 0.230388f
C3468 VPWR _221_/a_68_297# 0.016887f
C3469 counter\[2\] net16 0.201782f
C3470 _353_/a_381_47# _078_ 0.016597f
C3471 _004_ _328_/a_193_47# 0.079151f
C3472 _074_ clk 0.135815f
C3473 _138_ counter\[8\] 0.01262f
C3474 _251_/a_27_47# VGND 0.033341f
C3475 net2 _084_ 0.011758f
C3476 _084_ net9 0.037624f
C3477 _114_ _066_ 0.030787f
C3478 VGND _023_ 0.195975f
C3479 _066_ counter\[14\] 0.086357f
C3480 r2r_out[5] clk 0.29032f
C3481 _326_/a_466_413# _002_ 0.030904f
C3482 net17 _193_/a_113_297# 0.104964f
C3483 _149_ _108_ 0.073789f
C3484 _356_/a_1059_315# hold8/a_391_47# 0.015536f
C3485 divider\[2\] clknet_2_2__leaf_clk 0.228032f
C3486 r2r_out[1] _333_/a_27_47# 0.449199f
C3487 _340_/a_193_47# clknet_2_3__leaf_clk 0.016978f
C3488 VGND hold5/a_49_47# -0.017056f
C3489 counter\[12\] _041_ 0.014031f
C3490 _010_ _065_ 0.434106f
C3491 data[0] net12 0.064401f
C3492 _160_ counter\[8\] 0.157151f
C3493 _149_ _347_/a_1059_315# 0.055527f
C3494 _006_ _156_ 0.015616f
C3495 _136_ _054_ 0.294467f
C3496 _320_/a_80_21# _070_ 0.032984f
C3497 _121_ _117_ 0.493656f
C3498 VPWR _013_ 0.463192f
C3499 _274_/a_27_413# VPWR 0.028114f
C3500 _057_ counter\[14\] 0.09819f
C3501 net7 _262_/a_109_93# 0.043066f
C3502 _065_ _344_/a_27_47# 0.036575f
C3503 _125_ _228_/a_27_47# 0.11833f
C3504 counter\[5\] _216_/a_59_75# 0.025341f
C3505 counter\[0\] counter\[3\] 0.222218f
C3506 _060_ clknet_2_3__leaf_clk 0.501311f
C3507 _066_ _106_ 0.128945f
C3508 net18 _118_ 0.095735f
C3509 VGND counter\[2\] 1.464005f
C3510 _269_/a_27_413# rst 0.017024f
C3511 _187_/a_79_21# _093_ 0.021759f
C3512 clknet_0_clk _145_ 0.028186f
C3513 _003_ VGND 0.081134f
C3514 _065_ _108_ 0.090003f
C3515 counter\[0\] clkbuf_2_1__f_clk/a_110_47# 0.053135f
C3516 _161_ net5 0.057463f
C3517 _054_ net1 0.356094f
C3518 _356_/a_466_413# VGND 0.022292f
C3519 _054_ net5 0.053009f
C3520 _224_/a_59_75# _349_/a_1059_315# 0.014902f
C3521 VGND _233_/a_80_21# 0.046942f
C3522 counter\[0\] hold4/a_391_47# 0.054068f
C3523 _097_ hold4/a_285_47# 0.023984f
C3524 _053_ _093_ 0.051197f
C3525 _152_ _148_ 0.164636f
C3526 _278_/a_219_297# divider\[1\] 0.017631f
C3527 VPWR _342_/a_1059_315# 0.041376f
C3528 _144_ counter\[12\] 0.237567f
C3529 _238_/a_227_47# _035_ 0.01447f
C3530 _167_/a_27_47# VGND 0.029018f
C3531 _053_ _069_ 0.270794f
C3532 _258_/a_27_47# data[6] 0.012002f
C3533 VPWR counter\[9\] 1.888922f
C3534 _071_ net2 0.017982f
C3535 _073_ _337_/a_27_47# 0.01339f
C3536 VGND _269_/a_215_297# -0.017442f
C3537 VPWR _269_/a_27_413# 0.033116f
C3538 _023_ _066_ 0.028048f
C3539 _356_/a_466_413# counter\[15\] 0.031814f
C3540 VPWR clkbuf_2_3__f_clk/a_110_47# 0.112015f
C3541 counter\[1\] counter\[3\] 0.031192f
C3542 _213_/a_109_93# _117_ 0.01755f
C3543 VPWR hold9/a_49_47# 0.048993f
C3544 counter\[1\] _190_/a_206_369# 0.02925f
C3545 net4 _033_ 0.1435f
C3546 _311_/a_109_297# net2 0.024448f
C3547 _154_ _329_/a_27_47# 0.085562f
C3548 r2r_out[3] VPWR 1.592986f
C3549 VPWR _289_/a_489_413# 0.034027f
C3550 _149_ counter\[0\] 0.032993f
C3551 _319_/a_29_53# net9 0.025937f
C3552 _346_/a_891_413# VPWR 0.026337f
C3553 _053_ _009_ 0.141157f
C3554 _339_/a_193_47# _015_ 0.065484f
C3555 _136_ _243_/a_93_21# 0.023294f
C3556 _053_ _339_/a_193_47# 0.048858f
C3557 VGND _082_ 0.346132f
C3558 divider\[6\] _331_/a_193_47# 0.065414f
C3559 _347_/a_27_47# clknet_2_0__leaf_clk 0.112119f
C3560 _039_ VGND 0.473746f
C3561 VPWR _248_/a_77_199# 0.017263f
C3562 clknet_2_1__leaf_clk _333_/a_27_47# 0.022252f
C3563 VGND _318_/a_27_47# 0.032298f
C3564 VPWR _002_ 0.102178f
C3565 _049_ _038_ 0.310812f
C3566 _187_/a_297_47# net19 0.011336f
C3567 _065_ _128_ 0.03682f
C3568 _053_ hold10/a_391_47# 0.036088f
C3569 _353_/a_193_47# _029_ 0.23795f
C3570 _347_/a_634_159# _023_ 0.048438f
C3571 net2 _060_ 0.025124f
C3572 _251_/a_27_47# clkbuf_0_clk/a_110_47# 0.010123f
C3573 counter\[1\] hold4/a_391_47# 0.052169f
C3574 _060_ net9 0.904494f
C3575 net16 _103_ 0.18985f
C3576 hold5/a_285_47# _065_ 0.020006f
C3577 _212_/a_80_21# counter\[4\] 0.043944f
C3578 rst _340_/a_891_413# 0.013717f
C3579 _057_ _169_/a_149_47# 0.030537f
C3580 counter\[7\] VPWR 1.267232f
C3581 _094_ counter\[4\] 0.491041f
C3582 _040_ _046_ 0.064352f
C3583 _131_ counter\[11\] 0.143496f
C3584 counter\[15\] _255_/a_80_21# 0.013769f
C3585 clknet_2_3__leaf_clk net1 0.049971f
C3586 VPWR _147_ 0.283237f
C3587 _140_ _078_ 0.034132f
C3588 _159_ counter\[8\] 0.027563f
C3589 _326_/a_466_413# VPWR 0.024344f
C3590 net5 clknet_2_3__leaf_clk 0.028944f
C3591 _328_/a_193_47# divider\[2\] 0.03758f
C3592 _159_ _141_ 0.031882f
C3593 _094_ _219_/a_77_199# 0.010493f
C3594 VPWR _046_ 0.240692f
C3595 _336_/a_1062_300# clk 0.070416f
C3596 counter\[14\] counter\[9\] 0.039027f
C3597 counter\[13\] counter\[9\] 0.72165f
C3598 _039_ _037_ 0.030465f
C3599 _149_ counter\[1\] 0.078218f
C3600 net7 net3 0.323118f
C3601 _266_/a_215_53# divider\[2\] 0.027811f
C3602 counter\[0\] _065_ 0.05819f
C3603 counter\[0\] _341_/a_193_47# 0.050538f
C3604 _081_ _181_/a_250_297# 0.011952f
C3605 net6 _081_ 0.232132f
C3606 r2r_out[4] clk 0.528824f
C3607 _353_/a_466_413# VPWR 0.017821f
C3608 _066_ _233_/a_80_21# 0.043671f
C3609 counter\[6\] hold1/a_49_47# 0.083074f
C3610 counter\[10\] counter\[12\] 0.059368f
C3611 VGND _327_/a_634_159# -0.012168f
C3612 VPWR _327_/a_193_47# 0.012028f
C3613 _101_ _211_/a_27_47# 0.132963f
C3614 _346_/a_1059_315# _208_/a_76_199# 0.017544f
C3615 _094_ _118_ 0.101205f
C3616 VGND _350_/a_891_413# 0.024308f
C3617 VPWR _350_/a_1059_315# 0.017497f
C3618 clk _337_/a_1062_300# 0.021598f
C3619 divider\[4\] _268_/a_109_93# 0.021455f
C3620 net6 _005_ 0.03688f
C3621 clknet_0_clk _054_ 0.025323f
C3622 _345_/a_466_413# _021_ 0.046888f
C3623 counter\[13\] _248_/a_77_199# 0.041799f
C3624 clknet_2_3__leaf_clk _088_ 0.100474f
C3625 clknet_2_0__leaf_clk counter\[4\] 0.184451f
C3626 _240_/a_68_297# _054_ 0.015641f
C3627 _237_/a_27_47# _133_ 0.03328f
C3628 VPWR _279_/a_207_413# 0.046934f
C3629 _343_/a_1059_315# VGND 0.010373f
C3630 _072_ _073_ 0.208969f
C3631 _259_/a_27_47# rst 0.080949f
C3632 _103_ _102_ 0.346614f
C3633 VGND _357_/a_761_289# 0.013868f
C3634 VPWR _357_/a_193_47# 0.056746f
C3635 VGND _354_/a_1059_315# 0.017272f
C3636 VPWR _354_/a_466_413# 0.013039f
C3637 _352_/a_193_47# counter\[11\] 0.049594f
C3638 _307_/a_59_75# _078_ 0.046256f
C3639 _094_ _129_ 0.099169f
C3640 VGND _103_ 0.058211f
C3641 net13 counter\[6\] 0.104958f
C3642 _015_ VGND 0.220353f
C3643 _307_/a_59_75# _051_ 0.042457f
C3644 hold9/a_285_47# _335_/a_891_413# 0.015813f
C3645 _168_/a_76_199# net9 0.014954f
C3646 _053_ VGND 3.588297f
C3647 clknet_0_clk _225_/a_75_212# 0.020077f
C3648 clknet_2_1__leaf_clk _100_ 0.358519f
C3649 _053_ _324_/a_68_297# 0.05629f
C3650 _261_/a_215_297# net1 0.070826f
C3651 hold9/a_391_47# r2r_out[2] 0.057534f
C3652 counter\[14\] _046_ 0.024829f
C3653 _349_/a_1059_315# counter\[8\] 0.053201f
C3654 counter\[13\] _046_ 0.227349f
C3655 _136_ _121_ 0.02766f
C3656 VGND _292_/a_516_297# 0.015688f
C3657 _224_/a_59_75# counter\[8\] 0.055112f
C3658 _092_ rst 0.044497f
C3659 VPWR _126_ 0.319357f
C3660 VPWR rst 2.358003f
C3661 counter\[1\] _065_ 0.185157f
C3662 VPWR _030_ 0.355935f
C3663 VGND hold7/a_285_47# 0.074198f
C3664 _346_/a_381_47# _022_ 0.02431f
C3665 VPWR _272_/a_27_413# 0.060257f
C3666 _318_/a_27_47# r2r_out[0] 0.034203f
C3667 net2 net1 0.120247f
C3668 _011_ _335_/a_193_47# 0.065484f
C3669 input5/a_27_47# rst 0.010374f
C3670 _287_/a_215_53# VGND -0.01719f
C3671 net9 net1 0.022748f
C3672 net2 net5 0.041079f
C3673 _063_ _064_ 0.024657f
C3674 r2r_out[1] _058_ 0.087847f
C3675 VPWR _259_/a_27_47# 0.096003f
C3676 VPWR _325_/a_193_47# 0.037886f
C3677 _078_ _200_/a_77_199# 0.018359f
C3678 r2r_out[1] _071_ 0.416823f
C3679 VGND _291_/a_27_47# 0.012005f
C3680 VPWR _241_/a_59_75# 0.01619f
C3681 _291_/a_27_47# divider\[3\] 0.034625f
C3682 _135_ _078_ 0.0403f
C3683 _251_/a_27_47# counter\[9\] 0.015116f
C3684 _057_ _255_/a_80_21# 0.017168f
C3685 _032_ clknet_2_3__leaf_clk 0.038427f
C3686 VGND _298_/a_103_199# 0.042187f
C3687 _355_/a_634_159# VGND -0.013359f
C3688 _355_/a_193_47# VPWR 0.042708f
C3689 _342_/a_27_47# clknet_2_1__leaf_clk 0.092f
C3690 _325_/a_27_47# net8 0.437392f
C3691 net7 divider\[2\] 0.023675f
C3692 divider\[7\] net10 0.166807f
C3693 VPWR _332_/a_634_159# 0.02371f
C3694 VGND _332_/a_466_413# 0.017037f
C3695 _149_ _127_ 0.029551f
C3696 _117_ _133_ 0.250423f
C3697 divider\[1\] net4 0.919465f
C3698 _040_ VPWR 0.624263f
C3699 _348_/a_1059_315# clknet_2_0__leaf_clk 0.067436f
C3700 _149_ _001_ 0.377058f
C3701 _094_ _238_/a_77_199# 0.030207f
C3702 _069_ _068_ 0.127097f
C3703 VPWR _107_ 0.141626f
C3704 divider\[6\] _158_ 0.045124f
C3705 net14 _107_ 0.122694f
C3706 net1 net12 0.010559f
C3707 VGND _190_/a_489_47# 0.038838f
C3708 clknet_0_clk _243_/a_93_21# 0.012799f
C3709 _092_ VPWR 0.023096f
C3710 VGND _104_ 0.025686f
C3711 _054_ _078_ 0.210507f
C3712 _287_/a_215_53# _037_ 0.018942f
C3713 net14 VPWR 0.08492f
C3714 _332_/a_193_47# _008_ 0.094372f
C3715 _353_/a_1059_315# _066_ 0.019963f
C3716 _212_/a_80_21# _113_ 0.03093f
C3717 input5/a_27_47# VPWR 0.0802f
C3718 clkbuf_2_0__f_clk/a_110_47# hold6/a_285_47# 0.020048f
C3719 net9 _088_ 0.151564f
C3720 VPWR _171_/a_27_47# 0.049702f
C3721 r2r_out[1] _060_ 0.2048f
C3722 _268_/a_215_53# clknet_2_2__leaf_clk 0.090727f
C3723 VPWR _014_ 0.172228f
C3724 net5 clknet_2_2__leaf_clk 0.080116f
C3725 r2r_out[6] _084_ 0.042286f
C3726 VGND net8 1.417822f
C3727 _149_ net10 0.250714f
C3728 _170_/a_81_21# r2r_out[5] 0.0605f
C3729 VGND _008_ 0.15395f
C3730 divider\[3\] net8 0.162487f
C3731 _015_ _087_ 0.029612f
C3732 _053_ _087_ 0.098039f
C3733 _333_/a_381_47# _009_ 0.017746f
C3734 counter\[10\] _128_ 0.234076f
C3735 input10/a_27_47# load_divider 0.054459f
C3736 _094_ _035_ 0.014273f
C3737 _053_ _075_ 0.085908f
C3738 VPWR _080_ 0.244599f
C3739 _040_ _294_/a_78_199# 0.07876f
C3740 divider\[4\] _329_/a_891_413# 0.027893f
C3741 net10 _271_/a_29_53# 0.040891f
C3742 _076_ clknet_2_3__leaf_clk 0.045994f
C3743 _325_/a_27_47# net6 0.085025f
C3744 counter\[6\] _101_ 0.278897f
C3745 counter\[10\] _059_ 0.016126f
C3746 _336_/a_475_413# net21 0.010515f
C3747 _267_/a_215_297# _148_ 0.010244f
C3748 _334_/a_634_183# VPWR 0.044454f
C3749 _151_ net1 0.017194f
C3750 _053_ _066_ 0.213373f
C3751 _188_/a_27_47# VPWR 0.04233f
C3752 _273_/a_215_53# net10 0.038173f
C3753 _343_/a_891_413# _065_ 0.019736f
C3754 _053_ r2r_out[0] 0.035528f
C3755 _339_/a_475_413# _057_ 0.026322f
C3756 _353_/a_1059_315# clkbuf_0_clk/a_110_47# 0.017258f
C3757 _127_ _065_ 0.418467f
C3758 _155_ divider\[2\] 0.015444f
C3759 _284_/a_207_413# divider\[6\] 0.012894f
C3760 _040_ counter\[13\] 0.038153f
C3761 _314_/a_113_297# _064_ 0.044413f
C3762 VGND _181_/a_250_297# 0.019034f
C3763 VPWR _181_/a_93_21# 0.010833f
C3764 _140_ counter\[11\] 0.02421f
C3765 divider\[6\] _148_ 0.149346f
C3766 VGND net6 2.747798f
C3767 VPWR _116_ 0.019382f
C3768 _114_ VPWR 1.08376f
C3769 VGND _049_ 0.607384f
C3770 clknet_2_0__leaf_clk _350_/a_634_159# 0.010932f
C3771 divider\[3\] net6 0.028925f
C3772 _048_ _078_ 0.12228f
C3773 VPWR counter\[14\] 2.109343f
C3774 input8/a_27_47# VPWR 0.07305f
C3775 VPWR _330_/a_27_47# 0.132146f
C3776 VGND _330_/a_193_47# -0.049433f
C3777 _010_ VGND 0.100824f
C3778 VPWR counter\[13\] 1.504833f
C3779 VGND counter\[12\] 0.7846f
C3780 _351_/a_193_47# _027_ 0.051695f
C3781 _355_/a_1059_315# net4 0.060121f
C3782 _048_ _051_ 0.031638f
C3783 _320_/a_80_21# _054_ 0.015109f
C3784 _053_ _057_ 1.780349f
C3785 _173_/a_193_297# _077_ 0.030041f
C3786 divider\[0\] net3 0.026424f
C3787 _338_/a_193_47# r2r_out[5] 0.249495f
C3788 counter\[9\] _228_/a_27_47# 0.015738f
C3789 _078_ clknet_2_3__leaf_clk 0.132218f
C3790 clknet_2_1__leaf_clk _058_ 0.269554f
C3791 clknet_0_clk net9 1.660018f
C3792 _083_ r2r_out[5] 0.059941f
C3793 counter\[10\] _233_/a_217_297# 0.027124f
C3794 _355_/a_634_159# _066_ 0.023671f
C3795 divider\[4\] _034_ 0.011101f
C3796 _243_/a_93_21# _078_ 0.019908f
C3797 VGND _344_/a_27_47# 0.046168f
C3798 _160_ _281_/a_27_47# 0.016356f
C3799 _049_ counter\[15\] 0.038917f
C3800 _262_/a_215_53# net3 0.0597f
C3801 _094_ counter\[3\] 0.186836f
C3802 _094_ _190_/a_206_369# 0.031728f
C3803 _334_/a_193_47# _010_ 0.034146f
C3804 VGND _349_/a_27_47# 0.032326f
C3805 _148_ net4 0.209143f
C3806 _083_ _077_ 0.076043f
C3807 _141_ counter\[8\] 0.017817f
C3808 r2r_out[3] hold9/a_285_47# 0.097959f
C3809 VPWR _106_ 0.054243f
C3810 VGND _108_ 0.336763f
C3811 _141_ _143_ 0.329789f
C3812 VGND _068_ 0.020616f
C3813 _329_/a_381_47# net10 0.01692f
C3814 _053_ _336_/a_381_47# 0.019928f
C3815 _060_ clknet_2_1__leaf_clk 0.323053f
C3816 r2r_out[6] _340_/a_193_47# 0.010265f
C3817 VGND _341_/a_1059_315# -0.015239f
C3818 divider\[4\] _045_ 0.02206f
C3819 _329_/a_1059_315# clknet_2_2__leaf_clk 0.057928f
C3820 _094_ hold4/a_391_47# 0.051221f
C3821 counter\[13\] counter\[14\] 0.046545f
C3822 hold8/a_285_47# _054_ 0.071956f
C3823 _053_ _013_ 0.02328f
C3824 VPWR _347_/a_466_413# 0.018651f
C3825 net11 net12 0.013215f
C3826 _003_ _327_/a_193_47# 0.066565f
C3827 _152_ _327_/a_891_413# 0.016414f
C3828 _250_/a_113_297# _143_ 0.054228f
C3829 VPWR _122_ 0.095068f
C3830 _343_/a_466_413# counter\[2\] 0.034061f
C3831 _329_/a_466_413# _329_/a_27_47# -0.013083f
C3832 _155_ _042_ 0.024691f
C3833 divider\[4\] _289_/a_76_199# 0.027786f
C3834 _083_ _338_/a_381_47# 0.014758f
C3835 counter\[5\] _207_/a_35_297# 0.093803f
C3836 _326_/a_27_47# clknet_2_3__leaf_clk 0.099555f
C3837 counter\[0\] net16 0.250305f
C3838 _345_/a_891_413# hold2/a_285_47# 0.012799f
C3839 net4 _145_ 0.027022f
C3840 _315_/a_27_47# _078_ 0.017942f
C3841 _060_ r2r_out[6] 0.02414f
C3842 _274_/a_215_297# rst 0.016849f
C3843 _071_ _322_/a_27_47# 0.033467f
C3844 _251_/a_27_47# VPWR 0.035484f
C3845 _063_ clkbuf_2_1__f_clk/a_110_47# 0.014173f
C3846 _149_ _212_/a_80_21# 0.023464f
C3847 counter\[15\] _280_/a_27_413# 0.038462f
C3848 net6 _066_ 0.087528f
C3849 _149_ _094_ 0.084011f
C3850 net17 _098_ 0.273652f
C3851 VPWR _023_ 0.202663f
C3852 net2 _078_ 1.555665f
C3853 _330_/a_1059_315# _156_ 0.036443f
C3854 _066_ counter\[12\] 0.049707f
C3855 _078_ net9 0.389367f
C3856 VGND _169_/a_240_47# -0.015806f
C3857 _326_/a_1059_315# _002_ 0.034836f
C3858 _051_ net9 0.092015f
C3859 _208_/a_76_199# _066_ 0.027691f
C3860 VGND _128_ 0.033575f
C3861 counter\[4\] hold2/a_49_47# 0.030966f
C3862 _335_/a_27_47# _335_/a_193_47# -0.01246f
C3863 r2r_out[1] _333_/a_193_47# 0.03118f
C3864 _003_ rst 0.018535f
C3865 VPWR hold5/a_49_47# 0.038232f
C3866 VGND hold5/a_285_47# -0.021411f
C3867 _071_ _072_ 0.018806f
C3868 net10 data[3] 0.107727f
C3869 r2r_out[4] _170_/a_81_21# 0.055548f
C3870 _152_ clknet_2_2__leaf_clk 0.27968f
C3871 VGND _059_ 0.344493f
C3872 _287_/a_109_93# _038_ 0.019022f
C3873 _126_ _233_/a_80_21# 0.093279f
C3874 _149_ _347_/a_891_413# 0.014503f
C3875 _253_/a_215_47# counter\[14\] 0.045051f
C3876 _320_/a_80_21# _067_ 0.031786f
C3877 _074_ _054_ 0.042202f
C3878 _274_/a_215_297# VPWR 0.019346f
C3879 _078_ _098_ 0.091848f
C3880 _109_ counter\[4\] 0.048461f
C3881 _071_ _011_ 0.022346f
C3882 _057_ counter\[12\] 0.04775f
C3883 _149_ clk 0.08376f
C3884 counter\[1\] net16 0.106988f
C3885 _238_/a_77_199# _131_ 0.012756f
C3886 _065_ _344_/a_193_47# 0.027739f
C3887 _105_ counter\[4\] 0.02119f
C3888 counter\[12\] clkbuf_0_clk/a_110_47# 0.036954f
C3889 _274_/a_27_413# net8 0.022762f
C3890 _053_ r2r_out[3] 0.276552f
C3891 counter\[0\] _102_ 0.032268f
C3892 _097_ counter\[3\] 0.18194f
C3893 _149_ clknet_2_0__leaf_clk 0.440391f
C3894 _066_ _108_ 0.22079f
C3895 net8 _276_/a_215_297# 0.034297f
C3896 net18 _119_ 0.036572f
C3897 _159_ _281_/a_27_47# 0.043222f
C3898 _125_ _124_ 0.311994f
C3899 _306_/a_113_297# _056_ 0.016965f
C3900 _072_ _060_ 0.024914f
C3901 _068_ r2r_out[0] 0.024949f
C3902 _051_ clknet_2_2__leaf_clk 0.025602f
C3903 VPWR counter\[2\] 0.207038f
C3904 _251_/a_27_47# counter\[14\] 0.016864f
C3905 VGND counter\[0\] 1.408198f
C3906 clknet_2_1__leaf_clk net1 0.021589f
C3907 _269_/a_215_297# rst 0.055617f
C3908 _251_/a_27_47# counter\[13\] 0.0107f
C3909 _094_ _065_ 0.182006f
C3910 _114_ _023_ 0.010318f
C3911 _090_ clknet_2_3__leaf_clk 0.024071f
C3912 divider\[4\] _035_ 0.121254f
C3913 _053_ _002_ 0.012958f
C3914 _003_ VPWR 0.159594f
C3915 counter\[1\] _195_/a_227_47# 0.099259f
C3916 VGND load_divider 0.064691f
C3917 _097_ clkbuf_2_1__f_clk/a_110_47# 0.035465f
C3918 _057_ _252_/a_81_21# 0.068668f
C3919 _326_/a_27_47# net2 0.010637f
C3920 _347_/a_1059_315# _066_ 0.015225f
C3921 _356_/a_1059_315# VGND 0.013684f
C3922 _057_ _349_/a_27_47# 0.01812f
C3923 _097_ hold4/a_391_47# 0.014596f
C3924 _256_/a_266_47# _146_ 0.044727f
C3925 VGND _331_/a_27_47# 0.04811f
C3926 _246_/a_113_297# _133_ 0.017461f
C3927 _159_ divider\[2\] 0.420752f
C3928 VPWR _342_/a_891_413# 0.023948f
C3929 _005_ net10 0.03138f
C3930 _163_/a_27_47# _054_ 0.042256f
C3931 counter\[4\] _211_/a_27_47# 0.032488f
C3932 net7 net1 0.022171f
C3933 data[7] data[6] 0.042577f
C3934 _057_ _333_/a_381_47# 0.010749f
C3935 _208_/a_489_47# counter\[5\] 0.045606f
C3936 net7 net5 1.062037f
C3937 _167_/a_27_47# VPWR 0.161408f
C3938 divider\[4\] _292_/a_85_193# 0.036876f
C3939 VGND _124_ 0.041812f
C3940 _065_ clk 0.024574f
C3941 VPWR _263_/a_27_413# 0.060003f
C3942 VPWR _269_/a_215_297# 0.023665f
C3943 _356_/a_1059_315# counter\[15\] 0.070391f
C3944 counter\[1\] _102_ 0.094375f
C3945 r2r_out[6] _179_/a_79_21# 0.063499f
C3946 _261_/a_27_413# _150_ 0.05294f
C3947 clknet_2_0__leaf_clk _065_ 0.116992f
C3948 _213_/a_215_53# _118_ 0.026758f
C3949 VPWR hold9/a_285_47# 0.011088f
C3950 net4 _161_ 0.014872f
C3951 r2r_out[7] clk 0.528315f
C3952 VGND counter\[1\] 1.1994f
C3953 net4 _054_ 0.122201f
C3954 _149_ _097_ 0.028051f
C3955 _144_ _252_/a_299_297# 0.016912f
C3956 _053_ _339_/a_634_183# 0.011336f
C3957 VPWR _082_ 0.103401f
C3958 _224_/a_59_75# _120_ 0.062843f
C3959 VPWR _255_/a_80_21# 0.099493f
C3960 divider\[6\] _331_/a_634_159# 0.016074f
C3961 _347_/a_193_47# clknet_2_0__leaf_clk 0.087403f
C3962 counter\[4\] _205_/a_109_93# 0.010519f
C3963 _039_ VPWR 0.15011f
C3964 VPWR _318_/a_27_47# 0.027541f
C3965 clknet_2_1__leaf_clk _333_/a_193_47# 0.012493f
C3966 _084_ _085_ 0.054237f
C3967 _066_ _059_ 0.025974f
C3968 divider\[2\] _283_/a_78_199# 0.026286f
C3969 r2r_out[5] clknet_2_3__leaf_clk 0.350947f
C3970 _065_ _130_ 0.029885f
C3971 net2 hold8/a_285_47# 0.013293f
C3972 _356_/a_891_413# _149_ 0.019388f
C3973 _353_/a_634_159# _029_ 0.047991f
C3974 _347_/a_466_413# _023_ 0.043116f
C3975 _286_/a_219_297# divider\[6\] 0.036233f
C3976 hold5/a_391_47# _065_ 0.02134f
C3977 net10 _327_/a_27_47# 0.012527f
C3978 _082_ _080_ 0.039193f
C3979 _057_ _169_/a_240_47# 0.039812f
C3980 _089_ _060_ 0.011743f
C3981 _127_ _026_ 0.056433f
C3982 _136_ _138_ 0.190751f
C3983 _334_/a_193_47# counter\[1\] 0.012217f
C3984 _090_ net9 0.075749f
C3985 _052_ _124_ 0.02658f
C3986 _326_/a_1059_315# VPWR 0.027417f
C3987 _077_ clknet_2_3__leaf_clk 0.250394f
C3988 _229_/a_77_199# _125_ 0.063729f
C3989 _140_ _045_ 0.072592f
C3990 _167_/a_27_47# counter\[13\] 0.022082f
C3991 net6 _269_/a_27_413# 0.010061f
C3992 _336_/a_891_413# clk 0.040322f
C3993 counter\[12\] counter\[9\] 0.378942f
C3994 r2r_out[1] _061_ 0.07588f
C3995 _057_ _059_ 0.028015f
C3996 _053_ rst 0.650342f
C3997 VGND _238_/a_227_47# 0.034253f
C3998 _354_/a_27_47# clknet_2_2__leaf_clk 0.256695f
C3999 _291_/a_193_297# _035_ 0.012809f
C4000 _059_ clkbuf_0_clk/a_110_47# 0.011207f
C4001 _101_ _216_/a_59_75# 0.026193f
C4002 counter\[0\] _341_/a_634_159# 0.042893f
C4003 _227_/a_59_75# counter\[8\] 0.031254f
C4004 _149_ _186_/a_113_297# 0.011205f
C4005 clknet_0_clk clknet_2_1__leaf_clk 0.159174f
C4006 _325_/a_27_47# _001_ 0.026425f
C4007 _353_/a_1059_315# VPWR 0.017704f
C4008 _066_ _233_/a_217_297# 0.057871f
C4009 counter\[6\] hold1/a_285_47# 0.076316f
C4010 _025_ _349_/a_466_413# 0.029008f
C4011 _339_/a_1062_300# VGND 0.076786f
C4012 counter\[14\] _255_/a_80_21# 0.015048f
C4013 _094_ _119_ 0.059069f
C4014 VGND _062_ 0.03586f
C4015 net4 clknet_2_3__leaf_clk 0.34554f
C4016 counter\[5\] _021_ 0.016652f
C4017 _343_/a_1059_315# VPWR 0.030193f
C4018 _044_ _035_ 0.02158f
C4019 VGND _229_/a_77_199# 0.012444f
C4020 VPWR _357_/a_761_289# 0.040595f
C4021 divider\[5\] _156_ 0.222194f
C4022 VPWR _354_/a_1059_315# 0.060512f
C4023 _352_/a_634_159# counter\[11\] 0.01588f
C4024 _149_ divider\[4\] 0.027615f
C4025 VGND _127_ 0.196633f
C4026 counter\[6\] counter\[4\] 0.111818f
C4027 VPWR _103_ 0.268164f
C4028 VGND _001_ 0.044342f
C4029 counter\[12\] _137_ 0.240177f
C4030 _076_ _337_/a_27_47# 0.048866f
C4031 VGND _352_/a_27_47# 0.047411f
C4032 _015_ VPWR 0.16253f
C4033 _053_ VPWR 4.966164f
C4034 _155_ _156_ 0.01483f
C4035 counter\[1\] _066_ 0.010684f
C4036 _325_/a_27_47# _325_/a_466_413# -0.013083f
C4037 _332_/a_27_47# _158_ 0.08344f
C4038 _256_/a_81_21# _143_ 0.013006f
C4039 clkbuf_2_0__f_clk/a_110_47# _078_ 0.031406f
C4040 VGND input9/a_27_47# 0.024753f
C4041 _053_ _014_ 0.0742f
C4042 counter\[10\] _094_ 0.095794f
C4043 _349_/a_891_413# counter\[8\] 0.016042f
C4044 _148_ _150_ 0.125312f
C4045 _113_ _211_/a_27_47# 0.020727f
C4046 VPWR _292_/a_516_297# 0.062496f
C4047 counter\[9\] _280_/a_27_413# 0.025858f
C4048 VGND net10 2.01754f
C4049 _044_ _292_/a_85_193# 0.012619f
C4050 VGND hold7/a_391_47# 0.037064f
C4051 VPWR _272_/a_215_297# 0.047712f
C4052 VGND _029_ 0.484419f
C4053 divider\[3\] net10 0.20497f
C4054 net21 _335_/a_475_413# 0.010993f
C4055 _115_ _237_/a_27_47# 0.048301f
C4056 _287_/a_109_93# VGND -0.012163f
C4057 _287_/a_215_53# VPWR 0.01193f
C4058 divider\[6\] net9 0.220007f
C4059 _149_ _261_/a_27_413# 0.047449f
C4060 _149_ divider\[1\] 0.338226f
C4061 _067_ net4 0.069097f
C4062 _077_ net9 0.029812f
C4063 _351_/a_381_47# clknet_2_0__leaf_clk 0.015919f
C4064 VGND net18 0.035527f
C4065 net8 rst 0.047715f
C4066 hold7/a_49_47# _303_/a_113_297# 0.021797f
C4067 _040_ _298_/a_103_199# 0.082141f
C4068 net8 _272_/a_27_413# 0.03731f
C4069 VPWR _325_/a_634_159# 0.042254f
C4070 _291_/a_109_297# divider\[3\] 0.010312f
C4071 VPWR _298_/a_103_199# 0.04748f
C4072 _355_/a_634_159# VPWR 0.022051f
C4073 _025_ clknet_2_1__leaf_clk 0.010575f
C4074 _342_/a_193_47# clknet_2_1__leaf_clk 0.462626f
C4075 divider\[7\] _158_ 0.082896f
C4076 _325_/a_193_47# net8 0.080981f
C4077 counter\[15\] net10 0.111829f
C4078 _140_ _035_ 0.214833f
C4079 divider\[4\] _041_ 0.729783f
C4080 clknet_2_1__leaf_clk _078_ 1.630148f
C4081 VPWR _332_/a_466_413# 0.02017f
C4082 VGND _332_/a_1059_315# 0.042582f
C4083 _078_ _133_ 1.077864f
C4084 _149_ net20 0.029783f
C4085 _120_ counter\[8\] 0.070754f
C4086 _018_ clknet_2_1__leaf_clk 0.110206f
C4087 _348_/a_891_413# clknet_2_0__leaf_clk 0.035776f
C4088 _071_ _317_/a_113_297# 0.021169f
C4089 divider\[0\] net1 0.507471f
C4090 _355_/a_27_47# _031_ 0.053694f
C4091 _051_ _133_ 0.166574f
C4092 counter\[10\] clknet_2_0__leaf_clk 0.010415f
C4093 _152_ net7 0.023734f
C4094 divider\[0\] net5 0.122827f
C4095 _053_ counter\[14\] 0.011876f
C4096 VPWR _104_ 0.031894f
C4097 _274_/a_27_413# _331_/a_27_47# 0.012449f
C4098 net2 net4 0.018976f
C4099 _281_/a_27_47# counter\[8\] 0.011933f
C4100 _212_/a_209_297# _113_ 0.037145f
C4101 divider\[6\] clknet_2_2__leaf_clk 0.069732f
C4102 net4 net9 0.098623f
C4103 _262_/a_215_53# net1 0.016131f
C4104 _268_/a_109_93# clknet_2_2__leaf_clk 0.06573f
C4105 _084_ _086_ 0.243254f
C4106 _089_ _088_ 0.098203f
C4107 _031_ VGND 0.051344f
C4108 _091_ _178_/a_75_199# 0.012092f
C4109 net6 rst 0.194724f
C4110 counter\[9\] _059_ 0.083628f
C4111 VPWR net8 3.493228f
C4112 VPWR _008_ 0.182402f
C4113 net6 _272_/a_27_413# 0.052922f
C4114 _170_/a_299_297# r2r_out[5] 0.039427f
C4115 _294_/a_78_199# _298_/a_103_199# 0.014491f
C4116 counter\[10\] _130_ 0.110538f
C4117 _062_ r2r_out[0] 0.014939f
C4118 _069_ clk 0.069365f
C4119 divider\[4\] _329_/a_381_47# 0.016435f
C4120 _066_ _229_/a_77_199# 0.010555f
C4121 r2r_out[4] clknet_2_3__leaf_clk 0.248185f
C4122 _115_ _117_ 0.766136f
C4123 clknet_0_clk _138_ 0.138014f
C4124 _066_ _127_ 0.041482f
C4125 _325_/a_193_47# net6 0.259108f
C4126 _285_/a_35_297# divider\[7\] 0.050432f
C4127 _342_/a_27_47# _096_ 0.017222f
C4128 _094_ net16 0.035238f
C4129 _072_ _076_ 0.030757f
C4130 _334_/a_1062_300# VGND 0.080483f
C4131 _334_/a_475_413# VPWR 0.044728f
C4132 _273_/a_109_93# net10 0.042658f
C4133 _339_/a_1062_300# _057_ 0.016274f
C4134 _353_/a_634_159# clk 0.013493f
C4135 _298_/a_103_199# counter\[13\] 0.021107f
C4136 net4 clknet_2_2__leaf_clk 0.064675f
C4137 clk _340_/a_1062_300# 0.014989f
C4138 _101_ _192_/a_27_47# 0.017022f
C4139 _094_ _125_ 0.229874f
C4140 VGND _338_/a_27_47# 0.043643f
C4141 VPWR _181_/a_250_297# 0.044908f
C4142 _066_ _029_ 0.05961f
C4143 VPWR net6 0.748355f
C4144 VPWR _049_ 0.21445f
C4145 _123_ counter\[8\] 0.21375f
C4146 clknet_2_0__leaf_clk _350_/a_466_413# 0.01806f
C4147 _149_ _105_ 0.069346f
C4148 VPWR _330_/a_193_47# 0.080895f
C4149 _117_ counter\[8\] 0.163072f
C4150 _010_ VPWR 0.323876f
C4151 VPWR counter\[12\] 1.104291f
C4152 _356_/a_27_47# clknet_2_3__leaf_clk 0.013308f
C4153 _355_/a_891_413# net4 0.045366f
C4154 counter\[6\] _113_ 0.030627f
C4155 VGND _258_/a_27_47# 0.03222f
C4156 VPWR _208_/a_76_199# 0.01861f
C4157 _353_/a_27_47# clknet_2_1__leaf_clk 0.012644f
C4158 _149_ _148_ 0.911095f
C4159 _338_/a_634_183# r2r_out[5] 0.021871f
C4160 _065_ _091_ 0.030984f
C4161 VGND _205_/a_215_53# -0.022139f
C4162 net6 _080_ 0.061665f
C4163 _342_/a_1059_315# counter\[1\] 0.014163f
C4164 _355_/a_466_413# _066_ 0.025128f
C4165 _243_/a_250_297# _078_ 0.087496f
C4166 counter\[9\] _124_ 0.171385f
C4167 _169_/a_51_297# net9 0.015596f
C4168 _348_/a_27_47# _348_/a_466_413# -0.013083f
C4169 _348_/a_193_47# _348_/a_634_159# -0.016573f
C4170 VGND _344_/a_193_47# -0.10547f
C4171 VPWR _344_/a_27_47# -0.193055f
C4172 clknet_2_0__leaf_clk _026_ 0.38766f
C4173 _262_/a_109_93# net3 0.019806f
C4174 VPWR _252_/a_81_21# 0.022243f
C4175 _054_ _056_ 0.040096f
C4176 _264_/a_215_53# data[3] 0.054346f
C4177 _094_ _102_ 0.092074f
C4178 VGND _212_/a_80_21# 0.027746f
C4179 _343_/a_27_47# clknet_2_1__leaf_clk 0.031236f
C4180 _328_/a_891_413# rst 0.010711f
C4181 VPWR _349_/a_27_47# 0.089131f
C4182 VGND _349_/a_193_47# -0.033802f
C4183 VGND _094_ 1.397535f
C4184 data[6] net9 0.059095f
C4185 r2r_out[3] hold9/a_391_47# 0.066577f
C4186 _060_ _079_ 0.552293f
C4187 VPWR _108_ 0.064121f
C4188 VPWR _068_ 0.19504f
C4189 _031_ _066_ 0.035498f
C4190 _138_ _078_ 0.023948f
C4191 net6 _181_/a_93_21# 0.055647f
C4192 _348_/a_27_47# _024_ 0.032939f
C4193 net19 clknet_2_1__leaf_clk 0.19679f
C4194 _065_ _020_ 0.294559f
C4195 VPWR _341_/a_1059_315# 0.011201f
C4196 VGND _341_/a_891_413# -0.010827f
C4197 _044_ _041_ 0.167564f
C4198 VGND _146_ 0.228656f
C4199 _329_/a_891_413# clknet_2_2__leaf_clk 0.044436f
C4200 _112_ _094_ 0.018126f
C4201 _049_ counter\[14\] 0.063143f
C4202 counter\[12\] counter\[14\] 0.064401f
C4203 hold8/a_391_47# _054_ 0.059626f
C4204 counter\[13\] counter\[12\] 0.286627f
C4205 VGND _280_/a_207_413# 0.015658f
C4206 VPWR _347_/a_1059_315# 0.015293f
C4207 _244_/a_59_75# _139_ 0.024102f
C4208 net11 _000_ 0.260829f
C4209 _343_/a_1059_315# counter\[2\] 0.059166f
C4210 _020_ 0 0.139788f
C4211 _104_ 0 0.143482f
C4212 counter\[6\] 0 0.511237f
C4213 _023_ 0 0.172897f
C4214 _347_/a_381_47# 0 0.015369f
C4215 _347_/a_891_413# 0 0.161052f
C4216 _347_/a_1059_315# 0 0.248849f
C4217 _347_/a_466_413# 0 0.133203f
C4218 _347_/a_634_159# 0 0.142309f
C4219 _347_/a_193_47# 0 0.284262f
C4220 _347_/a_27_47# 0 0.449511f
C4221 VPWR 0 0.494483p
C4222 VGND 0 0.156041p
C4223 _160_ 0 0.129815f
C4224 divider\[1\] 0 0.412489f
C4225 _278_/a_27_53# 0 0.175308f
C4226 _278_/a_219_297# 0 0.137194f
C4227 _105_ 0 0.124266f
C4228 net14 0 0.119432f
C4229 counter\[7\] 0 0.594844f
C4230 _024_ 0 0.184261f
C4231 _348_/a_381_47# 0 0.015369f
C4232 _348_/a_891_413# 0 0.161052f
C4233 _348_/a_1059_315# 0 0.248849f
C4234 _348_/a_466_413# 0 0.133203f
C4235 _348_/a_634_159# 0 0.142309f
C4236 _348_/a_193_47# 0 0.284262f
C4237 _348_/a_27_47# 0 0.449511f
C4238 divider\[0\] 0 0.284172f
C4239 _279_/a_207_413# 0 0.137402f
C4240 _279_/a_27_413# 0 0.196502f
C4241 _049_ 0 0.195114f
C4242 _296_/a_27_53# 0 0.175308f
C4243 _296_/a_219_297# 0 0.137194f
C4244 _349_/a_381_47# 0 0.015369f
C4245 _349_/a_891_413# 0 0.161052f
C4246 _349_/a_1059_315# 0 0.248849f
C4247 _349_/a_466_413# 0 0.133203f
C4248 _349_/a_634_159# 0 0.142309f
C4249 _349_/a_193_47# 0 0.284262f
C4250 _349_/a_27_47# 0 0.449511f
C4251 _050_ 0 0.147091f
C4252 _297_/a_215_47# 0 0.01011f
C4253 _297_/a_79_21# 0 0.225128f
C4254 _101_ 0 0.916798f
C4255 _120_ 0 0.14294f
C4256 _221_/a_68_297# 0 0.153866f
C4257 _043_ 0 0.242838f
C4258 _047_ 0 0.088296f
C4259 _298_/a_253_47# 0 0.011031f
C4260 _298_/a_103_199# 0 0.196442f
C4261 _108_ 0 0.133143f
C4262 _106_ 0 0.142206f
C4263 _205_/a_109_93# 0 0.160708f
C4264 _205_/a_215_53# 0 0.142592f
C4265 _121_ 0 0.275415f
C4266 _045_ 0 0.263731f
C4267 _051_ 0 0.296787f
C4268 _080_ 0 0.119111f
C4269 r2r_out[5] 0 0.773589f
C4270 _170_/a_299_297# 0 0.034794f
C4271 _170_/a_81_21# 0 0.147141f
C4272 _206_/a_113_297# 0 0.034004f
C4273 _054_ 0 1.597855f
C4274 _059_ 0 0.350294f
C4275 _223_/a_250_297# 0 0.02777f
C4276 _223_/a_93_21# 0 0.150721f
C4277 _135_ 0 0.110228f
C4278 _240_/a_68_297# 0 0.153866f
C4279 _171_/a_27_47# 0 0.177187f
C4280 _109_ 0 0.104062f
C4281 _107_ 0 0.345335f
C4282 _207_/a_35_297# 0 0.254573f
C4283 hold9/a_391_47# 0 0.127705f
C4284 hold9/a_285_47# 0 0.29867f
C4285 hold9/a_49_47# 0 0.306903f
C4286 _122_ 0 0.14449f
C4287 _057_ 0 1.413733f
C4288 _224_/a_59_75# 0 0.177062f
C4289 _136_ 0 0.27487f
C4290 _241_/a_59_75# 0 0.177062f
C4291 _082_ 0 0.106064f
C4292 _081_ 0 0.474985f
C4293 clkbuf_2_3__f_clk/a_110_47# 0 1.73295f
C4294 _094_ 0 1.195606f
C4295 _066_ 0 1.46872f
C4296 _208_/a_489_47# 0 0.037211f
C4297 _208_/a_206_369# 0 0.153769f
C4298 _208_/a_76_199# 0 0.136541f
C4299 hold8/a_391_47# 0 0.127705f
C4300 hold8/a_285_47# 0 0.29867f
C4301 hold8/a_49_47# 0 0.306903f
C4302 _025_ 0 0.180417f
C4303 _123_ 0 0.170328f
C4304 _225_/a_75_212# 0 0.210264f
C4305 net2 0 0.285409f
C4306 _062_ 0 0.111631f
C4307 _311_/a_27_297# 0 0.190287f
C4308 _083_ 0 0.132825f
C4309 net6 0 0.371254f
C4310 _173_/a_27_47# 0 0.216317f
C4311 _095_ 0 0.141562f
C4312 _190_/a_489_47# 0 0.037211f
C4313 _190_/a_206_369# 0 0.153769f
C4314 _190_/a_76_199# 0 0.136541f
C4315 _022_ 0 0.190239f
C4316 _065_ 0 1.814524f
C4317 _110_ 0 0.200614f
C4318 hold7/a_391_47# 0 0.127705f
C4319 hold7/a_285_47# 0 0.29867f
C4320 hold7/a_49_47# 0 0.306903f
C4321 _124_ 0 0.248471f
C4322 counter\[9\] 0 0.84899f
C4323 _138_ 0 0.14067f
C4324 _137_ 0 0.102851f
C4325 _243_/a_250_297# 0 0.02777f
C4326 _243_/a_93_21# 0 0.150721f
C4327 _063_ 0 0.161343f
C4328 _014_ 0 0.165446f
C4329 _174_/a_215_47# 0 0.01011f
C4330 _174_/a_79_21# 0 0.225128f
C4331 _018_ 0 0.175898f
C4332 _096_ 0 0.212547f
C4333 _260_/a_109_93# 0 0.160708f
C4334 _260_/a_215_53# 0 0.142592f
C4335 hold6/a_391_47# 0 0.127705f
C4336 hold6/a_285_47# 0 0.29867f
C4337 hold6/a_49_47# 0 0.306903f
C4338 _227_/a_59_75# 0 0.177062f
C4339 _139_ 0 0.137918f
C4340 _244_/a_59_75# 0 0.177062f
C4341 _313_/a_27_47# 0 0.542977f
C4342 _084_ 0 0.2838f
C4343 r2r_out[6] 0 0.965787f
C4344 _097_ 0 0.335599f
C4345 counter\[0\] 0 0.951161f
C4346 counter\[2\] 0 0.576308f
C4347 _192_/a_27_47# 0 0.177187f
C4348 _006_ 0 0.180268f
C4349 _330_/a_381_47# 0 0.015369f
C4350 _330_/a_891_413# 0 0.161052f
C4351 _330_/a_1059_315# 0 0.248849f
C4352 _330_/a_466_413# 0 0.133203f
C4353 _330_/a_634_159# 0 0.142309f
C4354 _330_/a_193_47# 0 0.284262f
C4355 _330_/a_27_47# 0 0.449511f
C4356 _001_ 0 0.158742f
C4357 _150_ 0 0.184778f
C4358 _261_/a_215_297# 0 0.152836f
C4359 _261_/a_27_413# 0 0.171579f
C4360 net17 0 0.217366f
C4361 hold5/a_391_47# 0 0.127705f
C4362 hold5/a_285_47# 0 0.29867f
C4363 hold5/a_49_47# 0 0.306903f
C4364 counter\[8\] 0 0.733786f
C4365 _228_/a_27_47# 0 0.177187f
C4366 _029_ 0 0.194126f
C4367 _245_/a_75_212# 0 0.210264f
C4368 _064_ 0 0.111564f
C4369 _061_ 0 0.121096f
C4370 _314_/a_113_297# 0 0.034004f
C4371 _176_/a_68_297# 0 0.153866f
C4372 _193_/a_113_297# 0 0.034004f
C4373 _151_ 0 0.217983f
C4374 _262_/a_109_93# 0 0.160708f
C4375 _262_/a_215_53# 0 0.142592f
C4376 _007_ 0 0.164432f
C4377 _331_/a_381_47# 0 0.015369f
C4378 _331_/a_891_413# 0 0.161052f
C4379 _331_/a_1059_315# 0 0.248849f
C4380 _331_/a_466_413# 0 0.133203f
C4381 _331_/a_634_159# 0 0.142309f
C4382 _331_/a_193_47# 0 0.284262f
C4383 _331_/a_27_47# 0 0.449511f
C4384 hold4/a_391_47# 0 0.127705f
C4385 hold4/a_285_47# 0 0.29867f
C4386 hold4/a_49_47# 0 0.306903f
C4387 _126_ 0 0.471049f
C4388 _125_ 0 0.103379f
C4389 _229_/a_227_47# 0 0.030865f
C4390 _229_/a_77_199# 0 0.146762f
C4391 _140_ 0 0.115252f
C4392 counter\[12\] 0 0.850806f
C4393 counter\[13\] 0 1.031976f
C4394 _246_/a_113_297# 0 0.034004f
C4395 _315_/a_27_47# 0 0.542977f
C4396 _086_ 0 0.13159f
C4397 net7 0 0.367186f
C4398 _177_/a_59_75# 0 0.177062f
C4399 _008_ 0 0.166318f
C4400 _332_/a_381_47# 0 0.015369f
C4401 _332_/a_891_413# 0 0.161052f
C4402 _332_/a_1059_315# 0 0.248849f
C4403 _332_/a_466_413# 0 0.133203f
C4404 _332_/a_634_159# 0 0.142309f
C4405 _332_/a_193_47# 0 0.284262f
C4406 _332_/a_27_47# 0 0.449511f
C4407 _002_ 0 0.154364f
C4408 _263_/a_215_297# 0 0.152836f
C4409 _263_/a_27_413# 0 0.171579f
C4410 _280_/a_207_413# 0 0.137402f
C4411 _280_/a_27_413# 0 0.196502f
C4412 net15 0 0.143914f
C4413 hold3/a_391_47# 0 0.127705f
C4414 hold3/a_285_47# 0 0.29867f
C4415 hold3/a_49_47# 0 0.306903f
C4416 _087_ 0 0.115233f
C4417 _085_ 0 0.131682f
C4418 _178_/a_75_199# 0 0.20459f
C4419 _141_ 0 0.372285f
C4420 _247_/a_27_47# 0 0.177187f
C4421 net3 0 0.308777f
C4422 _333_/a_381_47# 0 0.016397f
C4423 _333_/a_891_413# 0 0.160892f
C4424 _333_/a_1062_300# 0 0.529662f
C4425 _333_/a_475_413# 0 0.137184f
C4426 _333_/a_634_183# 0 0.150209f
C4427 _333_/a_193_47# 0 0.271178f
C4428 _333_/a_27_47# 0 0.468295f
C4429 _099_ 0 0.143522f
C4430 _098_ 0 0.092047f
C4431 _195_/a_227_47# 0 0.030865f
C4432 _195_/a_77_199# 0 0.146762f
C4433 _264_/a_109_93# 0 0.160708f
C4434 _264_/a_215_53# 0 0.142592f
C4435 _026_ 0 0.206154f
C4436 _350_/a_381_47# 0 0.015369f
C4437 _350_/a_891_413# 0 0.161052f
C4438 _350_/a_1059_315# 0 0.248849f
C4439 _350_/a_466_413# 0 0.133203f
C4440 _350_/a_634_159# 0 0.142309f
C4441 _350_/a_193_47# 0 0.284262f
C4442 _350_/a_27_47# 0 0.449511f
C4443 _034_ 0 0.149276f
C4444 divider\[2\] 0 0.471944f
C4445 _161_ 0 0.121029f
C4446 _033_ 0 0.122585f
C4447 _281_/a_27_47# 0 0.216317f
C4448 hold2/a_391_47# 0 0.127705f
C4449 hold2/a_285_47# 0 0.29867f
C4450 hold2/a_49_47# 0 0.306903f
C4451 clkbuf_2_2__f_clk/a_110_47# 0 1.73295f
C4452 _068_ 0 0.102682f
C4453 r2r_out[2] 0 1.574642f
C4454 _317_/a_113_297# 0 0.034004f
C4455 _046_ 0 0.267328f
C4456 _248_/a_227_47# 0 0.030865f
C4457 _248_/a_77_199# 0 0.146762f
C4458 _179_/a_215_47# 0 0.01011f
C4459 _179_/a_79_21# 0 0.225128f
C4460 _019_ 0 0.166532f
C4461 _100_ 0 0.138217f
C4462 _003_ 0 0.16738f
C4463 _152_ 0 0.266852f
C4464 _265_/a_215_297# 0 0.152836f
C4465 _265_/a_27_413# 0 0.171579f
C4466 r2r_out[1] 0 1.313779f
C4467 _010_ 0 0.133868f
C4468 _334_/a_381_47# 0 0.016397f
C4469 _334_/a_891_413# 0 0.160892f
C4470 _334_/a_1062_300# 0 0.529662f
C4471 _334_/a_475_413# 0 0.137184f
C4472 _334_/a_634_183# 0 0.150209f
C4473 _334_/a_193_47# 0 0.271178f
C4474 _334_/a_27_47# 0 0.468295f
C4475 counter\[10\] 0 0.882194f
C4476 _027_ 0 0.144188f
C4477 _351_/a_381_47# 0 0.015369f
C4478 _351_/a_891_413# 0 0.161052f
C4479 _351_/a_1059_315# 0 0.248849f
C4480 _351_/a_466_413# 0 0.133203f
C4481 _351_/a_634_159# 0 0.142309f
C4482 _351_/a_193_47# 0 0.284262f
C4483 _351_/a_27_47# 0 0.449511f
C4484 hold1/a_391_47# 0 0.127705f
C4485 hold1/a_285_47# 0 0.29867f
C4486 hold1/a_49_47# 0 0.306903f
C4487 _069_ 0 0.293164f
C4488 _318_/a_27_47# 0 0.177187f
C4489 _142_ 0 0.163771f
C4490 _335_/a_381_47# 0 0.016397f
C4491 _335_/a_891_413# 0 0.160892f
C4492 _335_/a_1062_300# 0 0.529662f
C4493 _335_/a_475_413# 0 0.137184f
C4494 _335_/a_634_183# 0 0.150209f
C4495 _335_/a_193_47# 0 0.271178f
C4496 _335_/a_27_47# 0 0.468295f
C4497 _197_/a_27_47# 0 0.265166f
C4498 _153_ 0 0.215368f
C4499 _266_/a_109_93# 0 0.160708f
C4500 _266_/a_215_53# 0 0.142592f
C4501 counter\[11\] 0 0.496373f
C4502 _028_ 0 0.151063f
C4503 clknet_2_2__leaf_clk 0 1.365083f
C4504 _352_/a_381_47# 0 0.015369f
C4505 _352_/a_891_413# 0 0.161052f
C4506 _352_/a_1059_315# 0 0.248849f
C4507 _352_/a_466_413# 0 0.133203f
C4508 _352_/a_634_159# 0 0.142309f
C4509 _352_/a_193_47# 0 0.284262f
C4510 _352_/a_27_47# 0 0.449511f
C4511 _283_/a_215_47# 0 0.035725f
C4512 _283_/a_78_199# 0 0.15408f
C4513 ext_data 0 0.381423f
C4514 input9/a_27_47# 0 0.320141f
C4515 net9 0 0.897162f
C4516 _319_/a_29_53# 0 0.180006f
C4517 n_rst 0 0.373534f
C4518 input11/a_75_212# 0 0.210264f
C4519 _102_ 0 0.109635f
C4520 counter\[3\] 0 0.413211f
C4521 _012_ 0 0.164656f
C4522 clknet_2_3__leaf_clk 0 1.677769f
C4523 _336_/a_381_47# 0 0.016397f
C4524 _336_/a_891_413# 0 0.160892f
C4525 _336_/a_1062_300# 0 0.529662f
C4526 _336_/a_475_413# 0 0.137184f
C4527 _336_/a_634_183# 0 0.150209f
C4528 _336_/a_193_47# 0 0.271178f
C4529 _336_/a_27_47# 0 0.468295f
C4530 _004_ 0 0.157955f
C4531 _148_ 0 1.037932f
C4532 _267_/a_215_297# 0 0.152836f
C4533 _267_/a_27_413# 0 0.171579f
C4534 data[7] 0 0.370638f
C4535 input8/a_27_47# 0 0.207781f
C4536 _353_/a_381_47# 0 0.015369f
C4537 _353_/a_891_413# 0 0.161052f
C4538 _353_/a_1059_315# 0 0.248849f
C4539 _353_/a_466_413# 0 0.133203f
C4540 _353_/a_634_159# 0 0.142309f
C4541 _353_/a_193_47# 0 0.284262f
C4542 _353_/a_27_47# 0 0.449511f
C4543 _037_ 0 0.154114f
C4544 divider\[6\] 0 0.416701f
C4545 _284_/a_207_413# 0 0.137402f
C4546 _284_/a_27_413# 0 0.196502f
C4547 load_divider 0 0.467461f
C4548 input10/a_27_47# 0 0.320141f
C4549 _103_ 0 0.131058f
C4550 net16 0 0.228252f
C4551 _337_/a_381_47# 0 0.016397f
C4552 _337_/a_891_413# 0 0.160892f
C4553 _337_/a_1062_300# 0 0.529662f
C4554 _337_/a_475_413# 0 0.137184f
C4555 _337_/a_634_183# 0 0.150209f
C4556 _337_/a_193_47# 0 0.271178f
C4557 _337_/a_27_47# 0 0.468295f
C4558 _268_/a_109_93# 0 0.160708f
C4559 _268_/a_215_53# 0 0.142592f
C4560 data[6] 0 0.387893f
C4561 input7/a_27_47# 0 0.207781f
C4562 _030_ 0 0.188667f
C4563 _354_/a_381_47# 0 0.015369f
C4564 _354_/a_891_413# 0 0.161052f
C4565 _354_/a_1059_315# 0 0.248849f
C4566 _354_/a_466_413# 0 0.133203f
C4567 _354_/a_634_159# 0 0.142309f
C4568 _354_/a_193_47# 0 0.284262f
C4569 _354_/a_27_47# 0 0.449511f
C4570 _038_ 0 0.232612f
C4571 counter\[15\] 0 0.659376f
C4572 divider\[7\] 0 0.609766f
C4573 _285_/a_35_297# 0 0.254573f
C4574 _338_/a_381_47# 0 0.016397f
C4575 _338_/a_891_413# 0 0.160892f
C4576 _338_/a_1062_300# 0 0.529662f
C4577 _338_/a_475_413# 0 0.137184f
C4578 _338_/a_634_183# 0 0.150209f
C4579 _338_/a_193_47# 0 0.271178f
C4580 _338_/a_27_47# 0 0.468295f
C4581 _005_ 0 0.168656f
C4582 _154_ 0 0.230824f
C4583 _269_/a_215_297# 0 0.152836f
C4584 _269_/a_27_413# 0 0.171579f
C4585 data[5] 0 0.413225f
C4586 input6/a_27_47# 0 0.207781f
C4587 _031_ 0 0.167774f
C4588 _355_/a_381_47# 0 0.015369f
C4589 _355_/a_891_413# 0 0.161052f
C4590 _355_/a_1059_315# 0 0.248849f
C4591 _355_/a_466_413# 0 0.133203f
C4592 _355_/a_634_159# 0 0.142309f
C4593 _355_/a_193_47# 0 0.284262f
C4594 _355_/a_27_47# 0 0.449511f
C4595 _039_ 0 0.259719f
C4596 _286_/a_27_53# 0 0.175308f
C4597 _286_/a_219_297# 0 0.137194f
C4598 _357__12/LO 0 0.165803f
C4599 _015_ 0 0.176197f
C4600 _339_/a_381_47# 0 0.016397f
C4601 _339_/a_891_413# 0 0.160892f
C4602 _339_/a_1062_300# 0 0.529662f
C4603 _339_/a_475_413# 0 0.137184f
C4604 _339_/a_634_183# 0 0.150209f
C4605 _339_/a_193_47# 0 0.271178f
C4606 _339_/a_27_47# 0 0.468295f
C4607 net13 0 0.11668f
C4608 _040_ 0 0.230406f
C4609 _287_/a_109_93# 0 0.160708f
C4610 _287_/a_215_53# 0 0.142592f
C4611 _356_/a_381_47# 0 0.015369f
C4612 _356_/a_891_413# 0 0.161052f
C4613 _356_/a_1059_315# 0 0.248849f
C4614 _356_/a_466_413# 0 0.133203f
C4615 _356_/a_634_159# 0 0.142309f
C4616 _356_/a_193_47# 0 0.284262f
C4617 _356_/a_27_47# 0 0.449511f
C4618 data[4] 0 0.361738f
C4619 input5/a_27_47# 0 0.207781f
C4620 _112_ 0 0.334037f
C4621 _211_/a_27_47# 0 0.174893f
C4622 clkbuf_2_1__f_clk/a_110_47# 0 1.73295f
C4623 _041_ 0 0.351716f
C4624 _000_ 0 0.230562f
C4625 net12 0 0.361147f
C4626 _357_/a_448_47# 0 0.013901f
C4627 _357_/a_1108_47# 0 0.13732f
C4628 _357_/a_1283_21# 0 0.389264f
C4629 _357_/a_543_47# 0 0.157869f
C4630 _357_/a_761_289# 0 0.120848f
C4631 _357_/a_193_47# 0 0.273213f
C4632 _357_/a_27_47# 0 0.495752f
C4633 data[3] 0 0.37078f
C4634 input4/a_27_47# 0 0.207781f
C4635 _113_ 0 0.151554f
C4636 _212_/a_80_21# 0 0.211154f
C4637 _042_ 0 0.105845f
C4638 _155_ 0 0.219748f
C4639 _289_/a_489_413# 0 0.025434f
C4640 _289_/a_226_47# 0 0.162324f
C4641 _289_/a_76_199# 0 0.140862f
C4642 data[2] 0 0.413922f
C4643 input3/a_27_47# 0 0.207781f
C4644 _052_ 0 0.521989f
C4645 _213_/a_109_93# 0 0.160708f
C4646 _213_/a_215_53# 0 0.142592f
C4647 data[1] 0 0.359718f
C4648 input2/a_27_47# 0 0.207781f
C4649 _127_ 0 0.146809f
C4650 _114_ 0 0.136883f
C4651 _111_ 0 0.159998f
C4652 _149_ 0 1.534441f
C4653 _214_/a_113_297# 0 0.034004f
C4654 data[0] 0 0.363997f
C4655 input1/a_27_47# 0 0.207781f
C4656 _053_ 0 1.334401f
C4657 _300_/a_27_47# 0 0.542977f
C4658 _075_ 0 0.114664f
C4659 net4 0 0.309257f
C4660 _073_ 0 0.212728f
C4661 _163_/a_27_47# 0 0.216317f
C4662 _301_/a_27_47# 0 0.28447f
C4663 r2r_out[7] 0 1.160314f
C4664 _116_ 0 0.1519f
C4665 _216_/a_59_75# 0 0.177062f
C4666 _129_ 0 0.089789f
C4667 _233_/a_80_21# 0 0.209712f
C4668 r2r_out[0] 0 2.317233f
C4669 _164_/a_215_47# 0 0.01011f
C4670 _164_/a_79_21# 0 0.225128f
C4671 _143_ 0 0.211409f
C4672 _250_/a_113_297# 0 0.034004f
C4673 _088_ 0 0.133974f
C4674 _181_/a_250_297# 0 0.02777f
C4675 _181_/a_93_21# 0 0.150721f
C4676 _217_/a_27_47# 0 0.174893f
C4677 _130_ 0 0.116032f
C4678 _128_ 0 0.110616f
C4679 _234_/a_113_297# 0 0.034004f
C4680 net1 0 0.368816f
C4681 _303_/a_113_297# 0 0.034004f
C4682 _071_ 0 0.159373f
C4683 _067_ 0 0.132817f
C4684 _070_ 0 0.104523f
C4685 _320_/a_80_21# 0 0.211154f
C4686 _144_ 0 0.131641f
C4687 _251_/a_27_47# 0 0.177187f
C4688 _090_ 0 0.12904f
C4689 _089_ 0 0.180024f
C4690 clknet_0_clk 0 1.846245f
C4691 clkbuf_2_0__f_clk/a_110_47# 0 1.73295f
C4692 net18 0 0.207903f
C4693 _131_ 0 0.112788f
C4694 _235_/a_113_297# 0 0.034004f
C4695 _011_ 0 0.175267f
C4696 net21 0 0.136787f
C4697 _321_/a_448_47# 0 0.032359f
C4698 _321_/a_222_93# 0 0.158855f
C4699 _321_/a_79_199# 0 0.148299f
C4700 _145_ 0 0.10199f
C4701 counter\[14\] 0 0.698601f
C4702 _252_/a_299_297# 0 0.034794f
C4703 _252_/a_81_21# 0 0.147141f
C4704 _091_ 0 0.132233f
C4705 _183_/a_59_75# 0 0.177062f
C4706 clk 0 0.459614f
C4707 clkbuf_0_clk/a_110_47# 0 1.73295f
C4708 _119_ 0 0.14516f
C4709 _118_ 0 0.140742f
C4710 _078_ 0 1.392431f
C4711 _117_ 0 0.667154f
C4712 _115_ 0 0.186166f
C4713 _219_/a_227_47# 0 0.030865f
C4714 _219_/a_77_199# 0 0.146762f
C4715 _236_/a_27_47# 0 0.174893f
C4716 _305_/a_27_47# 0 0.031143f
C4717 _048_ 0 0.292809f
C4718 _167_/a_27_47# 0 0.542977f
C4719 _253_/a_215_47# 0 0.01011f
C4720 _253_/a_79_21# 0 0.225128f
C4721 _092_ 0 0.151309f
C4722 net22 0 0.156584f
C4723 _184_/a_27_47# 0 0.031143f
C4724 _072_ 0 0.539387f
C4725 r2r_out[3] 0 0.796864f
C4726 _322_/a_27_47# 0 0.174893f
C4727 _009_ 0 0.140339f
C4728 _056_ 0 0.226233f
C4729 _058_ 0 0.158282f
C4730 _306_/a_113_297# 0 0.034004f
C4731 _133_ 0 0.537427f
C4732 _132_ 0 0.274153f
C4733 _237_/a_27_47# 0 0.177187f
C4734 _077_ 0 0.165882f
C4735 net5 0 0.418495f
C4736 _168_/a_505_21# 0 0.246761f
C4737 _168_/a_76_199# 0 0.139466f
C4738 net20 0 0.262933f
C4739 _185_/a_113_297# 0 0.034004f
C4740 _156_ 0 0.222705f
C4741 _271_/a_29_53# 0 0.180006f
C4742 _016_ 0 0.148404f
C4743 _340_/a_381_47# 0 0.016397f
C4744 _340_/a_891_413# 0 0.160892f
C4745 _340_/a_1062_300# 0 0.529662f
C4746 _340_/a_475_413# 0 0.137184f
C4747 _340_/a_634_183# 0 0.150209f
C4748 _340_/a_193_47# 0 0.271178f
C4749 _340_/a_27_47# 0 0.468295f
C4750 _307_/a_59_75# 0 0.177062f
C4751 _134_ 0 0.191206f
C4752 _035_ 0 0.373861f
C4753 _238_/a_227_47# 0 0.030865f
C4754 _238_/a_77_199# 0 0.146762f
C4755 _013_ 0 0.186012f
C4756 r2r_out[4] 0 1.242296f
C4757 _076_ 0 0.105215f
C4758 _079_ 0 0.107529f
C4759 _169_/a_240_47# 0 0.013847f
C4760 _169_/a_51_297# 0 0.206675f
C4761 _093_ 0 0.10698f
C4762 _186_/a_113_297# 0 0.034004f
C4763 _074_ 0 0.119032f
C4764 _324_/a_68_297# 0 0.153866f
C4765 _147_ 0 0.114846f
C4766 _255_/a_80_21# 0 0.211154f
C4767 _341_/a_381_47# 0 0.015369f
C4768 _341_/a_891_413# 0 0.161052f
C4769 _341_/a_1059_315# 0 0.248849f
C4770 _341_/a_466_413# 0 0.133203f
C4771 _341_/a_634_159# 0 0.142309f
C4772 _341_/a_193_47# 0 0.284262f
C4773 _341_/a_27_47# 0 0.449511f
C4774 _272_/a_215_297# 0 0.152836f
C4775 _272_/a_27_413# 0 0.171579f
C4776 _308_/a_27_47# 0 0.542977f
C4777 _017_ 0 0.166374f
C4778 net19 0 0.149634f
C4779 _060_ 0 1.243661f
C4780 _187_/a_297_47# 0 0.034813f
C4781 _187_/a_79_21# 0 0.158207f
C4782 _032_ 0 0.191735f
C4783 _146_ 0 0.11411f
C4784 _256_/a_81_21# 0 0.214691f
C4785 _325_/a_381_47# 0 0.015369f
C4786 _325_/a_891_413# 0 0.161052f
C4787 _325_/a_1059_315# 0 0.248849f
C4788 _325_/a_466_413# 0 0.133203f
C4789 _325_/a_634_159# 0 0.142309f
C4790 _325_/a_193_47# 0 0.284262f
C4791 _325_/a_27_47# 0 0.449511f
C4792 counter\[1\] 0 0.691615f
C4793 _342_/a_381_47# 0 0.015369f
C4794 _342_/a_891_413# 0 0.161052f
C4795 _342_/a_1059_315# 0 0.248849f
C4796 _342_/a_466_413# 0 0.133203f
C4797 _342_/a_634_159# 0 0.142309f
C4798 _342_/a_193_47# 0 0.284262f
C4799 _342_/a_27_47# 0 0.449511f
C4800 _273_/a_109_93# 0 0.160708f
C4801 _273_/a_215_53# 0 0.142592f
C4802 _290_/a_207_413# 0 0.137402f
C4803 _290_/a_27_413# 0 0.196502f
C4804 _055_ 0 0.209131f
C4805 _309_/a_27_47# 0 0.031143f
C4806 _188_/a_27_47# 0 0.28447f
C4807 _326_/a_381_47# 0 0.015369f
C4808 _326_/a_891_413# 0 0.161052f
C4809 _326_/a_1059_315# 0 0.248849f
C4810 _326_/a_466_413# 0 0.133203f
C4811 _326_/a_634_159# 0 0.142309f
C4812 _326_/a_193_47# 0 0.284262f
C4813 _326_/a_27_47# 0 0.449511f
C4814 net11 0 0.273023f
C4815 _343_/a_381_47# 0 0.015369f
C4816 _343_/a_891_413# 0 0.161052f
C4817 _343_/a_1059_315# 0 0.248849f
C4818 _343_/a_466_413# 0 0.133203f
C4819 _343_/a_634_159# 0 0.142309f
C4820 _343_/a_193_47# 0 0.284262f
C4821 _343_/a_27_47# 0 0.449511f
C4822 _157_ 0 0.232165f
C4823 _274_/a_215_297# 0 0.152836f
C4824 _274_/a_27_413# 0 0.171579f
C4825 _044_ 0 0.121697f
C4826 divider\[3\] 0 0.358831f
C4827 _291_/a_27_47# 0 0.216317f
C4828 hold10/a_391_47# 0 0.127705f
C4829 hold10/a_285_47# 0 0.29867f
C4830 hold10/a_49_47# 0 0.306903f
C4831 _189_/a_285_47# 0 0.017425f
C4832 _189_/a_47_47# 0 0.199276f
C4833 _258_/a_27_47# 0 0.28447f
C4834 _327_/a_381_47# 0 0.015369f
C4835 _327_/a_891_413# 0 0.161052f
C4836 _327_/a_1059_315# 0 0.248849f
C4837 _327_/a_466_413# 0 0.133203f
C4838 _327_/a_634_159# 0 0.142309f
C4839 _327_/a_193_47# 0 0.284262f
C4840 _327_/a_27_47# 0 0.449511f
C4841 _344_/a_381_47# 0 0.015369f
C4842 _344_/a_891_413# 0 0.161052f
C4843 _344_/a_1059_315# 0 0.248849f
C4844 _344_/a_466_413# 0 0.133203f
C4845 _344_/a_634_159# 0 0.142309f
C4846 _344_/a_193_47# 0 0.284262f
C4847 _344_/a_27_47# 0 0.449511f
C4848 _158_ 0 0.294234f
C4849 net10 0 0.999061f
C4850 rst 0 0.938187f
C4851 _275_/a_109_93# 0 0.160708f
C4852 _275_/a_215_53# 0 0.142592f
C4853 _036_ 0 0.144652f
C4854 _292_/a_516_297# 0 0.035006f
C4855 _292_/a_85_193# 0 0.166604f
C4856 _328_/a_381_47# 0 0.015369f
C4857 _328_/a_891_413# 0 0.161052f
C4858 _328_/a_1059_315# 0 0.248849f
C4859 _328_/a_466_413# 0 0.133203f
C4860 _328_/a_634_159# 0 0.142309f
C4861 _328_/a_193_47# 0 0.284262f
C4862 _328_/a_27_47# 0 0.449511f
C4863 _259_/a_27_47# 0 0.542977f
C4864 counter\[4\] 0 0.80553f
C4865 _021_ 0 0.17623f
C4866 clknet_2_1__leaf_clk 0 1.550415f
C4867 _345_/a_381_47# 0 0.015369f
C4868 _345_/a_891_413# 0 0.161052f
C4869 _345_/a_1059_315# 0 0.248849f
C4870 _345_/a_466_413# 0 0.133203f
C4871 _345_/a_634_159# 0 0.142309f
C4872 _345_/a_193_47# 0 0.284262f
C4873 _345_/a_27_47# 0 0.449511f
C4874 net8 0 0.322867f
C4875 _276_/a_215_297# 0 0.152836f
C4876 _276_/a_27_413# 0 0.171579f
C4877 _329_/a_381_47# 0 0.015369f
C4878 _329_/a_891_413# 0 0.161052f
C4879 _329_/a_1059_315# 0 0.248849f
C4880 _329_/a_466_413# 0 0.133203f
C4881 _329_/a_634_159# 0 0.142309f
C4882 _329_/a_193_47# 0 0.284262f
C4883 _329_/a_27_47# 0 0.449511f
C4884 _200_/a_227_47# 0 0.030865f
C4885 _200_/a_77_199# 0 0.146762f
C4886 _159_ 0 0.283177f
C4887 counter\[5\] 0 0.645322f
C4888 clknet_2_0__leaf_clk 0 1.259837f
C4889 _346_/a_381_47# 0 0.015369f
C4890 _346_/a_891_413# 0 0.161052f
C4891 _346_/a_1059_315# 0 0.248849f
C4892 _346_/a_466_413# 0 0.133203f
C4893 _346_/a_634_159# 0 0.142309f
C4894 _346_/a_193_47# 0 0.284262f
C4895 _346_/a_27_47# 0 0.449511f
C4896 divider\[5\] 0 0.461407f
C4897 divider\[4\] 0 0.550471f
C4898 _294_/a_215_47# 0 0.035725f
C4899 _294_/a_78_199# 0 0.15408f
.ends

.subckt sky130_fd_pr__res_high_po_0p35_3KK54B a_n35_n4432# a_n35_4000# a_n165_n4562#
X0 a_n35_4000# a_n35_n4432# a_n165_n4562# sky130_fd_pr__res_high_po_0p35 l=40
C0 a_n35_n4432# a_n165_n4562# 0.597536f
C1 a_n35_4000# a_n165_n4562# 0.597536f
.ends

.subckt sky130_fd_pr__res_high_po_0p35_QPS5FG a_n165_n2562# a_n35_n2432# a_n35_2000#
X0 a_n35_2000# a_n35_n2432# a_n165_n2562# sky130_fd_pr__res_high_po_0p35 l=20
C0 a_n35_n2432# a_n165_n2562# 0.597536f
C1 a_n35_2000# a_n165_n2562# 0.597536f
.ends

.subckt r2r b0 b1 b2 b3 b4 b5 b6 b7 GND m1_n1840_11060# VSUBS out
XXR1 m1_n1840_11060# b0 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR10 VSUBS m1_n1040_2660# m1_n440_7180# sky130_fd_pr__res_high_po_0p35_QPS5FG
XXR2 m1_n1040_2660# b1 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR11 VSUBS m1_160_2660# m1_n440_7180# sky130_fd_pr__res_high_po_0p35_QPS5FG
XXR3 m1_n440_7180# b2 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR5 m1_760_7180# b4 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR12 VSUBS m1_160_2660# m1_760_7180# sky130_fd_pr__res_high_po_0p35_QPS5FG
XXR4 m1_160_2660# b3 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR14 VSUBS m1_1360_2660# m1_1960_7180# sky130_fd_pr__res_high_po_0p35_QPS5FG
XXR6 m1_1360_2660# b5 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR13 VSUBS m1_1360_2660# m1_760_7180# sky130_fd_pr__res_high_po_0p35_QPS5FG
XXR15 VSUBS out m1_1960_7180# sky130_fd_pr__res_high_po_0p35_QPS5FG
XXR7 m1_1960_7180# b6 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR8 out b7 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR16 GND m1_n1840_11060# VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR9 VSUBS m1_n1040_2660# m1_n1840_11060# sky130_fd_pr__res_high_po_0p35_QPS5FG
C0 b2 b1 0.098267f
C1 m1_160_2660# m1_760_7180# 0.131455f
C2 out m1_1360_2660# 0.151802f
C3 m1_n440_7180# m1_160_2660# 0.209321f
C4 m1_160_2660# m1_n1040_2660# 0.182372f
C5 m1_1360_2660# m1_160_2660# 0.182372f
C6 b2 b3 0.098267f
C7 m1_1360_2660# m1_1960_7180# 0.131485f
C8 out m1_1960_7180# 0.106769f
C9 b6 b7 0.098267f
C10 b5 b4 0.098267f
C11 m1_n1040_2660# GND 0.023658f
C12 m1_n1040_2660# m1_n1840_11060# 0.20932f
C13 b4 b3 0.098267f
C14 m1_1360_2660# m1_760_7180# 0.209322f
C15 b5 b6 0.098267f
C16 b1 b0 0.098267f
C17 m1_n440_7180# m1_n1040_2660# 0.131455f
C18 m1_n1040_2660# VSUBS 4.058431f
C19 GND VSUBS 0.991775f
C20 b7 VSUBS 0.971434f
C21 b6 VSUBS 0.866416f
C22 out VSUBS 4.202785f
C23 m1_1360_2660# VSUBS 3.909692f
C24 b5 VSUBS 0.866416f
C25 m1_1960_7180# VSUBS 2.022547f
C26 b3 VSUBS 0.866416f
C27 m1_760_7180# VSUBS 1.959661f
C28 b4 VSUBS 0.866416f
C29 b2 VSUBS 0.866416f
C30 m1_160_2660# VSUBS 3.875238f
C31 b1 VSUBS 0.866416f
C32 m1_n440_7180# VSUBS 1.959661f
C33 m1_n1840_11060# VSUBS 3.79668f
C34 b0 VSUBS 0.971437f
.ends

.subckt tt_um_mattvenn_r2r_dac clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VPWR VGND
Xr2r_dac_control_0 clk ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6]
+ ui_in[7] uio_in[0] uio_in[1] rst_n r2r_0/b0 r2r_0/b1 r2r_0/b2 r2r_0/b3 r2r_0/b4
+ r2r_0/b5 r2r_0/b6 r2r_0/b7 VPWR VGND r2r_dac_control
Xr2r_0 r2r_0/b0 r2r_0/b1 r2r_0/b2 r2r_0/b3 r2r_0/b4 r2r_0/b5 r2r_0/b6 r2r_0/b7 VGND
+ r2r_0/m1_n1840_11060# VGND ua[0] r2r
C0 uio_out[5] uio_out[6] 0.023797f
C1 ui_in[7] ui_in[6] 5.41126f
C2 ui_in[3] ui_in[2] 5.310389f
C3 ui_in[1] ui_in[2] 4.496709f
C4 uo_out[4] uo_out[5] 0.023797f
C5 r2r_0/b2 r2r_0/b3 0.287249f
C6 uio_out[5] uio_out[4] 0.023797f
C7 uio_out[0] uo_out[7] 0.023797f
C8 uio_in[0] uio_in[1] 6.209905f
C9 VGND clk 0.022177f
C10 r2r_0/b1 VGND 0.013869f
C11 ui_in[5] ui_in[6] 4.918385f
C12 uio_out[3] uio_out[4] 0.023797f
C13 uio_in[6] uio_in[5] 0.023797f
C14 uio_out[3] uio_out[2] 0.023797f
C15 uo_out[4] uo_out[3] 0.023797f
C16 uo_out[1] uo_out[2] 0.023797f
C17 VGND r2r_0/b0 0.010392f
C18 VGND VPWR 9.442356f
C19 VPWR ui_in[0] 0.03106f
C20 r2r_0/b1 r2r_0/b0 0.123983f
C21 uo_out[3] uo_out[2] 0.023797f
C22 VGND uio_oe[3] 0.016443f
C23 uio_in[3] uio_in[4] 0.023797f
C24 r2r_0/b1 r2r_0/b2 0.280483f
C25 r2r_0/b5 r2r_0/b6 1.032367f
C26 uo_out[6] uo_out[7] 0.023797f
C27 ui_in[3] ui_in[4] 4.3829f
C28 uio_in[1] uio_in[2] 0.024975f
C29 ui_in[0] rst_n 4.713152f
C30 clk rst_n 4.541323f
C31 ui_in[7] uio_in[0] 6.181085f
C32 uio_in[4] uio_in[5] 0.023797f
C33 VPWR rst_n 0.020143f
C34 r2r_0/b7 r2r_0/b6 1.281466f
C35 uo_out[6] uo_out[5] 0.023797f
C36 clk ena 0.023816f
C37 VGND uio_in[1] 0.178487f
C38 VGND r2r_0/m1_n1840_11060# 0.047088f
C39 r2r_0/b5 r2r_0/b4 0.780769f
C40 uio_in[3] uio_in[2] 0.023797f
C41 ui_in[5] ui_in[4] 4.521664f
C42 uio_oe[5] uio_oe[4] 0.023797f
C43 uio_out[7] uio_out[6] 0.023797f
C44 VGND uio_out[7] 0.023797f
C45 uo_out[0] uo_out[1] 0.023797f
C46 VGND uio_in[0] 0.015812f
C47 ui_in[0] ui_in[1] 4.916256f
C48 VGND uio_oe[2] 0.040241f
C49 uio_out[0] uio_out[1] 0.023797f
C50 uo_out[0] uio_in[7] 0.023797f
C51 VPWR ua[7] 0.010285f
C52 uio_oe[6] uio_oe[7] 0.023797f
C53 VPWR ui_in[1] 0.011936f
C54 uio_in[6] uio_in[7] 0.023797f
C55 uio_oe[2] uio_oe[3] 0.023797f
C56 r2r_0/b7 clk 0.352877f
C57 uio_oe[5] uio_oe[6] 0.023797f
C58 uio_out[1] uio_out[2] 0.023797f
C59 r2r_0/b3 r2r_0/b4 0.528153f
C60 uio_oe[4] uio_oe[3] 0.023797f
C61 ua[1] 0 0.122428f
C62 ua[2] 0 0.122428f
C63 ua[3] 0 0.122428f
C64 ua[4] 0 0.122428f
C65 ua[5] 0 0.122428f
C66 ua[6] 0 0.122428f
C67 ua[7] 0 0.111009f
C68 ena 0 0.073288f
C69 uio_in[2] 0 0.047383f
C70 uio_in[3] 0 0.047383f
C71 uio_in[4] 0 0.047383f
C72 uio_in[5] 0 0.047383f
C73 uio_in[6] 0 0.047383f
C74 uio_in[7] 0 0.047383f
C75 uo_out[0] 0 0.047383f
C76 uo_out[1] 0 0.047383f
C77 uo_out[2] 0 0.047383f
C78 uo_out[3] 0 0.047383f
C79 uo_out[4] 0 0.047383f
C80 uo_out[5] 0 0.047383f
C81 uo_out[6] 0 0.047383f
C82 uo_out[7] 0 0.047383f
C83 uio_out[0] 0 0.047383f
C84 uio_out[1] 0 0.047383f
C85 uio_out[2] 0 0.047354f
C86 uio_out[3] 0 0.047516f
C87 uio_out[4] 0 0.047679f
C88 uio_out[5] 0 0.047679f
C89 uio_out[6] 0 0.047878f
C90 uio_out[7] 0 0.047878f
C91 uio_oe[2] 0 0.03903f
C92 uio_oe[3] 0 0.03903f
C93 uio_oe[4] 0 0.043789f
C94 uio_oe[5] 0 0.043789f
C95 uio_oe[6] 0 0.0487f
C96 uio_oe[7] 0 0.073297f
C97 r2r_0/m1_n1040_2660# 0 3.629388f
C98 ua[0] 0 14.659142f
C99 r2r_0/m1_1360_2660# 0 3.477601f
C100 r2r_0/m1_1960_7180# 0 1.900238f
C101 r2r_0/m1_760_7180# 0 1.838729f
C102 r2r_0/m1_160_2660# 0 3.443148f
C103 r2r_0/m1_n440_7180# 0 1.838729f
C104 r2r_0/m1_n1840_11060# 0 3.562639f
C105 r2r_dac_control_0/_020_ 0 0.139788f
C106 r2r_dac_control_0/_104_ 0 0.143482f
C107 r2r_dac_control_0/counter\[6\] 0 0.511237f
C108 r2r_dac_control_0/_023_ 0 0.172897f
C109 r2r_dac_control_0/_347_/a_381_47# 0 0.015369f
C110 r2r_dac_control_0/_347_/a_891_413# 0 0.161052f
C111 r2r_dac_control_0/_347_/a_1059_315# 0 0.248849f
C112 r2r_dac_control_0/_347_/a_466_413# 0 0.133203f
C113 r2r_dac_control_0/_347_/a_634_159# 0 0.142309f
C114 r2r_dac_control_0/_347_/a_193_47# 0 0.284262f
C115 r2r_dac_control_0/_347_/a_27_47# 0 0.449511f
C116 VPWR 0 0.507816p
C117 VGND 0 0.172048p
C118 r2r_dac_control_0/_160_ 0 0.129815f
C119 r2r_dac_control_0/divider\[1\] 0 0.412489f
C120 r2r_dac_control_0/_278_/a_27_53# 0 0.175308f
C121 r2r_dac_control_0/_278_/a_219_297# 0 0.137194f
C122 r2r_dac_control_0/_105_ 0 0.124266f
C123 r2r_dac_control_0/net14 0 0.119432f
C124 r2r_dac_control_0/counter\[7\] 0 0.594844f
C125 r2r_dac_control_0/_024_ 0 0.184261f
C126 r2r_dac_control_0/_348_/a_381_47# 0 0.015369f
C127 r2r_dac_control_0/_348_/a_891_413# 0 0.161052f
C128 r2r_dac_control_0/_348_/a_1059_315# 0 0.248849f
C129 r2r_dac_control_0/_348_/a_466_413# 0 0.133203f
C130 r2r_dac_control_0/_348_/a_634_159# 0 0.142309f
C131 r2r_dac_control_0/_348_/a_193_47# 0 0.284262f
C132 r2r_dac_control_0/_348_/a_27_47# 0 0.449511f
C133 r2r_dac_control_0/divider\[0\] 0 0.284172f
C134 r2r_dac_control_0/_279_/a_207_413# 0 0.137402f
C135 r2r_dac_control_0/_279_/a_27_413# 0 0.196502f
C136 r2r_dac_control_0/_049_ 0 0.195114f
C137 r2r_dac_control_0/_296_/a_27_53# 0 0.175308f
C138 r2r_dac_control_0/_296_/a_219_297# 0 0.137194f
C139 r2r_dac_control_0/_349_/a_381_47# 0 0.015369f
C140 r2r_dac_control_0/_349_/a_891_413# 0 0.161052f
C141 r2r_dac_control_0/_349_/a_1059_315# 0 0.248849f
C142 r2r_dac_control_0/_349_/a_466_413# 0 0.133203f
C143 r2r_dac_control_0/_349_/a_634_159# 0 0.142309f
C144 r2r_dac_control_0/_349_/a_193_47# 0 0.284262f
C145 r2r_dac_control_0/_349_/a_27_47# 0 0.449511f
C146 r2r_dac_control_0/_050_ 0 0.147091f
C147 r2r_dac_control_0/_297_/a_215_47# 0 0.01011f
C148 r2r_dac_control_0/_297_/a_79_21# 0 0.225128f
C149 r2r_dac_control_0/_101_ 0 0.916798f
C150 r2r_dac_control_0/_120_ 0 0.14294f
C151 r2r_dac_control_0/_221_/a_68_297# 0 0.153866f
C152 r2r_dac_control_0/_043_ 0 0.242838f
C153 r2r_dac_control_0/_047_ 0 0.088296f
C154 r2r_dac_control_0/_298_/a_253_47# 0 0.011031f
C155 r2r_dac_control_0/_298_/a_103_199# 0 0.196442f
C156 r2r_dac_control_0/_108_ 0 0.133143f
C157 r2r_dac_control_0/_106_ 0 0.142206f
C158 r2r_dac_control_0/_205_/a_109_93# 0 0.160708f
C159 r2r_dac_control_0/_205_/a_215_53# 0 0.142592f
C160 r2r_dac_control_0/_121_ 0 0.275415f
C161 r2r_dac_control_0/_045_ 0 0.263731f
C162 r2r_dac_control_0/_051_ 0 0.296787f
C163 r2r_dac_control_0/_080_ 0 0.119111f
C164 r2r_0/b5 0 6.00686f
C165 r2r_dac_control_0/_170_/a_299_297# 0 0.034794f
C166 r2r_dac_control_0/_170_/a_81_21# 0 0.147141f
C167 r2r_dac_control_0/_206_/a_113_297# 0 0.034004f
C168 r2r_dac_control_0/_054_ 0 1.597855f
C169 r2r_dac_control_0/_059_ 0 0.350294f
C170 r2r_dac_control_0/_223_/a_250_297# 0 0.02777f
C171 r2r_dac_control_0/_223_/a_93_21# 0 0.150721f
C172 r2r_dac_control_0/_135_ 0 0.110228f
C173 r2r_dac_control_0/_240_/a_68_297# 0 0.153866f
C174 r2r_dac_control_0/_171_/a_27_47# 0 0.177187f
C175 r2r_dac_control_0/_109_ 0 0.104062f
C176 r2r_dac_control_0/_107_ 0 0.345335f
C177 r2r_dac_control_0/_207_/a_35_297# 0 0.254573f
C178 r2r_dac_control_0/hold9/a_391_47# 0 0.127705f
C179 r2r_dac_control_0/hold9/a_285_47# 0 0.29867f
C180 r2r_dac_control_0/hold9/a_49_47# 0 0.306903f
C181 r2r_dac_control_0/_122_ 0 0.14449f
C182 r2r_dac_control_0/_057_ 0 1.413733f
C183 r2r_dac_control_0/_224_/a_59_75# 0 0.177062f
C184 r2r_dac_control_0/_136_ 0 0.27487f
C185 r2r_dac_control_0/_241_/a_59_75# 0 0.177062f
C186 r2r_dac_control_0/_082_ 0 0.106064f
C187 r2r_dac_control_0/_081_ 0 0.474985f
C188 r2r_dac_control_0/clkbuf_2_3__f_clk/a_110_47# 0 1.73295f
C189 r2r_dac_control_0/_094_ 0 1.195606f
C190 r2r_dac_control_0/_066_ 0 1.46872f
C191 r2r_dac_control_0/_208_/a_489_47# 0 0.037211f
C192 r2r_dac_control_0/_208_/a_206_369# 0 0.153769f
C193 r2r_dac_control_0/_208_/a_76_199# 0 0.136541f
C194 r2r_dac_control_0/hold8/a_391_47# 0 0.127705f
C195 r2r_dac_control_0/hold8/a_285_47# 0 0.29867f
C196 r2r_dac_control_0/hold8/a_49_47# 0 0.306903f
C197 r2r_dac_control_0/_025_ 0 0.180417f
C198 r2r_dac_control_0/_123_ 0 0.170328f
C199 r2r_dac_control_0/_225_/a_75_212# 0 0.210264f
C200 r2r_dac_control_0/net2 0 0.285409f
C201 r2r_dac_control_0/_062_ 0 0.111631f
C202 r2r_dac_control_0/_311_/a_27_297# 0 0.190287f
C203 r2r_dac_control_0/_083_ 0 0.132825f
C204 r2r_dac_control_0/net6 0 0.371254f
C205 r2r_dac_control_0/_173_/a_27_47# 0 0.216317f
C206 r2r_dac_control_0/_095_ 0 0.141562f
C207 r2r_dac_control_0/_190_/a_489_47# 0 0.037211f
C208 r2r_dac_control_0/_190_/a_206_369# 0 0.153769f
C209 r2r_dac_control_0/_190_/a_76_199# 0 0.136541f
C210 r2r_dac_control_0/_022_ 0 0.190239f
C211 r2r_dac_control_0/_065_ 0 1.814524f
C212 r2r_dac_control_0/_110_ 0 0.200614f
C213 r2r_dac_control_0/hold7/a_391_47# 0 0.127705f
C214 r2r_dac_control_0/hold7/a_285_47# 0 0.29867f
C215 r2r_dac_control_0/hold7/a_49_47# 0 0.306903f
C216 r2r_dac_control_0/_124_ 0 0.248471f
C217 r2r_dac_control_0/counter\[9\] 0 0.84899f
C218 r2r_dac_control_0/_138_ 0 0.14067f
C219 r2r_dac_control_0/_137_ 0 0.102851f
C220 r2r_dac_control_0/_243_/a_250_297# 0 0.02777f
C221 r2r_dac_control_0/_243_/a_93_21# 0 0.150721f
C222 r2r_dac_control_0/_063_ 0 0.161343f
C223 r2r_dac_control_0/_014_ 0 0.165446f
C224 r2r_dac_control_0/_174_/a_215_47# 0 0.01011f
C225 r2r_dac_control_0/_174_/a_79_21# 0 0.225128f
C226 r2r_dac_control_0/_018_ 0 0.175898f
C227 r2r_dac_control_0/_096_ 0 0.212547f
C228 r2r_dac_control_0/_260_/a_109_93# 0 0.160708f
C229 r2r_dac_control_0/_260_/a_215_53# 0 0.142592f
C230 r2r_dac_control_0/hold6/a_391_47# 0 0.127705f
C231 r2r_dac_control_0/hold6/a_285_47# 0 0.29867f
C232 r2r_dac_control_0/hold6/a_49_47# 0 0.306903f
C233 r2r_dac_control_0/_227_/a_59_75# 0 0.177062f
C234 r2r_dac_control_0/_139_ 0 0.137918f
C235 r2r_dac_control_0/_244_/a_59_75# 0 0.177062f
C236 r2r_dac_control_0/_313_/a_27_47# 0 0.542977f
C237 r2r_dac_control_0/_084_ 0 0.2838f
C238 r2r_0/b6 0 6.834352f
C239 r2r_dac_control_0/_097_ 0 0.335599f
C240 r2r_dac_control_0/counter\[0\] 0 0.951161f
C241 r2r_dac_control_0/counter\[2\] 0 0.576308f
C242 r2r_dac_control_0/_192_/a_27_47# 0 0.177187f
C243 r2r_dac_control_0/_006_ 0 0.180268f
C244 r2r_dac_control_0/_330_/a_381_47# 0 0.015369f
C245 r2r_dac_control_0/_330_/a_891_413# 0 0.161052f
C246 r2r_dac_control_0/_330_/a_1059_315# 0 0.248849f
C247 r2r_dac_control_0/_330_/a_466_413# 0 0.133203f
C248 r2r_dac_control_0/_330_/a_634_159# 0 0.142309f
C249 r2r_dac_control_0/_330_/a_193_47# 0 0.284262f
C250 r2r_dac_control_0/_330_/a_27_47# 0 0.449511f
C251 r2r_dac_control_0/_001_ 0 0.158742f
C252 r2r_dac_control_0/_150_ 0 0.184778f
C253 r2r_dac_control_0/_261_/a_215_297# 0 0.152836f
C254 r2r_dac_control_0/_261_/a_27_413# 0 0.171579f
C255 r2r_dac_control_0/net17 0 0.217366f
C256 r2r_dac_control_0/hold5/a_391_47# 0 0.127705f
C257 r2r_dac_control_0/hold5/a_285_47# 0 0.29867f
C258 r2r_dac_control_0/hold5/a_49_47# 0 0.306903f
C259 r2r_dac_control_0/counter\[8\] 0 0.733786f
C260 r2r_dac_control_0/_228_/a_27_47# 0 0.177187f
C261 r2r_dac_control_0/_029_ 0 0.194126f
C262 r2r_dac_control_0/_245_/a_75_212# 0 0.210264f
C263 r2r_dac_control_0/_064_ 0 0.111564f
C264 r2r_dac_control_0/_061_ 0 0.121096f
C265 r2r_dac_control_0/_314_/a_113_297# 0 0.034004f
C266 r2r_dac_control_0/_176_/a_68_297# 0 0.153866f
C267 r2r_dac_control_0/_193_/a_113_297# 0 0.034004f
C268 r2r_dac_control_0/_151_ 0 0.217983f
C269 r2r_dac_control_0/_262_/a_109_93# 0 0.160708f
C270 r2r_dac_control_0/_262_/a_215_53# 0 0.142592f
C271 r2r_dac_control_0/_007_ 0 0.164432f
C272 r2r_dac_control_0/_331_/a_381_47# 0 0.015369f
C273 r2r_dac_control_0/_331_/a_891_413# 0 0.161052f
C274 r2r_dac_control_0/_331_/a_1059_315# 0 0.248849f
C275 r2r_dac_control_0/_331_/a_466_413# 0 0.133203f
C276 r2r_dac_control_0/_331_/a_634_159# 0 0.142309f
C277 r2r_dac_control_0/_331_/a_193_47# 0 0.284262f
C278 r2r_dac_control_0/_331_/a_27_47# 0 0.449511f
C279 r2r_dac_control_0/hold4/a_391_47# 0 0.127705f
C280 r2r_dac_control_0/hold4/a_285_47# 0 0.29867f
C281 r2r_dac_control_0/hold4/a_49_47# 0 0.306903f
C282 r2r_dac_control_0/_126_ 0 0.471049f
C283 r2r_dac_control_0/_125_ 0 0.103379f
C284 r2r_dac_control_0/_229_/a_227_47# 0 0.030865f
C285 r2r_dac_control_0/_229_/a_77_199# 0 0.146762f
C286 r2r_dac_control_0/_140_ 0 0.115252f
C287 r2r_dac_control_0/counter\[12\] 0 0.850806f
C288 r2r_dac_control_0/counter\[13\] 0 1.031976f
C289 r2r_dac_control_0/_246_/a_113_297# 0 0.034004f
C290 r2r_dac_control_0/_315_/a_27_47# 0 0.542977f
C291 r2r_dac_control_0/_086_ 0 0.13159f
C292 r2r_dac_control_0/net7 0 0.367186f
C293 r2r_dac_control_0/_177_/a_59_75# 0 0.177062f
C294 r2r_dac_control_0/_008_ 0 0.166318f
C295 r2r_dac_control_0/_332_/a_381_47# 0 0.015369f
C296 r2r_dac_control_0/_332_/a_891_413# 0 0.161052f
C297 r2r_dac_control_0/_332_/a_1059_315# 0 0.248849f
C298 r2r_dac_control_0/_332_/a_466_413# 0 0.133203f
C299 r2r_dac_control_0/_332_/a_634_159# 0 0.142309f
C300 r2r_dac_control_0/_332_/a_193_47# 0 0.284262f
C301 r2r_dac_control_0/_332_/a_27_47# 0 0.449511f
C302 r2r_dac_control_0/_002_ 0 0.154364f
C303 r2r_dac_control_0/_263_/a_215_297# 0 0.152836f
C304 r2r_dac_control_0/_263_/a_27_413# 0 0.171579f
C305 r2r_dac_control_0/_280_/a_207_413# 0 0.137402f
C306 r2r_dac_control_0/_280_/a_27_413# 0 0.196502f
C307 r2r_dac_control_0/net15 0 0.143914f
C308 r2r_dac_control_0/hold3/a_391_47# 0 0.127705f
C309 r2r_dac_control_0/hold3/a_285_47# 0 0.29867f
C310 r2r_dac_control_0/hold3/a_49_47# 0 0.306903f
C311 r2r_dac_control_0/_087_ 0 0.115233f
C312 r2r_dac_control_0/_085_ 0 0.131682f
C313 r2r_dac_control_0/_178_/a_75_199# 0 0.20459f
C314 r2r_dac_control_0/_141_ 0 0.372285f
C315 r2r_dac_control_0/_247_/a_27_47# 0 0.177187f
C316 r2r_dac_control_0/net3 0 0.308777f
C317 r2r_dac_control_0/_333_/a_381_47# 0 0.016397f
C318 r2r_dac_control_0/_333_/a_891_413# 0 0.160892f
C319 r2r_dac_control_0/_333_/a_1062_300# 0 0.529662f
C320 r2r_dac_control_0/_333_/a_475_413# 0 0.137184f
C321 r2r_dac_control_0/_333_/a_634_183# 0 0.150209f
C322 r2r_dac_control_0/_333_/a_193_47# 0 0.271178f
C323 r2r_dac_control_0/_333_/a_27_47# 0 0.468295f
C324 r2r_dac_control_0/_099_ 0 0.143522f
C325 r2r_dac_control_0/_098_ 0 0.092047f
C326 r2r_dac_control_0/_195_/a_227_47# 0 0.030865f
C327 r2r_dac_control_0/_195_/a_77_199# 0 0.146762f
C328 r2r_dac_control_0/_264_/a_109_93# 0 0.160708f
C329 r2r_dac_control_0/_264_/a_215_53# 0 0.142592f
C330 r2r_dac_control_0/_026_ 0 0.206154f
C331 r2r_dac_control_0/_350_/a_381_47# 0 0.015369f
C332 r2r_dac_control_0/_350_/a_891_413# 0 0.161052f
C333 r2r_dac_control_0/_350_/a_1059_315# 0 0.248849f
C334 r2r_dac_control_0/_350_/a_466_413# 0 0.133203f
C335 r2r_dac_control_0/_350_/a_634_159# 0 0.142309f
C336 r2r_dac_control_0/_350_/a_193_47# 0 0.284262f
C337 r2r_dac_control_0/_350_/a_27_47# 0 0.449511f
C338 r2r_dac_control_0/_034_ 0 0.149276f
C339 r2r_dac_control_0/divider\[2\] 0 0.471944f
C340 r2r_dac_control_0/_161_ 0 0.121029f
C341 r2r_dac_control_0/_033_ 0 0.122585f
C342 r2r_dac_control_0/_281_/a_27_47# 0 0.216317f
C343 r2r_dac_control_0/hold2/a_391_47# 0 0.127705f
C344 r2r_dac_control_0/hold2/a_285_47# 0 0.29867f
C345 r2r_dac_control_0/hold2/a_49_47# 0 0.306903f
C346 r2r_dac_control_0/clkbuf_2_2__f_clk/a_110_47# 0 1.73295f
C347 r2r_dac_control_0/_068_ 0 0.102682f
C348 r2r_0/b2 0 4.163335f
C349 r2r_dac_control_0/_317_/a_113_297# 0 0.034004f
C350 r2r_dac_control_0/_046_ 0 0.267328f
C351 r2r_dac_control_0/_248_/a_227_47# 0 0.030865f
C352 r2r_dac_control_0/_248_/a_77_199# 0 0.146762f
C353 r2r_dac_control_0/_179_/a_215_47# 0 0.01011f
C354 r2r_dac_control_0/_179_/a_79_21# 0 0.225128f
C355 r2r_dac_control_0/_019_ 0 0.166532f
C356 r2r_dac_control_0/_100_ 0 0.138217f
C357 r2r_dac_control_0/_003_ 0 0.16738f
C358 r2r_dac_control_0/_152_ 0 0.266852f
C359 r2r_dac_control_0/_265_/a_215_297# 0 0.152836f
C360 r2r_dac_control_0/_265_/a_27_413# 0 0.171579f
C361 r2r_0/b1 0 4.018358f
C362 r2r_dac_control_0/_010_ 0 0.133868f
C363 r2r_dac_control_0/_334_/a_381_47# 0 0.016397f
C364 r2r_dac_control_0/_334_/a_891_413# 0 0.160892f
C365 r2r_dac_control_0/_334_/a_1062_300# 0 0.529662f
C366 r2r_dac_control_0/_334_/a_475_413# 0 0.137184f
C367 r2r_dac_control_0/_334_/a_634_183# 0 0.150209f
C368 r2r_dac_control_0/_334_/a_193_47# 0 0.271178f
C369 r2r_dac_control_0/_334_/a_27_47# 0 0.468295f
C370 r2r_dac_control_0/counter\[10\] 0 0.882194f
C371 r2r_dac_control_0/_027_ 0 0.144188f
C372 r2r_dac_control_0/_351_/a_381_47# 0 0.015369f
C373 r2r_dac_control_0/_351_/a_891_413# 0 0.161052f
C374 r2r_dac_control_0/_351_/a_1059_315# 0 0.248849f
C375 r2r_dac_control_0/_351_/a_466_413# 0 0.133203f
C376 r2r_dac_control_0/_351_/a_634_159# 0 0.142309f
C377 r2r_dac_control_0/_351_/a_193_47# 0 0.284262f
C378 r2r_dac_control_0/_351_/a_27_47# 0 0.449511f
C379 r2r_dac_control_0/hold1/a_391_47# 0 0.127705f
C380 r2r_dac_control_0/hold1/a_285_47# 0 0.29867f
C381 r2r_dac_control_0/hold1/a_49_47# 0 0.306903f
C382 r2r_dac_control_0/_069_ 0 0.293164f
C383 r2r_dac_control_0/_318_/a_27_47# 0 0.177187f
C384 r2r_dac_control_0/_142_ 0 0.163771f
C385 r2r_dac_control_0/_335_/a_381_47# 0 0.016397f
C386 r2r_dac_control_0/_335_/a_891_413# 0 0.160892f
C387 r2r_dac_control_0/_335_/a_1062_300# 0 0.529662f
C388 r2r_dac_control_0/_335_/a_475_413# 0 0.137184f
C389 r2r_dac_control_0/_335_/a_634_183# 0 0.150209f
C390 r2r_dac_control_0/_335_/a_193_47# 0 0.271178f
C391 r2r_dac_control_0/_335_/a_27_47# 0 0.468295f
C392 r2r_dac_control_0/_197_/a_27_47# 0 0.265166f
C393 r2r_dac_control_0/_153_ 0 0.215368f
C394 r2r_dac_control_0/_266_/a_109_93# 0 0.160708f
C395 r2r_dac_control_0/_266_/a_215_53# 0 0.142592f
C396 r2r_dac_control_0/counter\[11\] 0 0.496373f
C397 r2r_dac_control_0/_028_ 0 0.151063f
C398 r2r_dac_control_0/clknet_2_2__leaf_clk 0 1.365083f
C399 r2r_dac_control_0/_352_/a_381_47# 0 0.015369f
C400 r2r_dac_control_0/_352_/a_891_413# 0 0.161052f
C401 r2r_dac_control_0/_352_/a_1059_315# 0 0.248849f
C402 r2r_dac_control_0/_352_/a_466_413# 0 0.133203f
C403 r2r_dac_control_0/_352_/a_634_159# 0 0.142309f
C404 r2r_dac_control_0/_352_/a_193_47# 0 0.284262f
C405 r2r_dac_control_0/_352_/a_27_47# 0 0.449511f
C406 r2r_dac_control_0/_283_/a_215_47# 0 0.035725f
C407 r2r_dac_control_0/_283_/a_78_199# 0 0.15408f
C408 uio_in[0] 0 2.775601f
C409 r2r_dac_control_0/input9/a_27_47# 0 0.320141f
C410 r2r_dac_control_0/net9 0 0.897162f
C411 r2r_dac_control_0/_319_/a_29_53# 0 0.180006f
C412 rst_n 0 2.05334f
C413 r2r_dac_control_0/input11/a_75_212# 0 0.210264f
C414 r2r_dac_control_0/_102_ 0 0.109635f
C415 r2r_dac_control_0/counter\[3\] 0 0.413211f
C416 r2r_dac_control_0/_012_ 0 0.164656f
C417 r2r_dac_control_0/clknet_2_3__leaf_clk 0 1.677769f
C418 r2r_dac_control_0/_336_/a_381_47# 0 0.016397f
C419 r2r_dac_control_0/_336_/a_891_413# 0 0.160892f
C420 r2r_dac_control_0/_336_/a_1062_300# 0 0.529662f
C421 r2r_dac_control_0/_336_/a_475_413# 0 0.137184f
C422 r2r_dac_control_0/_336_/a_634_183# 0 0.150209f
C423 r2r_dac_control_0/_336_/a_193_47# 0 0.271178f
C424 r2r_dac_control_0/_336_/a_27_47# 0 0.468295f
C425 r2r_dac_control_0/_004_ 0 0.157955f
C426 r2r_dac_control_0/_148_ 0 1.037932f
C427 r2r_dac_control_0/_267_/a_215_297# 0 0.152836f
C428 r2r_dac_control_0/_267_/a_27_413# 0 0.171579f
C429 ui_in[7] 0 2.74616f
C430 r2r_dac_control_0/input8/a_27_47# 0 0.207781f
C431 r2r_dac_control_0/_353_/a_381_47# 0 0.015369f
C432 r2r_dac_control_0/_353_/a_891_413# 0 0.161052f
C433 r2r_dac_control_0/_353_/a_1059_315# 0 0.248849f
C434 r2r_dac_control_0/_353_/a_466_413# 0 0.133203f
C435 r2r_dac_control_0/_353_/a_634_159# 0 0.142309f
C436 r2r_dac_control_0/_353_/a_193_47# 0 0.284262f
C437 r2r_dac_control_0/_353_/a_27_47# 0 0.449511f
C438 r2r_dac_control_0/_037_ 0 0.154114f
C439 r2r_dac_control_0/divider\[6\] 0 0.416701f
C440 r2r_dac_control_0/_284_/a_207_413# 0 0.137402f
C441 r2r_dac_control_0/_284_/a_27_413# 0 0.196502f
C442 uio_in[1] 0 6.447606f
C443 r2r_dac_control_0/input10/a_27_47# 0 0.320141f
C444 r2r_dac_control_0/_103_ 0 0.131058f
C445 r2r_dac_control_0/net16 0 0.228252f
C446 r2r_dac_control_0/_337_/a_381_47# 0 0.016397f
C447 r2r_dac_control_0/_337_/a_891_413# 0 0.160892f
C448 r2r_dac_control_0/_337_/a_1062_300# 0 0.529662f
C449 r2r_dac_control_0/_337_/a_475_413# 0 0.137184f
C450 r2r_dac_control_0/_337_/a_634_183# 0 0.150209f
C451 r2r_dac_control_0/_337_/a_193_47# 0 0.271178f
C452 r2r_dac_control_0/_337_/a_27_47# 0 0.468295f
C453 r2r_dac_control_0/_268_/a_109_93# 0 0.160708f
C454 r2r_dac_control_0/_268_/a_215_53# 0 0.142592f
C455 ui_in[6] 0 2.802236f
C456 r2r_dac_control_0/input7/a_27_47# 0 0.207781f
C457 r2r_dac_control_0/_030_ 0 0.188667f
C458 r2r_dac_control_0/_354_/a_381_47# 0 0.015369f
C459 r2r_dac_control_0/_354_/a_891_413# 0 0.161052f
C460 r2r_dac_control_0/_354_/a_1059_315# 0 0.248849f
C461 r2r_dac_control_0/_354_/a_466_413# 0 0.133203f
C462 r2r_dac_control_0/_354_/a_634_159# 0 0.142309f
C463 r2r_dac_control_0/_354_/a_193_47# 0 0.284262f
C464 r2r_dac_control_0/_354_/a_27_47# 0 0.449511f
C465 r2r_dac_control_0/_038_ 0 0.232612f
C466 r2r_dac_control_0/counter\[15\] 0 0.659376f
C467 r2r_dac_control_0/divider\[7\] 0 0.609766f
C468 r2r_dac_control_0/_285_/a_35_297# 0 0.254573f
C469 r2r_dac_control_0/_338_/a_381_47# 0 0.016397f
C470 r2r_dac_control_0/_338_/a_891_413# 0 0.160892f
C471 r2r_dac_control_0/_338_/a_1062_300# 0 0.529662f
C472 r2r_dac_control_0/_338_/a_475_413# 0 0.137184f
C473 r2r_dac_control_0/_338_/a_634_183# 0 0.150209f
C474 r2r_dac_control_0/_338_/a_193_47# 0 0.271178f
C475 r2r_dac_control_0/_338_/a_27_47# 0 0.468295f
C476 r2r_dac_control_0/_005_ 0 0.168656f
C477 r2r_dac_control_0/_154_ 0 0.230824f
C478 r2r_dac_control_0/_269_/a_215_297# 0 0.152836f
C479 r2r_dac_control_0/_269_/a_27_413# 0 0.171579f
C480 ui_in[5] 0 2.825069f
C481 r2r_dac_control_0/input6/a_27_47# 0 0.207781f
C482 r2r_dac_control_0/_031_ 0 0.167774f
C483 r2r_dac_control_0/_355_/a_381_47# 0 0.015369f
C484 r2r_dac_control_0/_355_/a_891_413# 0 0.161052f
C485 r2r_dac_control_0/_355_/a_1059_315# 0 0.248849f
C486 r2r_dac_control_0/_355_/a_466_413# 0 0.133203f
C487 r2r_dac_control_0/_355_/a_634_159# 0 0.142309f
C488 r2r_dac_control_0/_355_/a_193_47# 0 0.284262f
C489 r2r_dac_control_0/_355_/a_27_47# 0 0.449511f
C490 r2r_dac_control_0/_039_ 0 0.259719f
C491 r2r_dac_control_0/_286_/a_27_53# 0 0.175308f
C492 r2r_dac_control_0/_286_/a_219_297# 0 0.137194f
C493 r2r_dac_control_0/_357__12/LO 0 0.165803f
C494 r2r_dac_control_0/_015_ 0 0.176197f
C495 r2r_dac_control_0/_339_/a_381_47# 0 0.016397f
C496 r2r_dac_control_0/_339_/a_891_413# 0 0.160892f
C497 r2r_dac_control_0/_339_/a_1062_300# 0 0.529662f
C498 r2r_dac_control_0/_339_/a_475_413# 0 0.137184f
C499 r2r_dac_control_0/_339_/a_634_183# 0 0.150209f
C500 r2r_dac_control_0/_339_/a_193_47# 0 0.271178f
C501 r2r_dac_control_0/_339_/a_27_47# 0 0.468295f
C502 r2r_dac_control_0/net13 0 0.11668f
C503 r2r_dac_control_0/_040_ 0 0.230406f
C504 r2r_dac_control_0/_287_/a_109_93# 0 0.160708f
C505 r2r_dac_control_0/_287_/a_215_53# 0 0.142592f
C506 r2r_dac_control_0/_356_/a_381_47# 0 0.015369f
C507 r2r_dac_control_0/_356_/a_891_413# 0 0.161052f
C508 r2r_dac_control_0/_356_/a_1059_315# 0 0.248849f
C509 r2r_dac_control_0/_356_/a_466_413# 0 0.133203f
C510 r2r_dac_control_0/_356_/a_634_159# 0 0.142309f
C511 r2r_dac_control_0/_356_/a_193_47# 0 0.284262f
C512 r2r_dac_control_0/_356_/a_27_47# 0 0.449511f
C513 ui_in[4] 0 0.711328f
C514 r2r_dac_control_0/input5/a_27_47# 0 0.207781f
C515 r2r_dac_control_0/_112_ 0 0.334037f
C516 r2r_dac_control_0/_211_/a_27_47# 0 0.174893f
C517 r2r_dac_control_0/clkbuf_2_1__f_clk/a_110_47# 0 1.73295f
C518 r2r_dac_control_0/_041_ 0 0.351716f
C519 r2r_dac_control_0/_000_ 0 0.230562f
C520 r2r_dac_control_0/net12 0 0.361147f
C521 r2r_dac_control_0/_357_/a_448_47# 0 0.013901f
C522 r2r_dac_control_0/_357_/a_1108_47# 0 0.13732f
C523 r2r_dac_control_0/_357_/a_1283_21# 0 0.389264f
C524 r2r_dac_control_0/_357_/a_543_47# 0 0.157869f
C525 r2r_dac_control_0/_357_/a_761_289# 0 0.120848f
C526 r2r_dac_control_0/_357_/a_193_47# 0 0.273213f
C527 r2r_dac_control_0/_357_/a_27_47# 0 0.495752f
C528 ui_in[3] 0 2.064625f
C529 r2r_dac_control_0/input4/a_27_47# 0 0.207781f
C530 r2r_dac_control_0/_113_ 0 0.151554f
C531 r2r_dac_control_0/_212_/a_80_21# 0 0.211154f
C532 r2r_dac_control_0/_042_ 0 0.105845f
C533 r2r_dac_control_0/_155_ 0 0.219748f
C534 r2r_dac_control_0/_289_/a_489_413# 0 0.025434f
C535 r2r_dac_control_0/_289_/a_226_47# 0 0.162324f
C536 r2r_dac_control_0/_289_/a_76_199# 0 0.140862f
C537 ui_in[2] 0 2.085923f
C538 r2r_dac_control_0/input3/a_27_47# 0 0.207781f
C539 r2r_dac_control_0/_052_ 0 0.521989f
C540 r2r_dac_control_0/_213_/a_109_93# 0 0.160708f
C541 r2r_dac_control_0/_213_/a_215_53# 0 0.142592f
C542 ui_in[1] 0 2.062965f
C543 r2r_dac_control_0/input2/a_27_47# 0 0.207781f
C544 r2r_dac_control_0/_127_ 0 0.146809f
C545 r2r_dac_control_0/_114_ 0 0.136883f
C546 r2r_dac_control_0/_111_ 0 0.159998f
C547 r2r_dac_control_0/_149_ 0 1.534441f
C548 r2r_dac_control_0/_214_/a_113_297# 0 0.034004f
C549 ui_in[0] 0 2.001586f
C550 r2r_dac_control_0/input1/a_27_47# 0 0.207781f
C551 r2r_dac_control_0/_053_ 0 1.334401f
C552 r2r_dac_control_0/_300_/a_27_47# 0 0.542977f
C553 r2r_dac_control_0/_075_ 0 0.114664f
C554 r2r_dac_control_0/net4 0 0.309257f
C555 r2r_dac_control_0/_073_ 0 0.212728f
C556 r2r_dac_control_0/_163_/a_27_47# 0 0.216317f
C557 r2r_dac_control_0/_301_/a_27_47# 0 0.28447f
C558 r2r_0/b7 0 8.831756f
C559 r2r_dac_control_0/_116_ 0 0.1519f
C560 r2r_dac_control_0/_216_/a_59_75# 0 0.177062f
C561 r2r_dac_control_0/_129_ 0 0.089789f
C562 r2r_dac_control_0/_233_/a_80_21# 0 0.209712f
C563 r2r_0/b0 0 5.49168f
C564 r2r_dac_control_0/_164_/a_215_47# 0 0.01011f
C565 r2r_dac_control_0/_164_/a_79_21# 0 0.225128f
C566 r2r_dac_control_0/_143_ 0 0.211409f
C567 r2r_dac_control_0/_250_/a_113_297# 0 0.034004f
C568 r2r_dac_control_0/_088_ 0 0.133974f
C569 r2r_dac_control_0/_181_/a_250_297# 0 0.02777f
C570 r2r_dac_control_0/_181_/a_93_21# 0 0.150721f
C571 r2r_dac_control_0/_217_/a_27_47# 0 0.174893f
C572 r2r_dac_control_0/_130_ 0 0.116032f
C573 r2r_dac_control_0/_128_ 0 0.110616f
C574 r2r_dac_control_0/_234_/a_113_297# 0 0.034004f
C575 r2r_dac_control_0/net1 0 0.368816f
C576 r2r_dac_control_0/_303_/a_113_297# 0 0.034004f
C577 r2r_dac_control_0/_071_ 0 0.159373f
C578 r2r_dac_control_0/_067_ 0 0.132817f
C579 r2r_dac_control_0/_070_ 0 0.104523f
C580 r2r_dac_control_0/_320_/a_80_21# 0 0.211154f
C581 r2r_dac_control_0/_144_ 0 0.131641f
C582 r2r_dac_control_0/_251_/a_27_47# 0 0.177187f
C583 r2r_dac_control_0/_090_ 0 0.12904f
C584 r2r_dac_control_0/_089_ 0 0.180024f
C585 r2r_dac_control_0/clknet_0_clk 0 1.846245f
C586 r2r_dac_control_0/clkbuf_2_0__f_clk/a_110_47# 0 1.73295f
C587 r2r_dac_control_0/net18 0 0.207903f
C588 r2r_dac_control_0/_131_ 0 0.112788f
C589 r2r_dac_control_0/_235_/a_113_297# 0 0.034004f
C590 r2r_dac_control_0/_011_ 0 0.175267f
C591 r2r_dac_control_0/net21 0 0.136787f
C592 r2r_dac_control_0/_321_/a_448_47# 0 0.032359f
C593 r2r_dac_control_0/_321_/a_222_93# 0 0.158855f
C594 r2r_dac_control_0/_321_/a_79_199# 0 0.148299f
C595 r2r_dac_control_0/_145_ 0 0.10199f
C596 r2r_dac_control_0/counter\[14\] 0 0.698601f
C597 r2r_dac_control_0/_252_/a_299_297# 0 0.034794f
C598 r2r_dac_control_0/_252_/a_81_21# 0 0.147141f
C599 r2r_dac_control_0/_091_ 0 0.132233f
C600 r2r_dac_control_0/_183_/a_59_75# 0 0.177062f
C601 clk 0 3.946568f
C602 r2r_dac_control_0/clkbuf_0_clk/a_110_47# 0 1.73295f
C603 r2r_dac_control_0/_119_ 0 0.14516f
C604 r2r_dac_control_0/_118_ 0 0.140742f
C605 r2r_dac_control_0/_078_ 0 1.392431f
C606 r2r_dac_control_0/_117_ 0 0.667154f
C607 r2r_dac_control_0/_115_ 0 0.186166f
C608 r2r_dac_control_0/_219_/a_227_47# 0 0.030865f
C609 r2r_dac_control_0/_219_/a_77_199# 0 0.146762f
C610 r2r_dac_control_0/_236_/a_27_47# 0 0.174893f
C611 r2r_dac_control_0/_305_/a_27_47# 0 0.031143f
C612 r2r_dac_control_0/_048_ 0 0.292809f
C613 r2r_dac_control_0/_167_/a_27_47# 0 0.542977f
C614 r2r_dac_control_0/_253_/a_215_47# 0 0.01011f
C615 r2r_dac_control_0/_253_/a_79_21# 0 0.225128f
C616 r2r_dac_control_0/_092_ 0 0.151309f
C617 r2r_dac_control_0/net22 0 0.156584f
C618 r2r_dac_control_0/_184_/a_27_47# 0 0.031143f
C619 r2r_dac_control_0/_072_ 0 0.539387f
C620 r2r_0/b3 0 4.193635f
C621 r2r_dac_control_0/_322_/a_27_47# 0 0.174893f
C622 r2r_dac_control_0/_009_ 0 0.140339f
C623 r2r_dac_control_0/_056_ 0 0.226233f
C624 r2r_dac_control_0/_058_ 0 0.158282f
C625 r2r_dac_control_0/_306_/a_113_297# 0 0.034004f
C626 r2r_dac_control_0/_133_ 0 0.537427f
C627 r2r_dac_control_0/_132_ 0 0.274153f
C628 r2r_dac_control_0/_237_/a_27_47# 0 0.177187f
C629 r2r_dac_control_0/_077_ 0 0.165882f
C630 r2r_dac_control_0/net5 0 0.418495f
C631 r2r_dac_control_0/_168_/a_505_21# 0 0.246761f
C632 r2r_dac_control_0/_168_/a_76_199# 0 0.139466f
C633 r2r_dac_control_0/net20 0 0.262933f
C634 r2r_dac_control_0/_185_/a_113_297# 0 0.034004f
C635 r2r_dac_control_0/_156_ 0 0.222705f
C636 r2r_dac_control_0/_271_/a_29_53# 0 0.180006f
C637 r2r_dac_control_0/_016_ 0 0.148404f
C638 r2r_dac_control_0/_340_/a_381_47# 0 0.016397f
C639 r2r_dac_control_0/_340_/a_891_413# 0 0.160892f
C640 r2r_dac_control_0/_340_/a_1062_300# 0 0.529662f
C641 r2r_dac_control_0/_340_/a_475_413# 0 0.137184f
C642 r2r_dac_control_0/_340_/a_634_183# 0 0.150209f
C643 r2r_dac_control_0/_340_/a_193_47# 0 0.271178f
C644 r2r_dac_control_0/_340_/a_27_47# 0 0.468295f
C645 r2r_dac_control_0/_307_/a_59_75# 0 0.177062f
C646 r2r_dac_control_0/_134_ 0 0.191206f
C647 r2r_dac_control_0/_035_ 0 0.373861f
C648 r2r_dac_control_0/_238_/a_227_47# 0 0.030865f
C649 r2r_dac_control_0/_238_/a_77_199# 0 0.146762f
C650 r2r_dac_control_0/_013_ 0 0.186012f
C651 r2r_0/b4 0 5.871322f
C652 r2r_dac_control_0/_076_ 0 0.105215f
C653 r2r_dac_control_0/_079_ 0 0.107529f
C654 r2r_dac_control_0/_169_/a_240_47# 0 0.013847f
C655 r2r_dac_control_0/_169_/a_51_297# 0 0.206675f
C656 r2r_dac_control_0/_093_ 0 0.10698f
C657 r2r_dac_control_0/_186_/a_113_297# 0 0.034004f
C658 r2r_dac_control_0/_074_ 0 0.119032f
C659 r2r_dac_control_0/_324_/a_68_297# 0 0.153866f
C660 r2r_dac_control_0/_147_ 0 0.114846f
C661 r2r_dac_control_0/_255_/a_80_21# 0 0.211154f
C662 r2r_dac_control_0/_341_/a_381_47# 0 0.015369f
C663 r2r_dac_control_0/_341_/a_891_413# 0 0.161052f
C664 r2r_dac_control_0/_341_/a_1059_315# 0 0.248849f
C665 r2r_dac_control_0/_341_/a_466_413# 0 0.133203f
C666 r2r_dac_control_0/_341_/a_634_159# 0 0.142309f
C667 r2r_dac_control_0/_341_/a_193_47# 0 0.284262f
C668 r2r_dac_control_0/_341_/a_27_47# 0 0.449511f
C669 r2r_dac_control_0/_272_/a_215_297# 0 0.152836f
C670 r2r_dac_control_0/_272_/a_27_413# 0 0.171579f
C671 r2r_dac_control_0/_308_/a_27_47# 0 0.542977f
C672 r2r_dac_control_0/_017_ 0 0.166374f
C673 r2r_dac_control_0/net19 0 0.149634f
C674 r2r_dac_control_0/_060_ 0 1.243661f
C675 r2r_dac_control_0/_187_/a_297_47# 0 0.034813f
C676 r2r_dac_control_0/_187_/a_79_21# 0 0.158207f
C677 r2r_dac_control_0/_032_ 0 0.191735f
C678 r2r_dac_control_0/_146_ 0 0.11411f
C679 r2r_dac_control_0/_256_/a_81_21# 0 0.214691f
C680 r2r_dac_control_0/_325_/a_381_47# 0 0.015369f
C681 r2r_dac_control_0/_325_/a_891_413# 0 0.161052f
C682 r2r_dac_control_0/_325_/a_1059_315# 0 0.248849f
C683 r2r_dac_control_0/_325_/a_466_413# 0 0.133203f
C684 r2r_dac_control_0/_325_/a_634_159# 0 0.142309f
C685 r2r_dac_control_0/_325_/a_193_47# 0 0.284262f
C686 r2r_dac_control_0/_325_/a_27_47# 0 0.449511f
C687 r2r_dac_control_0/counter\[1\] 0 0.691615f
C688 r2r_dac_control_0/_342_/a_381_47# 0 0.015369f
C689 r2r_dac_control_0/_342_/a_891_413# 0 0.161052f
C690 r2r_dac_control_0/_342_/a_1059_315# 0 0.248849f
C691 r2r_dac_control_0/_342_/a_466_413# 0 0.133203f
C692 r2r_dac_control_0/_342_/a_634_159# 0 0.142309f
C693 r2r_dac_control_0/_342_/a_193_47# 0 0.284262f
C694 r2r_dac_control_0/_342_/a_27_47# 0 0.449511f
C695 r2r_dac_control_0/_273_/a_109_93# 0 0.160708f
C696 r2r_dac_control_0/_273_/a_215_53# 0 0.142592f
C697 r2r_dac_control_0/_290_/a_207_413# 0 0.137402f
C698 r2r_dac_control_0/_290_/a_27_413# 0 0.196502f
C699 r2r_dac_control_0/_055_ 0 0.209131f
C700 r2r_dac_control_0/_309_/a_27_47# 0 0.031143f
C701 r2r_dac_control_0/_188_/a_27_47# 0 0.28447f
C702 r2r_dac_control_0/_326_/a_381_47# 0 0.015369f
C703 r2r_dac_control_0/_326_/a_891_413# 0 0.161052f
C704 r2r_dac_control_0/_326_/a_1059_315# 0 0.248849f
C705 r2r_dac_control_0/_326_/a_466_413# 0 0.133203f
C706 r2r_dac_control_0/_326_/a_634_159# 0 0.142309f
C707 r2r_dac_control_0/_326_/a_193_47# 0 0.284262f
C708 r2r_dac_control_0/_326_/a_27_47# 0 0.449511f
C709 r2r_dac_control_0/net11 0 0.273023f
C710 r2r_dac_control_0/_343_/a_381_47# 0 0.015369f
C711 r2r_dac_control_0/_343_/a_891_413# 0 0.161052f
C712 r2r_dac_control_0/_343_/a_1059_315# 0 0.248849f
C713 r2r_dac_control_0/_343_/a_466_413# 0 0.133203f
C714 r2r_dac_control_0/_343_/a_634_159# 0 0.142309f
C715 r2r_dac_control_0/_343_/a_193_47# 0 0.284262f
C716 r2r_dac_control_0/_343_/a_27_47# 0 0.449511f
C717 r2r_dac_control_0/_157_ 0 0.232165f
C718 r2r_dac_control_0/_274_/a_215_297# 0 0.152836f
C719 r2r_dac_control_0/_274_/a_27_413# 0 0.171579f
C720 r2r_dac_control_0/_044_ 0 0.121697f
C721 r2r_dac_control_0/divider\[3\] 0 0.358831f
C722 r2r_dac_control_0/_291_/a_27_47# 0 0.216317f
C723 r2r_dac_control_0/hold10/a_391_47# 0 0.127705f
C724 r2r_dac_control_0/hold10/a_285_47# 0 0.29867f
C725 r2r_dac_control_0/hold10/a_49_47# 0 0.306903f
C726 r2r_dac_control_0/_189_/a_285_47# 0 0.017425f
C727 r2r_dac_control_0/_189_/a_47_47# 0 0.199276f
C728 r2r_dac_control_0/_258_/a_27_47# 0 0.28447f
C729 r2r_dac_control_0/_327_/a_381_47# 0 0.015369f
C730 r2r_dac_control_0/_327_/a_891_413# 0 0.161052f
C731 r2r_dac_control_0/_327_/a_1059_315# 0 0.248849f
C732 r2r_dac_control_0/_327_/a_466_413# 0 0.133203f
C733 r2r_dac_control_0/_327_/a_634_159# 0 0.142309f
C734 r2r_dac_control_0/_327_/a_193_47# 0 0.284262f
C735 r2r_dac_control_0/_327_/a_27_47# 0 0.449511f
C736 r2r_dac_control_0/_344_/a_381_47# 0 0.015369f
C737 r2r_dac_control_0/_344_/a_891_413# 0 0.161052f
C738 r2r_dac_control_0/_344_/a_1059_315# 0 0.248849f
C739 r2r_dac_control_0/_344_/a_466_413# 0 0.133203f
C740 r2r_dac_control_0/_344_/a_634_159# 0 0.142309f
C741 r2r_dac_control_0/_344_/a_193_47# 0 0.284262f
C742 r2r_dac_control_0/_344_/a_27_47# 0 0.449511f
C743 r2r_dac_control_0/_158_ 0 0.294234f
C744 r2r_dac_control_0/net10 0 0.999061f
C745 r2r_dac_control_0/rst 0 0.938187f
C746 r2r_dac_control_0/_275_/a_109_93# 0 0.160708f
C747 r2r_dac_control_0/_275_/a_215_53# 0 0.142592f
C748 r2r_dac_control_0/_036_ 0 0.144652f
C749 r2r_dac_control_0/_292_/a_516_297# 0 0.035006f
C750 r2r_dac_control_0/_292_/a_85_193# 0 0.166604f
C751 r2r_dac_control_0/_328_/a_381_47# 0 0.015369f
C752 r2r_dac_control_0/_328_/a_891_413# 0 0.161052f
C753 r2r_dac_control_0/_328_/a_1059_315# 0 0.248849f
C754 r2r_dac_control_0/_328_/a_466_413# 0 0.133203f
C755 r2r_dac_control_0/_328_/a_634_159# 0 0.142309f
C756 r2r_dac_control_0/_328_/a_193_47# 0 0.284262f
C757 r2r_dac_control_0/_328_/a_27_47# 0 0.449511f
C758 r2r_dac_control_0/_259_/a_27_47# 0 0.542977f
C759 r2r_dac_control_0/counter\[4\] 0 0.80553f
C760 r2r_dac_control_0/_021_ 0 0.17623f
C761 r2r_dac_control_0/clknet_2_1__leaf_clk 0 1.550415f
C762 r2r_dac_control_0/_345_/a_381_47# 0 0.015369f
C763 r2r_dac_control_0/_345_/a_891_413# 0 0.161052f
C764 r2r_dac_control_0/_345_/a_1059_315# 0 0.248849f
C765 r2r_dac_control_0/_345_/a_466_413# 0 0.133203f
C766 r2r_dac_control_0/_345_/a_634_159# 0 0.142309f
C767 r2r_dac_control_0/_345_/a_193_47# 0 0.284262f
C768 r2r_dac_control_0/_345_/a_27_47# 0 0.449511f
C769 r2r_dac_control_0/net8 0 0.322867f
C770 r2r_dac_control_0/_276_/a_215_297# 0 0.152836f
C771 r2r_dac_control_0/_276_/a_27_413# 0 0.171579f
C772 r2r_dac_control_0/_329_/a_381_47# 0 0.015369f
C773 r2r_dac_control_0/_329_/a_891_413# 0 0.161052f
C774 r2r_dac_control_0/_329_/a_1059_315# 0 0.248849f
C775 r2r_dac_control_0/_329_/a_466_413# 0 0.133203f
C776 r2r_dac_control_0/_329_/a_634_159# 0 0.142309f
C777 r2r_dac_control_0/_329_/a_193_47# 0 0.284262f
C778 r2r_dac_control_0/_329_/a_27_47# 0 0.449511f
C779 r2r_dac_control_0/_200_/a_227_47# 0 0.030865f
C780 r2r_dac_control_0/_200_/a_77_199# 0 0.146762f
C781 r2r_dac_control_0/_159_ 0 0.283177f
C782 r2r_dac_control_0/counter\[5\] 0 0.645322f
C783 r2r_dac_control_0/clknet_2_0__leaf_clk 0 1.259837f
C784 r2r_dac_control_0/_346_/a_381_47# 0 0.015369f
C785 r2r_dac_control_0/_346_/a_891_413# 0 0.161052f
C786 r2r_dac_control_0/_346_/a_1059_315# 0 0.248849f
C787 r2r_dac_control_0/_346_/a_466_413# 0 0.133203f
C788 r2r_dac_control_0/_346_/a_634_159# 0 0.142309f
C789 r2r_dac_control_0/_346_/a_193_47# 0 0.284262f
C790 r2r_dac_control_0/_346_/a_27_47# 0 0.449511f
C791 r2r_dac_control_0/divider\[5\] 0 0.461407f
C792 r2r_dac_control_0/divider\[4\] 0 0.550471f
C793 r2r_dac_control_0/_294_/a_215_47# 0 0.035725f
C794 r2r_dac_control_0/_294_/a_78_199# 0 0.15408f
.ends

