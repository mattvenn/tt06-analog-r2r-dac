magic
tech sky130A
magscale 1 2
timestamp 1709130371
<< metal1 >>
rect 26234 29400 26240 29521
rect 26361 29400 26367 29521
rect 21740 29166 21860 29172
rect 21860 29046 22160 29166
rect 22634 29160 22640 29280
rect 22760 29160 22766 29280
rect 23274 29180 23280 29300
rect 23400 29180 23406 29300
rect 23854 29200 23860 29320
rect 23980 29200 23986 29320
rect 21740 29040 21860 29046
rect 22040 28840 22160 29046
rect 22640 28840 22760 29160
rect 23280 28840 23400 29180
rect 23860 28840 23980 29200
rect 24454 29180 24460 29300
rect 24580 29180 24586 29300
rect 25054 29180 25060 29300
rect 25180 29180 25186 29300
rect 25654 29180 25660 29300
rect 25780 29180 25786 29300
rect 24460 28820 24580 29180
rect 25060 28840 25180 29180
rect 25660 28840 25780 29180
rect 26240 28840 26361 29400
rect 27260 19440 27700 19560
rect 20594 15540 20600 15740
rect 20800 15540 20806 15740
rect 20600 13980 20800 15540
rect 27580 7260 27700 19440
rect 27580 7134 27700 7140
<< via1 >>
rect 26240 29400 26361 29521
rect 21740 29046 21860 29166
rect 22640 29160 22760 29280
rect 23280 29180 23400 29300
rect 23860 29200 23980 29320
rect 24460 29180 24580 29300
rect 25060 29180 25180 29300
rect 25660 29180 25780 29300
rect 20600 15540 20800 15740
rect 27580 7140 27700 7260
<< metal2 >>
rect 3948 44538 4008 44547
rect 3948 44469 4008 44478
rect 3950 41864 4006 44469
rect 5250 44339 5310 44341
rect 5243 44283 5252 44339
rect 5308 44283 5317 44339
rect 5250 41703 5310 44283
rect 6515 44089 6524 44149
rect 6584 44089 6593 44149
rect 6526 41737 6582 44089
rect 7809 43931 7869 43933
rect 7802 43875 7811 43931
rect 7867 43875 7876 43931
rect 7809 41727 7869 43875
rect 9096 43700 9152 43707
rect 9094 43698 9154 43700
rect 9094 43642 9096 43698
rect 9152 43642 9154 43698
rect 9094 41815 9154 43642
rect 10388 43452 10448 43461
rect 10388 43383 10448 43392
rect 10390 41801 10446 43383
rect 11680 43202 11740 43204
rect 11673 43146 11682 43202
rect 11738 43146 11747 43202
rect 11680 41767 11740 43146
rect 12964 43012 13024 43021
rect 12964 42943 13024 42952
rect 12966 41857 13022 42943
rect 14242 42786 14302 42788
rect 14235 42730 14244 42786
rect 14300 42730 14309 42786
rect 14242 41759 14302 42730
rect 15540 42594 15600 42603
rect 15540 42525 15600 42534
rect 15542 41897 15598 42525
rect 16826 42397 16886 42399
rect 16819 42341 16828 42397
rect 16884 42341 16893 42397
rect 16826 41835 16886 42341
rect 18107 42144 18116 42204
rect 18176 42144 18185 42204
rect 18118 41872 18174 42144
rect 26240 29756 26361 29761
rect 26236 29645 26245 29756
rect 26356 29645 26365 29756
rect 26240 29521 26361 29645
rect 22640 29495 22760 29500
rect 23280 29495 23400 29500
rect 23860 29495 23980 29500
rect 24460 29495 24580 29500
rect 25060 29495 25180 29500
rect 25660 29495 25780 29500
rect 22636 29385 22645 29495
rect 22755 29385 22764 29495
rect 23276 29385 23285 29495
rect 23395 29385 23404 29495
rect 23856 29385 23865 29495
rect 23975 29385 23984 29495
rect 24456 29385 24465 29495
rect 24575 29385 24584 29495
rect 25056 29385 25065 29495
rect 25175 29385 25184 29495
rect 25656 29385 25665 29495
rect 25775 29385 25784 29495
rect 26240 29394 26361 29400
rect 22640 29280 22760 29385
rect 21465 29166 21575 29170
rect 21460 29161 21740 29166
rect 21460 29051 21465 29161
rect 21575 29051 21740 29161
rect 21460 29046 21740 29051
rect 21860 29046 21866 29166
rect 23280 29300 23400 29385
rect 23860 29320 23980 29385
rect 23860 29194 23980 29200
rect 24460 29300 24580 29385
rect 23280 29174 23400 29180
rect 24460 29174 24580 29180
rect 25060 29300 25180 29385
rect 25060 29174 25180 29180
rect 25660 29300 25780 29385
rect 25660 29174 25780 29180
rect 22640 29154 22760 29160
rect 21465 29042 21575 29046
rect 20600 16395 20800 16400
rect 20596 16205 20605 16395
rect 20795 16205 20804 16395
rect 20600 15740 20800 16205
rect 20600 15534 20800 15540
rect 27574 7140 27580 7260
rect 27700 7140 27706 7260
rect 27580 5280 27700 7140
rect 29465 5280 29575 5284
rect 27580 5275 29580 5280
rect 27580 5165 29465 5275
rect 29575 5165 29580 5275
rect 27580 5160 29580 5165
rect 29465 5156 29575 5160
<< via2 >>
rect 3948 44478 4008 44538
rect 5252 44283 5308 44339
rect 6524 44089 6584 44149
rect 7811 43875 7867 43931
rect 9096 43642 9152 43698
rect 10388 43392 10448 43452
rect 11682 43146 11738 43202
rect 12964 42952 13024 43012
rect 14244 42730 14300 42786
rect 15540 42534 15600 42594
rect 16828 42341 16884 42397
rect 18116 42144 18176 42204
rect 26245 29645 26356 29756
rect 22645 29385 22755 29495
rect 23285 29385 23395 29495
rect 23865 29385 23975 29495
rect 24465 29385 24575 29495
rect 25065 29385 25175 29495
rect 25665 29385 25775 29495
rect 21465 29051 21575 29161
rect 20605 16205 20795 16395
rect 29465 5165 29575 5275
<< metal3 >>
rect 3943 44538 4013 44543
rect 22870 44538 22876 44540
rect 3943 44478 3948 44538
rect 4008 44478 22876 44538
rect 3943 44473 4013 44478
rect 22870 44476 22876 44478
rect 22940 44476 22946 44540
rect 5247 44341 5313 44344
rect 23612 44343 23676 44349
rect 5247 44339 23612 44341
rect 5247 44283 5252 44339
rect 5308 44283 23612 44339
rect 5247 44281 23612 44283
rect 5247 44278 5313 44281
rect 23612 44273 23676 44279
rect 6519 44149 6589 44154
rect 24345 44151 24409 44157
rect 6519 44089 6524 44149
rect 6584 44089 24345 44149
rect 6519 44084 6589 44089
rect 24345 44081 24409 44087
rect 7806 43933 7872 43936
rect 25084 43935 25148 43941
rect 7806 43931 25084 43933
rect 7806 43875 7811 43931
rect 7867 43875 25084 43931
rect 7806 43873 25084 43875
rect 7806 43870 7872 43873
rect 25084 43865 25148 43871
rect 9091 43700 9157 43703
rect 25814 43700 25820 43702
rect 9091 43698 25820 43700
rect 9091 43642 9096 43698
rect 9152 43642 25820 43698
rect 9091 43640 25820 43642
rect 9091 43637 9157 43640
rect 25814 43638 25820 43640
rect 25884 43638 25890 43702
rect 10383 43452 10453 43457
rect 26552 43454 26616 43460
rect 10383 43392 10388 43452
rect 10448 43392 26552 43452
rect 10383 43387 10453 43392
rect 26552 43384 26616 43390
rect 11677 43204 11743 43207
rect 27292 43206 27356 43212
rect 11677 43202 27292 43204
rect 11677 43146 11682 43202
rect 11738 43146 27292 43202
rect 11677 43144 27292 43146
rect 11677 43141 11743 43144
rect 27292 43136 27356 43142
rect 12959 43012 13029 43017
rect 28018 43012 28024 43014
rect 12959 42952 12964 43012
rect 13024 42952 28024 43012
rect 12959 42947 13029 42952
rect 28018 42950 28024 42952
rect 28088 42950 28094 43014
rect 14239 42788 14305 42791
rect 28764 42790 28828 42796
rect 14239 42786 28764 42788
rect 14239 42730 14244 42786
rect 14300 42730 28764 42786
rect 14239 42728 28764 42730
rect 14239 42725 14305 42728
rect 28764 42720 28828 42726
rect 15535 42594 15605 42599
rect 29486 42594 29492 42596
rect 15535 42534 15540 42594
rect 15600 42534 29492 42594
rect 15535 42529 15605 42534
rect 29486 42532 29492 42534
rect 29556 42532 29562 42596
rect 16823 42399 16889 42402
rect 30236 42401 30300 42407
rect 16823 42397 30236 42399
rect 16823 42341 16828 42397
rect 16884 42341 30236 42397
rect 16823 42339 30236 42341
rect 16823 42336 16889 42339
rect 30236 42331 30300 42337
rect 18111 42204 18181 42209
rect 30973 42206 31037 42212
rect 18111 42144 18116 42204
rect 18176 42144 30973 42204
rect 18111 42139 18181 42144
rect 30973 42136 31037 42142
rect 18840 40460 26360 40580
rect 18880 38556 25780 38676
rect 18840 36652 25180 36772
rect 18840 34748 24580 34868
rect 18860 32844 23980 32964
rect 18960 30940 23400 31060
rect 19820 29680 22760 29800
rect 19820 29156 19940 29680
rect 22640 29495 22760 29680
rect 22640 29385 22645 29495
rect 22755 29385 22760 29495
rect 22640 29380 22760 29385
rect 23280 29495 23400 30940
rect 23280 29385 23285 29495
rect 23395 29385 23400 29495
rect 23280 29380 23400 29385
rect 23860 29495 23980 32844
rect 23860 29385 23865 29495
rect 23975 29385 23980 29495
rect 23860 29380 23980 29385
rect 24460 29495 24580 34748
rect 24460 29385 24465 29495
rect 24575 29385 24580 29495
rect 24460 29380 24580 29385
rect 25060 29495 25180 36652
rect 25060 29385 25065 29495
rect 25175 29385 25180 29495
rect 25060 29380 25180 29385
rect 25660 29495 25780 38556
rect 26240 29761 26360 40460
rect 26240 29756 26361 29761
rect 26240 29645 26245 29756
rect 26356 29645 26361 29756
rect 26240 29640 26361 29645
rect 25660 29385 25665 29495
rect 25775 29385 25780 29495
rect 25660 29380 25780 29385
rect 18920 29036 19940 29156
rect 20940 29161 21580 29166
rect 20940 29051 21465 29161
rect 21575 29051 21580 29161
rect 20940 29046 21580 29051
rect 20940 27252 21060 29046
rect 18940 27132 21060 27252
rect 5310 25300 5630 25306
rect 12760 25300 13080 25306
rect 182 24980 188 25300
rect 508 24980 5310 25300
rect 5630 24980 9056 25300
rect 9376 24980 12760 25300
rect 13080 24980 16450 25300
rect 16770 24980 16780 25300
rect 5310 24974 5630 24980
rect 12760 24974 13080 24980
rect 20600 24231 20800 24232
rect 20595 24033 20601 24231
rect 20799 24033 20805 24231
rect 20600 16395 20800 24033
rect 20600 16205 20605 16395
rect 20795 16205 20800 16395
rect 20600 16200 20800 16205
rect 31313 5280 31431 5285
rect 29460 5279 31432 5280
rect 29460 5275 31313 5279
rect 29460 5165 29465 5275
rect 29575 5165 31313 5275
rect 29460 5161 31313 5165
rect 31431 5161 31432 5279
rect 29460 5160 31432 5161
rect 31313 5155 31431 5160
<< via3 >>
rect 22876 44476 22940 44540
rect 23612 44279 23676 44343
rect 24345 44087 24409 44151
rect 25084 43871 25148 43935
rect 25820 43638 25884 43702
rect 26552 43390 26616 43454
rect 27292 43142 27356 43206
rect 28024 42950 28088 43014
rect 28764 42726 28828 42790
rect 29492 42532 29556 42596
rect 30236 42337 30300 42401
rect 30973 42142 31037 42206
rect 188 24980 508 25300
rect 5310 24980 5630 25300
rect 9056 24980 9376 25300
rect 12760 24980 13080 25300
rect 16450 24980 16770 25300
rect 20601 24033 20799 24231
rect 31313 5161 31431 5279
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44723 5274 45152
rect 5950 44723 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 3547 44663 6010 44723
rect 200 25301 500 44152
rect 1688 43545 1988 44256
rect 3547 43545 3607 44663
rect 22878 44541 22938 45152
rect 22875 44540 22941 44541
rect 22875 44476 22876 44540
rect 22940 44476 22941 44540
rect 22875 44475 22941 44476
rect 23614 44344 23674 45152
rect 24350 45117 24410 45152
rect 24347 44952 24410 45117
rect 23611 44343 23677 44344
rect 23611 44279 23612 44343
rect 23676 44279 23677 44343
rect 23611 44278 23677 44279
rect 24347 44152 24407 44952
rect 24344 44151 24410 44152
rect 24344 44087 24345 44151
rect 24409 44087 24410 44151
rect 24344 44086 24410 44087
rect 25086 43936 25146 45152
rect 25083 43935 25149 43936
rect 25083 43871 25084 43935
rect 25148 43871 25149 43935
rect 25083 43870 25149 43871
rect 25822 43703 25882 45152
rect 26558 45117 26618 45152
rect 26554 44952 26618 45117
rect 25819 43702 25885 43703
rect 25819 43638 25820 43702
rect 25884 43638 25885 43702
rect 25819 43637 25885 43638
rect 1668 43485 3607 43545
rect 187 25300 509 25301
rect 187 24980 188 25300
rect 508 24980 510 25300
rect 187 24979 509 24980
rect 200 1000 500 24979
rect 1688 24290 1988 43485
rect 26554 43455 26614 44952
rect 26551 43454 26617 43455
rect 26551 43390 26552 43454
rect 26616 43390 26617 43454
rect 26551 43389 26617 43390
rect 27294 43207 27354 45152
rect 28030 45117 28090 45152
rect 28026 44952 28090 45117
rect 27291 43206 27357 43207
rect 27291 43142 27292 43206
rect 27356 43142 27357 43206
rect 27291 43141 27357 43142
rect 28026 43015 28086 44952
rect 28023 43014 28089 43015
rect 28023 42950 28024 43014
rect 28088 42950 28089 43014
rect 28023 42949 28089 42950
rect 28766 42791 28826 45152
rect 29502 45125 29562 45152
rect 29494 44952 29562 45125
rect 28763 42790 28829 42791
rect 28763 42726 28764 42790
rect 28828 42726 28829 42790
rect 28763 42725 28829 42726
rect 29494 42597 29554 44952
rect 29491 42596 29557 42597
rect 29491 42532 29492 42596
rect 29556 42532 29557 42596
rect 29491 42531 29557 42532
rect 30238 42402 30298 45152
rect 30974 45074 31034 45152
rect 30974 44952 31035 45074
rect 31710 44952 31770 45152
rect 30235 42401 30301 42402
rect 30235 42337 30236 42401
rect 30300 42337 30301 42401
rect 30235 42336 30301 42337
rect 30975 42207 31035 44952
rect 30972 42206 31038 42207
rect 30972 42142 30973 42206
rect 31037 42142 31038 42206
rect 30972 42141 31038 42142
rect 5310 25301 5630 27340
rect 5309 25300 5631 25301
rect 5309 24980 5310 25300
rect 5630 24980 5631 25300
rect 5309 24979 5631 24980
rect 7190 24290 7490 27070
rect 9056 25301 9376 27418
rect 9055 25300 9377 25301
rect 9055 24980 9056 25300
rect 9376 24980 9377 25300
rect 9055 24979 9377 24980
rect 10930 24290 11230 27110
rect 12760 25301 13080 27494
rect 12759 25300 13081 25301
rect 12759 24980 12760 25300
rect 13080 24980 13081 25300
rect 12759 24979 13081 24980
rect 14590 24290 14890 27170
rect 16450 25301 16770 27550
rect 16449 25300 16771 25301
rect 16449 24980 16450 25300
rect 16770 24980 16771 25300
rect 16449 24979 16771 24980
rect 1688 24232 18790 24290
rect 1688 24231 20800 24232
rect 1688 24033 20601 24231
rect 20799 24033 20800 24231
rect 1688 24032 20800 24033
rect 1688 23990 18790 24032
rect 1688 1104 1988 23990
rect 31312 5279 31432 5280
rect 31312 5161 31313 5279
rect 31431 5161 31432 5279
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31312 0 31432 5161
use r2r  r2r_0
timestamp 1709129632
transform 1 0 23200 0 1 11400
box -2600 2400 4200 17600
use r2r_dac_control  r2r_dac_control_0
timestamp 1708507682
transform 1 0 3104 0 1 26036
box 514 496 16000 16000
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 1688 1104 1988 44256 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
