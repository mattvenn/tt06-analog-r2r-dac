magic
tech sky130A
timestamp 1708444847
<< xpolycontact >>
rect -17 50 17 266
rect -17 -266 17 -50
<< ppolyres >>
rect -17 -50 17 50
<< viali >>
rect -9 58 9 257
rect -9 -257 9 -58
<< metal1 >>
rect -12 257 12 263
rect -12 58 -9 257
rect 9 58 12 257
rect -12 52 12 58
rect -12 -58 12 -52
rect -12 -257 -9 -58
rect 9 -257 12 -58
rect -12 -263 12 -257
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 1.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 2.026k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
