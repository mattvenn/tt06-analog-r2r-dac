magic
tech sky130A
magscale 1 2
timestamp 1708461890
<< metal1 >>
rect 22480 31060 22600 31066
rect 23474 31060 23480 31180
rect 23600 31060 23606 31180
rect 22600 30940 22920 31060
rect 22480 30934 22600 30940
rect 21400 29800 21520 29806
rect 21520 29680 22640 29800
rect 21400 29674 21520 29680
rect 21340 29340 21460 29346
rect 21460 29220 22320 29340
rect 21340 29214 21460 29220
rect 22520 29200 22640 29680
rect 22800 29220 22920 30940
rect 23174 30500 23180 30620
rect 23300 30500 23306 30620
rect 23180 29220 23300 30500
rect 23480 29200 23600 31060
rect 23774 31040 23780 31160
rect 23900 31040 23906 31160
rect 23780 29200 23900 31040
rect 24074 31020 24080 31140
rect 24200 31020 24206 31140
rect 24080 29240 24200 31020
rect 24354 30820 24360 30940
rect 24480 30820 24486 30940
rect 24360 29800 24480 30820
rect 24360 29680 24580 29800
rect 24460 29240 24580 29680
rect 24296 27666 25140 27866
rect 24943 6080 25138 27666
rect 24943 5583 25140 6080
rect 25020 5280 25140 5583
rect 26060 5280 26180 5286
rect 25020 5160 26060 5280
rect 26060 5154 26180 5160
<< via1 >>
rect 23480 31060 23600 31180
rect 22480 30940 22600 31060
rect 21400 29680 21520 29800
rect 21340 29220 21460 29340
rect 23180 30500 23300 30620
rect 23780 31040 23900 31160
rect 24080 31020 24200 31140
rect 24360 30820 24480 30940
rect 26060 5160 26180 5280
<< metal2 >>
rect 23480 32335 23600 32340
rect 23476 32225 23485 32335
rect 23595 32225 23604 32335
rect 23180 31475 23300 31480
rect 23176 31365 23185 31475
rect 23295 31365 23304 31475
rect 21285 31060 21395 31064
rect 21280 31055 22480 31060
rect 21280 30945 21285 31055
rect 21395 30945 22480 31055
rect 21280 30940 22480 30945
rect 22600 30940 22606 31060
rect 21285 30936 21395 30940
rect 23180 30620 23300 31365
rect 23480 31180 23600 32225
rect 23780 32035 23900 32040
rect 23776 31925 23785 32035
rect 23895 31925 23904 32035
rect 23480 31054 23600 31060
rect 23780 31160 23900 31925
rect 24080 31815 24200 31820
rect 24076 31705 24085 31815
rect 24195 31705 24204 31815
rect 24360 31795 24480 31800
rect 23780 31034 23900 31040
rect 24080 31140 24200 31705
rect 24356 31685 24365 31795
rect 24475 31685 24484 31795
rect 24080 31014 24200 31020
rect 24360 30940 24480 31685
rect 24360 30814 24480 30820
rect 23180 30494 23300 30500
rect 20945 29800 21055 29804
rect 20940 29795 21400 29800
rect 20940 29685 20945 29795
rect 21055 29685 21400 29795
rect 20940 29680 21400 29685
rect 21520 29680 21526 29800
rect 20945 29676 21055 29680
rect 20945 29340 21055 29344
rect 20940 29335 21340 29340
rect 20940 29225 20945 29335
rect 21055 29225 21340 29335
rect 20940 29220 21340 29225
rect 21460 29220 21466 29340
rect 20945 29216 21055 29220
rect 29465 5280 29575 5284
rect 26054 5160 26060 5280
rect 26180 5275 29580 5280
rect 26180 5165 29465 5275
rect 29575 5165 29580 5275
rect 26180 5160 29580 5165
rect 29465 5156 29575 5160
<< via2 >>
rect 23485 32225 23595 32335
rect 23185 31365 23295 31475
rect 21285 30945 21395 31055
rect 23785 31925 23895 32035
rect 24085 31705 24195 31815
rect 24365 31685 24475 31795
rect 20945 29685 21055 29795
rect 20945 29225 21055 29335
rect 29465 5165 29575 5275
<< metal3 >>
rect 18840 40460 24480 40580
rect 18880 38556 24200 38676
rect 18840 36652 23900 36772
rect 18840 34748 23600 34868
rect 18860 32844 23300 32964
rect 23180 31475 23300 32844
rect 23480 32335 23600 34748
rect 23480 32225 23485 32335
rect 23595 32225 23600 32335
rect 23480 32220 23600 32225
rect 23780 32035 23900 36652
rect 23780 31925 23785 32035
rect 23895 31925 23900 32035
rect 23780 31920 23900 31925
rect 24080 31815 24200 38556
rect 24080 31705 24085 31815
rect 24195 31705 24200 31815
rect 24080 31700 24200 31705
rect 24360 31795 24480 40460
rect 24360 31685 24365 31795
rect 24475 31685 24480 31795
rect 24360 31680 24480 31685
rect 23180 31365 23185 31475
rect 23295 31365 23300 31475
rect 23180 31360 23300 31365
rect 18960 31055 21400 31060
rect 18960 30945 21285 31055
rect 21395 30945 21400 31055
rect 18960 30940 21400 30945
rect 19820 29795 21060 29800
rect 19820 29685 20945 29795
rect 21055 29685 21060 29795
rect 19820 29680 21060 29685
rect 19820 29156 19940 29680
rect 18920 29036 19940 29156
rect 20940 29335 21060 29340
rect 20940 29225 20945 29335
rect 21055 29225 21060 29335
rect 20940 27252 21060 29225
rect 18940 27132 21060 27252
rect 31313 5280 31431 5285
rect 29460 5279 31432 5280
rect 29460 5275 31313 5279
rect 29460 5165 29465 5275
rect 29575 5165 31313 5275
rect 29460 5161 31313 5165
rect 31431 5161 31432 5279
rect 29460 5160 31432 5161
rect 31313 5155 31431 5160
<< via3 >>
rect 31313 5161 31431 5279
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 25300 500 44152
rect 200 1000 500 24980
rect 1688 24290 1988 44256
rect 5340 25276 5660 27260
rect 5340 25004 5364 25276
rect 5636 25004 5660 25276
rect 5340 24980 5660 25004
rect 7190 24290 7490 27070
rect 9040 25276 9360 27260
rect 9040 25004 9064 25276
rect 9336 25004 9360 25276
rect 9040 24980 9360 25004
rect 10930 24290 11230 27110
rect 12760 25276 13080 27560
rect 12760 25004 12784 25276
rect 13056 25004 13080 25276
rect 12760 24980 13080 25004
rect 14590 24290 14890 27170
rect 16460 25276 16780 27700
rect 16460 25004 16484 25276
rect 16756 25004 16780 25276
rect 16460 24980 16780 25004
rect 1688 23990 18790 24290
rect 1688 1104 1988 23990
rect 31312 5279 31432 5280
rect 31312 5161 31313 5279
rect 31431 5161 31432 5279
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31312 0 31432 5161
<< via4 >>
rect 190 24980 510 25300
rect 5364 25004 5636 25276
rect 9064 25004 9336 25276
rect 12784 25004 13056 25276
rect 16484 25004 16756 25276
<< metal5 >>
rect 166 25300 534 25324
rect 166 24980 190 25300
rect 510 25276 18540 25300
rect 510 25004 5364 25276
rect 5636 25004 9064 25276
rect 9336 25004 12784 25276
rect 13056 25004 16484 25276
rect 16756 25004 18540 25276
rect 510 24980 18540 25004
rect 166 24956 534 24980
use r2r  r2r_0
timestamp 1708461036
transform 1 0 21996 0 1 27306
box 160 -600 2600 2080
use r2r_dac_control  r2r_dac_control_0
timestamp 1708461890
transform 1 0 3104 0 1 26036
box 514 496 16000 16000
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 1688 1104 1988 44256 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
