* NGSPICE file created from r2r_parax.ext - technology: sky130A

.subckt r2r_parax b0 b1 b2 b3 b4 b5 b6 b7 out VSUBS GND
X0 b7 out VSUBS.t2 sky130_fd_pr__res_high_po_0p35 l=40.16
X1 a_n434_6998# a_166_2566# VSUBS.t3 sky130_fd_pr__res_high_po_0p35 l=20.16
X2 a_766_6998# a_1366_2566# VSUBS.t6 sky130_fd_pr__res_high_po_0p35 l=20.16
X3 b0 a_n1834_10998# VSUBS.t5 sky130_fd_pr__res_high_po_0p35 l=40.16
X4 b6 a_1966_6998# VSUBS.t0 sky130_fd_pr__res_high_po_0p35 l=40.16
X5 b3 a_166_2566# VSUBS.t1 sky130_fd_pr__res_high_po_0p35 l=40.16
X6 b5 a_1366_2566# VSUBS.t4 sky130_fd_pr__res_high_po_0p35 l=40.16
X7 a_n1834_10998# a_n1034_2566# VSUBS.t5 sky130_fd_pr__res_high_po_0p35 l=20.16
X8 b1 a_n1034_2566# VSUBS.t7 sky130_fd_pr__res_high_po_0p35 l=40.16
X9 a_1966_6998# out VSUBS.t0 sky130_fd_pr__res_high_po_0p35 l=20.16
X10 a_n1834_10998# GND VSUBS.t8 sky130_fd_pr__res_high_po_0p35 l=40.16
X11 a_766_6998# a_166_2566# VSUBS.t1 sky130_fd_pr__res_high_po_0p35 l=20.16
X12 a_1966_6998# a_1366_2566# VSUBS.t4 sky130_fd_pr__res_high_po_0p35 l=20.16
X13 b2 a_n434_6998# VSUBS.t3 sky130_fd_pr__res_high_po_0p35 l=40.16
X14 b4 a_766_6998# VSUBS.t6 sky130_fd_pr__res_high_po_0p35 l=40.16
X15 a_n434_6998# a_n1034_2566# VSUBS.t7 sky130_fd_pr__res_high_po_0p35 l=20.16
R0 VSUBS.n134 VSUBS.n5 27093.3
R1 VSUBS.n138 VSUBS.n5 27093.3
R2 VSUBS.n134 VSUBS.n6 27093.3
R3 VSUBS.n138 VSUBS.n6 27093.3
R4 VSUBS.n120 VSUBS.n9 27093.3
R5 VSUBS.n124 VSUBS.n9 27093.3
R6 VSUBS.n120 VSUBS.n10 27093.3
R7 VSUBS.n124 VSUBS.n10 27093.3
R8 VSUBS.n106 VSUBS.n13 27093.3
R9 VSUBS.n110 VSUBS.n13 27093.3
R10 VSUBS.n106 VSUBS.n14 27093.3
R11 VSUBS.n110 VSUBS.n14 27093.3
R12 VSUBS.n92 VSUBS.n17 27093.3
R13 VSUBS.n96 VSUBS.n17 27093.3
R14 VSUBS.n92 VSUBS.n18 27093.3
R15 VSUBS.n96 VSUBS.n18 27093.3
R16 VSUBS.n78 VSUBS.n21 27093.3
R17 VSUBS.n82 VSUBS.n21 27093.3
R18 VSUBS.n78 VSUBS.n22 27093.3
R19 VSUBS.n82 VSUBS.n22 27093.3
R20 VSUBS.n64 VSUBS.n25 27093.3
R21 VSUBS.n68 VSUBS.n25 27093.3
R22 VSUBS.n64 VSUBS.n26 27093.3
R23 VSUBS.n68 VSUBS.n26 27093.3
R24 VSUBS.n50 VSUBS.n29 27093.3
R25 VSUBS.n54 VSUBS.n29 27093.3
R26 VSUBS.n50 VSUBS.n30 27093.3
R27 VSUBS.n54 VSUBS.n30 27093.3
R28 VSUBS.n40 VSUBS.n32 27093.3
R29 VSUBS.n36 VSUBS.n33 27093.3
R30 VSUBS.n40 VSUBS.n33 27093.3
R31 VSUBS.n142 VSUBS.n2 27093.3
R32 VSUBS.n144 VSUBS.n2 27093.3
R33 VSUBS.n144 VSUBS.n3 27093.3
R34 VSUBS.n132 VSUBS.n126 15505.1
R35 VSUBS.n126 VSUBS.n4 15505.1
R36 VSUBS.n132 VSUBS.n127 15505.1
R37 VSUBS.n127 VSUBS.n4 15505.1
R38 VSUBS.n118 VSUBS.n112 15505.1
R39 VSUBS.n112 VSUBS.n8 15505.1
R40 VSUBS.n118 VSUBS.n113 15505.1
R41 VSUBS.n113 VSUBS.n8 15505.1
R42 VSUBS.n104 VSUBS.n98 15505.1
R43 VSUBS.n98 VSUBS.n12 15505.1
R44 VSUBS.n104 VSUBS.n99 15505.1
R45 VSUBS.n99 VSUBS.n12 15505.1
R46 VSUBS.n90 VSUBS.n84 15505.1
R47 VSUBS.n84 VSUBS.n16 15505.1
R48 VSUBS.n90 VSUBS.n85 15505.1
R49 VSUBS.n85 VSUBS.n16 15505.1
R50 VSUBS.n76 VSUBS.n70 15505.1
R51 VSUBS.n70 VSUBS.n20 15505.1
R52 VSUBS.n76 VSUBS.n71 15505.1
R53 VSUBS.n71 VSUBS.n20 15505.1
R54 VSUBS.n62 VSUBS.n56 15505.1
R55 VSUBS.n56 VSUBS.n24 15505.1
R56 VSUBS.n62 VSUBS.n57 15505.1
R57 VSUBS.n57 VSUBS.n24 15505.1
R58 VSUBS.n48 VSUBS.n42 15505.1
R59 VSUBS.n42 VSUBS.n28 15505.1
R60 VSUBS.n48 VSUBS.n43 15505.1
R61 VSUBS.n43 VSUBS.n28 15505.1
R62 VSUBS.n135 VSUBS.n7 1760.38
R63 VSUBS.n137 VSUBS.n7 1760.38
R64 VSUBS.n136 VSUBS.n135 1760.38
R65 VSUBS.n137 VSUBS.n136 1760.38
R66 VSUBS.n121 VSUBS.n11 1760.38
R67 VSUBS.n123 VSUBS.n11 1760.38
R68 VSUBS.n122 VSUBS.n121 1760.38
R69 VSUBS.n123 VSUBS.n122 1760.38
R70 VSUBS.n107 VSUBS.n15 1760.38
R71 VSUBS.n109 VSUBS.n15 1760.38
R72 VSUBS.n108 VSUBS.n107 1760.38
R73 VSUBS.n109 VSUBS.n108 1760.38
R74 VSUBS.n93 VSUBS.n19 1760.38
R75 VSUBS.n95 VSUBS.n19 1760.38
R76 VSUBS.n94 VSUBS.n93 1760.38
R77 VSUBS.n95 VSUBS.n94 1760.38
R78 VSUBS.n79 VSUBS.n23 1760.38
R79 VSUBS.n81 VSUBS.n23 1760.38
R80 VSUBS.n80 VSUBS.n79 1760.38
R81 VSUBS.n81 VSUBS.n80 1760.38
R82 VSUBS.n65 VSUBS.n27 1760.38
R83 VSUBS.n67 VSUBS.n27 1760.38
R84 VSUBS.n66 VSUBS.n65 1760.38
R85 VSUBS.n67 VSUBS.n66 1760.38
R86 VSUBS.n51 VSUBS.n31 1760.38
R87 VSUBS.n53 VSUBS.n31 1760.38
R88 VSUBS.n52 VSUBS.n51 1760.38
R89 VSUBS.n53 VSUBS.n52 1760.38
R90 VSUBS.n37 VSUBS.n34 1760.38
R91 VSUBS.n39 VSUBS.n34 1760.38
R92 VSUBS.n38 VSUBS.n37 1760.38
R93 VSUBS.n39 VSUBS.n38 1760.38
R94 VSUBS.n141 VSUBS.n0 1760.38
R95 VSUBS.n141 VSUBS.n1 1760.38
R96 VSUBS.n145 VSUBS.n1 1760.38
R97 VSUBS.n146 VSUBS.n0 1432.47
R98 VSUBS.n131 VSUBS.n128 1007.44
R99 VSUBS.n129 VSUBS.n128 1007.44
R100 VSUBS.n131 VSUBS.n130 1007.44
R101 VSUBS.n130 VSUBS.n129 1007.44
R102 VSUBS.n117 VSUBS.n114 1007.44
R103 VSUBS.n115 VSUBS.n114 1007.44
R104 VSUBS.n117 VSUBS.n116 1007.44
R105 VSUBS.n116 VSUBS.n115 1007.44
R106 VSUBS.n103 VSUBS.n100 1007.44
R107 VSUBS.n101 VSUBS.n100 1007.44
R108 VSUBS.n103 VSUBS.n102 1007.44
R109 VSUBS.n102 VSUBS.n101 1007.44
R110 VSUBS.n89 VSUBS.n86 1007.44
R111 VSUBS.n87 VSUBS.n86 1007.44
R112 VSUBS.n89 VSUBS.n88 1007.44
R113 VSUBS.n88 VSUBS.n87 1007.44
R114 VSUBS.n75 VSUBS.n72 1007.44
R115 VSUBS.n73 VSUBS.n72 1007.44
R116 VSUBS.n75 VSUBS.n74 1007.44
R117 VSUBS.n74 VSUBS.n73 1007.44
R118 VSUBS.n61 VSUBS.n58 1007.44
R119 VSUBS.n59 VSUBS.n58 1007.44
R120 VSUBS.n61 VSUBS.n60 1007.44
R121 VSUBS.n60 VSUBS.n59 1007.44
R122 VSUBS.n47 VSUBS.n44 1007.44
R123 VSUBS.n45 VSUBS.n44 1007.44
R124 VSUBS.n47 VSUBS.n46 1007.44
R125 VSUBS.n46 VSUBS.n45 1007.44
R126 VSUBS.n46 VSUBS.n43 292.5
R127 VSUBS.n43 VSUBS.t0 292.5
R128 VSUBS.n44 VSUBS.n42 292.5
R129 VSUBS.n42 VSUBS.t0 292.5
R130 VSUBS.n60 VSUBS.n57 292.5
R131 VSUBS.n57 VSUBS.t4 292.5
R132 VSUBS.n58 VSUBS.n56 292.5
R133 VSUBS.n56 VSUBS.t4 292.5
R134 VSUBS.n74 VSUBS.n71 292.5
R135 VSUBS.n71 VSUBS.t6 292.5
R136 VSUBS.n72 VSUBS.n70 292.5
R137 VSUBS.n70 VSUBS.t6 292.5
R138 VSUBS.n88 VSUBS.n85 292.5
R139 VSUBS.n85 VSUBS.t1 292.5
R140 VSUBS.n86 VSUBS.n84 292.5
R141 VSUBS.n84 VSUBS.t1 292.5
R142 VSUBS.n102 VSUBS.n99 292.5
R143 VSUBS.n99 VSUBS.t3 292.5
R144 VSUBS.n100 VSUBS.n98 292.5
R145 VSUBS.n98 VSUBS.t3 292.5
R146 VSUBS.n116 VSUBS.n113 292.5
R147 VSUBS.n113 VSUBS.t7 292.5
R148 VSUBS.n114 VSUBS.n112 292.5
R149 VSUBS.n112 VSUBS.t7 292.5
R150 VSUBS.n130 VSUBS.n127 292.5
R151 VSUBS.n127 VSUBS.t5 292.5
R152 VSUBS.n128 VSUBS.n126 292.5
R153 VSUBS.n126 VSUBS.t5 292.5
R154 VSUBS.n38 VSUBS.n33 292.5
R155 VSUBS.n33 VSUBS.t2 292.5
R156 VSUBS.n34 VSUBS.n32 292.5
R157 VSUBS.n52 VSUBS.n30 292.5
R158 VSUBS.n30 VSUBS.t0 292.5
R159 VSUBS.n31 VSUBS.n29 292.5
R160 VSUBS.n29 VSUBS.t0 292.5
R161 VSUBS.n66 VSUBS.n26 292.5
R162 VSUBS.n26 VSUBS.t4 292.5
R163 VSUBS.n27 VSUBS.n25 292.5
R164 VSUBS.n25 VSUBS.t4 292.5
R165 VSUBS.n80 VSUBS.n22 292.5
R166 VSUBS.n22 VSUBS.t6 292.5
R167 VSUBS.n23 VSUBS.n21 292.5
R168 VSUBS.n21 VSUBS.t6 292.5
R169 VSUBS.n94 VSUBS.n18 292.5
R170 VSUBS.n18 VSUBS.t1 292.5
R171 VSUBS.n19 VSUBS.n17 292.5
R172 VSUBS.n17 VSUBS.t1 292.5
R173 VSUBS.n108 VSUBS.n14 292.5
R174 VSUBS.n14 VSUBS.t3 292.5
R175 VSUBS.n15 VSUBS.n13 292.5
R176 VSUBS.n13 VSUBS.t3 292.5
R177 VSUBS.n122 VSUBS.n10 292.5
R178 VSUBS.n10 VSUBS.t7 292.5
R179 VSUBS.n11 VSUBS.n9 292.5
R180 VSUBS.n9 VSUBS.t7 292.5
R181 VSUBS.n136 VSUBS.n6 292.5
R182 VSUBS.n6 VSUBS.t5 292.5
R183 VSUBS.n7 VSUBS.n5 292.5
R184 VSUBS.n5 VSUBS.t5 292.5
R185 VSUBS.n142 VSUBS.n141 292.5
R186 VSUBS.n145 VSUBS.n144 292.5
R187 VSUBS.n144 VSUBS.t8 292.5
R188 VSUBS.n35 VSUBS.n32 288.877
R189 VSUBS.n143 VSUBS.n142 288.877
R190 VSUBS.n146 VSUBS.n145 269.93
R191 VSUBS.n140 VSUBS.n139 145.895
R192 VSUBS.n49 VSUBS.n41 88.0005
R193 VSUBS.n63 VSUBS.n55 88.0005
R194 VSUBS.n77 VSUBS.n69 88.0005
R195 VSUBS.n91 VSUBS.n83 88.0005
R196 VSUBS.n105 VSUBS.n97 88.0005
R197 VSUBS.n119 VSUBS.n111 88.0005
R198 VSUBS.n133 VSUBS.n125 88.0005
R199 VSUBS.n36 VSUBS.n35 46.7228
R200 VSUBS.n143 VSUBS.n3 46.7228
R201 VSUBS.n41 VSUBS.t2 42.8426
R202 VSUBS.n49 VSUBS.t0 42.8426
R203 VSUBS.n55 VSUBS.t0 42.8426
R204 VSUBS.n63 VSUBS.t4 42.8426
R205 VSUBS.n69 VSUBS.t4 42.8426
R206 VSUBS.n77 VSUBS.t6 42.8426
R207 VSUBS.n83 VSUBS.t6 42.8426
R208 VSUBS.n91 VSUBS.t1 42.8426
R209 VSUBS.n97 VSUBS.t1 42.8426
R210 VSUBS.n105 VSUBS.t3 42.8426
R211 VSUBS.n111 VSUBS.t3 42.8426
R212 VSUBS.n119 VSUBS.t7 42.8426
R213 VSUBS.n125 VSUBS.t7 42.8426
R214 VSUBS.n133 VSUBS.t5 42.8426
R215 VSUBS.n139 VSUBS.t5 42.8426
R216 VSUBS.t8 VSUBS.n140 42.8426
R217 VSUBS.n45 VSUBS.n28 8.0142
R218 VSUBS.n55 VSUBS.n28 8.0142
R219 VSUBS.n48 VSUBS.n47 8.0142
R220 VSUBS.n49 VSUBS.n48 8.0142
R221 VSUBS.n59 VSUBS.n24 8.0142
R222 VSUBS.n69 VSUBS.n24 8.0142
R223 VSUBS.n62 VSUBS.n61 8.0142
R224 VSUBS.n63 VSUBS.n62 8.0142
R225 VSUBS.n73 VSUBS.n20 8.0142
R226 VSUBS.n83 VSUBS.n20 8.0142
R227 VSUBS.n76 VSUBS.n75 8.0142
R228 VSUBS.n77 VSUBS.n76 8.0142
R229 VSUBS.n87 VSUBS.n16 8.0142
R230 VSUBS.n97 VSUBS.n16 8.0142
R231 VSUBS.n90 VSUBS.n89 8.0142
R232 VSUBS.n91 VSUBS.n90 8.0142
R233 VSUBS.n101 VSUBS.n12 8.0142
R234 VSUBS.n111 VSUBS.n12 8.0142
R235 VSUBS.n104 VSUBS.n103 8.0142
R236 VSUBS.n105 VSUBS.n104 8.0142
R237 VSUBS.n115 VSUBS.n8 8.0142
R238 VSUBS.n125 VSUBS.n8 8.0142
R239 VSUBS.n118 VSUBS.n117 8.0142
R240 VSUBS.n119 VSUBS.n118 8.0142
R241 VSUBS.n129 VSUBS.n4 8.0142
R242 VSUBS.n139 VSUBS.n4 8.0142
R243 VSUBS.n132 VSUBS.n131 8.0142
R244 VSUBS.n133 VSUBS.n132 8.0142
R245 VSUBS.n40 VSUBS.n39 4.46615
R246 VSUBS.n41 VSUBS.n40 4.46615
R247 VSUBS.n37 VSUBS.n36 4.46615
R248 VSUBS.n54 VSUBS.n53 4.46615
R249 VSUBS.n55 VSUBS.n54 4.46615
R250 VSUBS.n51 VSUBS.n50 4.46615
R251 VSUBS.n50 VSUBS.n49 4.46615
R252 VSUBS.n68 VSUBS.n67 4.46615
R253 VSUBS.n69 VSUBS.n68 4.46615
R254 VSUBS.n65 VSUBS.n64 4.46615
R255 VSUBS.n64 VSUBS.n63 4.46615
R256 VSUBS.n82 VSUBS.n81 4.46615
R257 VSUBS.n83 VSUBS.n82 4.46615
R258 VSUBS.n79 VSUBS.n78 4.46615
R259 VSUBS.n78 VSUBS.n77 4.46615
R260 VSUBS.n96 VSUBS.n95 4.46615
R261 VSUBS.n97 VSUBS.n96 4.46615
R262 VSUBS.n93 VSUBS.n92 4.46615
R263 VSUBS.n92 VSUBS.n91 4.46615
R264 VSUBS.n110 VSUBS.n109 4.46615
R265 VSUBS.n111 VSUBS.n110 4.46615
R266 VSUBS.n107 VSUBS.n106 4.46615
R267 VSUBS.n106 VSUBS.n105 4.46615
R268 VSUBS.n124 VSUBS.n123 4.46615
R269 VSUBS.n125 VSUBS.n124 4.46615
R270 VSUBS.n121 VSUBS.n120 4.46615
R271 VSUBS.n120 VSUBS.n119 4.46615
R272 VSUBS.n138 VSUBS.n137 4.46615
R273 VSUBS.n139 VSUBS.n138 4.46615
R274 VSUBS.n135 VSUBS.n134 4.46615
R275 VSUBS.n134 VSUBS.n133 4.46615
R276 VSUBS.n3 VSUBS.n0 4.46615
R277 VSUBS.n2 VSUBS.n1 4.46615
R278 VSUBS.n140 VSUBS.n2 4.46615
R279 VSUBS VSUBS.n146 1.39508
R280 VSUBS.n35 VSUBS.t2 0.50541
R281 VSUBS.t8 VSUBS.n143 0.50541
C0 a_n1034_2566# a_n434_6998# 0.131455f
C1 a_n1034_2566# GND 0.023658f
C2 out a_1366_2566# 0.151801f
C3 a_1966_6998# a_1366_2566# 0.131485f
C4 b5 b6 0.098267f
C5 out a_1966_6998# 0.106769f
C6 b7 b6 0.098267f
C7 a_n1834_10998# a_n434_6998# 1.8e-21
C8 b5 b4 0.098267f
C9 a_n1034_2566# a_n1834_10998# 0.20932f
C10 b3 b2 0.098267f
C11 a_766_6998# a_166_2566# 0.131455f
C12 a_n434_6998# a_166_2566# 0.209322f
C13 b3 b4 0.098267f
C14 b1 b2 0.098267f
C15 b1 b0 0.098267f
C16 a_n1034_2566# a_166_2566# 0.182372f
C17 a_166_2566# a_1366_2566# 0.182372f
C18 a_766_6998# a_1366_2566# 0.209322f
.ends

