magic
tech sky130A
magscale 1 2
timestamp 1708085196
<< viali >>
rect 6837 3689 6871 3723
rect 6377 3553 6411 3587
rect 6561 3553 6595 3587
rect 10793 3553 10827 3587
rect 6285 3485 6319 3519
rect 6469 3485 6503 3519
rect 8125 3485 8159 3519
rect 8401 3485 8435 3519
rect 6101 3349 6135 3383
rect 10609 3349 10643 3383
rect 7849 3145 7883 3179
rect 4077 2941 4111 2975
rect 4353 2941 4387 2975
rect 5825 2941 5859 2975
rect 7665 2941 7699 2975
rect 9045 2941 9079 2975
rect 5641 2805 5675 2839
rect 7113 2805 7147 2839
rect 8125 2805 8159 2839
rect 8953 2805 8987 2839
rect 4721 2601 4755 2635
rect 6745 2601 6779 2635
rect 7113 2601 7147 2635
rect 8585 2533 8619 2567
rect 3893 2465 3927 2499
rect 4077 2465 4111 2499
rect 4997 2465 5031 2499
rect 5549 2465 5583 2499
rect 6653 2465 6687 2499
rect 6856 2465 6890 2499
rect 3801 2397 3835 2431
rect 3985 2397 4019 2431
rect 4353 2397 4387 2431
rect 6469 2397 6503 2431
rect 7021 2397 7055 2431
rect 8861 2397 8895 2431
rect 4905 2329 4939 2363
rect 6745 2329 6779 2363
rect 4261 2261 4295 2295
rect 4721 2261 4755 2295
rect 5917 2261 5951 2295
rect 4353 1989 4387 2023
rect 4537 1921 4571 1955
rect 4721 1921 4755 1955
rect 4077 1853 4111 1887
rect 4445 1853 4479 1887
rect 4629 1853 4663 1887
rect 4997 1853 5031 1887
rect 7481 1853 7515 1887
rect 4353 1785 4387 1819
rect 4169 1717 4203 1751
rect 6101 1717 6135 1751
rect 7297 1717 7331 1751
rect 5181 1513 5215 1547
rect 5825 1445 5859 1479
rect 5365 1377 5399 1411
rect 6009 1377 6043 1411
rect 6101 1377 6135 1411
rect 5549 1309 5583 1343
rect 5641 1309 5675 1343
rect 7665 1309 7699 1343
rect 7941 1309 7975 1343
rect 5825 1241 5859 1275
rect 6561 1173 6595 1207
rect 3709 969 3743 1003
rect 7205 969 7239 1003
rect 9689 969 9723 1003
rect 6653 833 6687 867
rect 7389 833 7423 867
rect 7297 765 7331 799
rect 7481 765 7515 799
rect 4997 697 5031 731
rect 8401 697 8435 731
<< metal1 >>
rect 552 11450 11568 11472
rect 552 11398 3112 11450
rect 3164 11398 3176 11450
rect 3228 11398 3240 11450
rect 3292 11398 3304 11450
rect 3356 11398 3368 11450
rect 3420 11398 5826 11450
rect 5878 11398 5890 11450
rect 5942 11398 5954 11450
rect 6006 11398 6018 11450
rect 6070 11398 6082 11450
rect 6134 11398 8540 11450
rect 8592 11398 8604 11450
rect 8656 11398 8668 11450
rect 8720 11398 8732 11450
rect 8784 11398 8796 11450
rect 8848 11398 11254 11450
rect 11306 11398 11318 11450
rect 11370 11398 11382 11450
rect 11434 11398 11446 11450
rect 11498 11398 11510 11450
rect 11562 11398 11568 11450
rect 552 11376 11568 11398
rect 552 10906 11408 10928
rect 552 10854 1755 10906
rect 1807 10854 1819 10906
rect 1871 10854 1883 10906
rect 1935 10854 1947 10906
rect 1999 10854 2011 10906
rect 2063 10854 4469 10906
rect 4521 10854 4533 10906
rect 4585 10854 4597 10906
rect 4649 10854 4661 10906
rect 4713 10854 4725 10906
rect 4777 10854 7183 10906
rect 7235 10854 7247 10906
rect 7299 10854 7311 10906
rect 7363 10854 7375 10906
rect 7427 10854 7439 10906
rect 7491 10854 9897 10906
rect 9949 10854 9961 10906
rect 10013 10854 10025 10906
rect 10077 10854 10089 10906
rect 10141 10854 10153 10906
rect 10205 10854 11408 10906
rect 552 10832 11408 10854
rect 552 10362 11568 10384
rect 552 10310 3112 10362
rect 3164 10310 3176 10362
rect 3228 10310 3240 10362
rect 3292 10310 3304 10362
rect 3356 10310 3368 10362
rect 3420 10310 5826 10362
rect 5878 10310 5890 10362
rect 5942 10310 5954 10362
rect 6006 10310 6018 10362
rect 6070 10310 6082 10362
rect 6134 10310 8540 10362
rect 8592 10310 8604 10362
rect 8656 10310 8668 10362
rect 8720 10310 8732 10362
rect 8784 10310 8796 10362
rect 8848 10310 11254 10362
rect 11306 10310 11318 10362
rect 11370 10310 11382 10362
rect 11434 10310 11446 10362
rect 11498 10310 11510 10362
rect 11562 10310 11568 10362
rect 552 10288 11568 10310
rect 552 9818 11408 9840
rect 552 9766 1755 9818
rect 1807 9766 1819 9818
rect 1871 9766 1883 9818
rect 1935 9766 1947 9818
rect 1999 9766 2011 9818
rect 2063 9766 4469 9818
rect 4521 9766 4533 9818
rect 4585 9766 4597 9818
rect 4649 9766 4661 9818
rect 4713 9766 4725 9818
rect 4777 9766 7183 9818
rect 7235 9766 7247 9818
rect 7299 9766 7311 9818
rect 7363 9766 7375 9818
rect 7427 9766 7439 9818
rect 7491 9766 9897 9818
rect 9949 9766 9961 9818
rect 10013 9766 10025 9818
rect 10077 9766 10089 9818
rect 10141 9766 10153 9818
rect 10205 9766 11408 9818
rect 552 9744 11408 9766
rect 552 9274 11568 9296
rect 552 9222 3112 9274
rect 3164 9222 3176 9274
rect 3228 9222 3240 9274
rect 3292 9222 3304 9274
rect 3356 9222 3368 9274
rect 3420 9222 5826 9274
rect 5878 9222 5890 9274
rect 5942 9222 5954 9274
rect 6006 9222 6018 9274
rect 6070 9222 6082 9274
rect 6134 9222 8540 9274
rect 8592 9222 8604 9274
rect 8656 9222 8668 9274
rect 8720 9222 8732 9274
rect 8784 9222 8796 9274
rect 8848 9222 11254 9274
rect 11306 9222 11318 9274
rect 11370 9222 11382 9274
rect 11434 9222 11446 9274
rect 11498 9222 11510 9274
rect 11562 9222 11568 9274
rect 552 9200 11568 9222
rect 552 8730 11408 8752
rect 552 8678 1755 8730
rect 1807 8678 1819 8730
rect 1871 8678 1883 8730
rect 1935 8678 1947 8730
rect 1999 8678 2011 8730
rect 2063 8678 4469 8730
rect 4521 8678 4533 8730
rect 4585 8678 4597 8730
rect 4649 8678 4661 8730
rect 4713 8678 4725 8730
rect 4777 8678 7183 8730
rect 7235 8678 7247 8730
rect 7299 8678 7311 8730
rect 7363 8678 7375 8730
rect 7427 8678 7439 8730
rect 7491 8678 9897 8730
rect 9949 8678 9961 8730
rect 10013 8678 10025 8730
rect 10077 8678 10089 8730
rect 10141 8678 10153 8730
rect 10205 8678 11408 8730
rect 552 8656 11408 8678
rect 552 8186 11568 8208
rect 552 8134 3112 8186
rect 3164 8134 3176 8186
rect 3228 8134 3240 8186
rect 3292 8134 3304 8186
rect 3356 8134 3368 8186
rect 3420 8134 5826 8186
rect 5878 8134 5890 8186
rect 5942 8134 5954 8186
rect 6006 8134 6018 8186
rect 6070 8134 6082 8186
rect 6134 8134 8540 8186
rect 8592 8134 8604 8186
rect 8656 8134 8668 8186
rect 8720 8134 8732 8186
rect 8784 8134 8796 8186
rect 8848 8134 11254 8186
rect 11306 8134 11318 8186
rect 11370 8134 11382 8186
rect 11434 8134 11446 8186
rect 11498 8134 11510 8186
rect 11562 8134 11568 8186
rect 552 8112 11568 8134
rect 552 7642 11408 7664
rect 552 7590 1755 7642
rect 1807 7590 1819 7642
rect 1871 7590 1883 7642
rect 1935 7590 1947 7642
rect 1999 7590 2011 7642
rect 2063 7590 4469 7642
rect 4521 7590 4533 7642
rect 4585 7590 4597 7642
rect 4649 7590 4661 7642
rect 4713 7590 4725 7642
rect 4777 7590 7183 7642
rect 7235 7590 7247 7642
rect 7299 7590 7311 7642
rect 7363 7590 7375 7642
rect 7427 7590 7439 7642
rect 7491 7590 9897 7642
rect 9949 7590 9961 7642
rect 10013 7590 10025 7642
rect 10077 7590 10089 7642
rect 10141 7590 10153 7642
rect 10205 7590 11408 7642
rect 552 7568 11408 7590
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 5534 7528 5540 7540
rect 2832 7500 5540 7528
rect 2832 7488 2838 7500
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 552 7098 11568 7120
rect 552 7046 3112 7098
rect 3164 7046 3176 7098
rect 3228 7046 3240 7098
rect 3292 7046 3304 7098
rect 3356 7046 3368 7098
rect 3420 7046 5826 7098
rect 5878 7046 5890 7098
rect 5942 7046 5954 7098
rect 6006 7046 6018 7098
rect 6070 7046 6082 7098
rect 6134 7046 8540 7098
rect 8592 7046 8604 7098
rect 8656 7046 8668 7098
rect 8720 7046 8732 7098
rect 8784 7046 8796 7098
rect 8848 7046 11254 7098
rect 11306 7046 11318 7098
rect 11370 7046 11382 7098
rect 11434 7046 11446 7098
rect 11498 7046 11510 7098
rect 11562 7046 11568 7098
rect 552 7024 11568 7046
rect 552 6554 11408 6576
rect 552 6502 1755 6554
rect 1807 6502 1819 6554
rect 1871 6502 1883 6554
rect 1935 6502 1947 6554
rect 1999 6502 2011 6554
rect 2063 6502 4469 6554
rect 4521 6502 4533 6554
rect 4585 6502 4597 6554
rect 4649 6502 4661 6554
rect 4713 6502 4725 6554
rect 4777 6502 7183 6554
rect 7235 6502 7247 6554
rect 7299 6502 7311 6554
rect 7363 6502 7375 6554
rect 7427 6502 7439 6554
rect 7491 6502 9897 6554
rect 9949 6502 9961 6554
rect 10013 6502 10025 6554
rect 10077 6502 10089 6554
rect 10141 6502 10153 6554
rect 10205 6502 11408 6554
rect 552 6480 11408 6502
rect 552 6010 11568 6032
rect 552 5958 3112 6010
rect 3164 5958 3176 6010
rect 3228 5958 3240 6010
rect 3292 5958 3304 6010
rect 3356 5958 3368 6010
rect 3420 5958 5826 6010
rect 5878 5958 5890 6010
rect 5942 5958 5954 6010
rect 6006 5958 6018 6010
rect 6070 5958 6082 6010
rect 6134 5958 8540 6010
rect 8592 5958 8604 6010
rect 8656 5958 8668 6010
rect 8720 5958 8732 6010
rect 8784 5958 8796 6010
rect 8848 5958 11254 6010
rect 11306 5958 11318 6010
rect 11370 5958 11382 6010
rect 11434 5958 11446 6010
rect 11498 5958 11510 6010
rect 11562 5958 11568 6010
rect 552 5936 11568 5958
rect 552 5466 11408 5488
rect 552 5414 1755 5466
rect 1807 5414 1819 5466
rect 1871 5414 1883 5466
rect 1935 5414 1947 5466
rect 1999 5414 2011 5466
rect 2063 5414 4469 5466
rect 4521 5414 4533 5466
rect 4585 5414 4597 5466
rect 4649 5414 4661 5466
rect 4713 5414 4725 5466
rect 4777 5414 7183 5466
rect 7235 5414 7247 5466
rect 7299 5414 7311 5466
rect 7363 5414 7375 5466
rect 7427 5414 7439 5466
rect 7491 5414 9897 5466
rect 9949 5414 9961 5466
rect 10013 5414 10025 5466
rect 10077 5414 10089 5466
rect 10141 5414 10153 5466
rect 10205 5414 11408 5466
rect 552 5392 11408 5414
rect 552 4922 11568 4944
rect 552 4870 3112 4922
rect 3164 4870 3176 4922
rect 3228 4870 3240 4922
rect 3292 4870 3304 4922
rect 3356 4870 3368 4922
rect 3420 4870 5826 4922
rect 5878 4870 5890 4922
rect 5942 4870 5954 4922
rect 6006 4870 6018 4922
rect 6070 4870 6082 4922
rect 6134 4870 8540 4922
rect 8592 4870 8604 4922
rect 8656 4870 8668 4922
rect 8720 4870 8732 4922
rect 8784 4870 8796 4922
rect 8848 4870 11254 4922
rect 11306 4870 11318 4922
rect 11370 4870 11382 4922
rect 11434 4870 11446 4922
rect 11498 4870 11510 4922
rect 11562 4870 11568 4922
rect 552 4848 11568 4870
rect 552 4378 11408 4400
rect 552 4326 1755 4378
rect 1807 4326 1819 4378
rect 1871 4326 1883 4378
rect 1935 4326 1947 4378
rect 1999 4326 2011 4378
rect 2063 4326 4469 4378
rect 4521 4326 4533 4378
rect 4585 4326 4597 4378
rect 4649 4326 4661 4378
rect 4713 4326 4725 4378
rect 4777 4326 7183 4378
rect 7235 4326 7247 4378
rect 7299 4326 7311 4378
rect 7363 4326 7375 4378
rect 7427 4326 7439 4378
rect 7491 4326 9897 4378
rect 9949 4326 9961 4378
rect 10013 4326 10025 4378
rect 10077 4326 10089 4378
rect 10141 4326 10153 4378
rect 10205 4326 11408 4378
rect 552 4304 11408 4326
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 11606 4128 11612 4140
rect 6880 4100 11612 4128
rect 6880 4088 6886 4100
rect 11606 4088 11612 4100
rect 11664 4088 11670 4140
rect 552 3834 11568 3856
rect 552 3782 3112 3834
rect 3164 3782 3176 3834
rect 3228 3782 3240 3834
rect 3292 3782 3304 3834
rect 3356 3782 3368 3834
rect 3420 3782 5826 3834
rect 5878 3782 5890 3834
rect 5942 3782 5954 3834
rect 6006 3782 6018 3834
rect 6070 3782 6082 3834
rect 6134 3782 8540 3834
rect 8592 3782 8604 3834
rect 8656 3782 8668 3834
rect 8720 3782 8732 3834
rect 8784 3782 8796 3834
rect 8848 3782 11254 3834
rect 11306 3782 11318 3834
rect 11370 3782 11382 3834
rect 11434 3782 11446 3834
rect 11498 3782 11510 3834
rect 11562 3782 11568 3834
rect 552 3760 11568 3782
rect 6822 3680 6828 3732
rect 6880 3680 6886 3732
rect 6270 3612 6276 3664
rect 6328 3612 6334 3664
rect 6288 3584 6316 3612
rect 6365 3587 6423 3593
rect 6365 3584 6377 3587
rect 6288 3556 6377 3584
rect 6365 3553 6377 3556
rect 6411 3553 6423 3587
rect 6365 3547 6423 3553
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 6840 3584 6868 3680
rect 6595 3556 6868 3584
rect 10781 3587 10839 3593
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 10781 3553 10793 3587
rect 10827 3553 10839 3587
rect 10781 3547 10839 3553
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 6273 3519 6331 3525
rect 6273 3516 6285 3519
rect 5776 3488 6285 3516
rect 5776 3476 5782 3488
rect 6273 3485 6285 3488
rect 6319 3485 6331 3519
rect 6273 3479 6331 3485
rect 6457 3519 6515 3525
rect 6457 3485 6469 3519
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 6472 3448 6500 3479
rect 8110 3476 8116 3528
rect 8168 3476 8174 3528
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 8938 3516 8944 3528
rect 8435 3488 8944 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 10796 3516 10824 3547
rect 11238 3516 11244 3528
rect 10796 3488 11244 3516
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 6380 3420 6500 3448
rect 6380 3392 6408 3420
rect 5626 3340 5632 3392
rect 5684 3380 5690 3392
rect 6089 3383 6147 3389
rect 6089 3380 6101 3383
rect 5684 3352 6101 3380
rect 5684 3340 5690 3352
rect 6089 3349 6101 3352
rect 6135 3349 6147 3383
rect 6089 3343 6147 3349
rect 6362 3340 6368 3392
rect 6420 3340 6426 3392
rect 10594 3340 10600 3392
rect 10652 3340 10658 3392
rect 552 3290 11408 3312
rect 552 3238 1755 3290
rect 1807 3238 1819 3290
rect 1871 3238 1883 3290
rect 1935 3238 1947 3290
rect 1999 3238 2011 3290
rect 2063 3238 4469 3290
rect 4521 3238 4533 3290
rect 4585 3238 4597 3290
rect 4649 3238 4661 3290
rect 4713 3238 4725 3290
rect 4777 3238 7183 3290
rect 7235 3238 7247 3290
rect 7299 3238 7311 3290
rect 7363 3238 7375 3290
rect 7427 3238 7439 3290
rect 7491 3238 9897 3290
rect 9949 3238 9961 3290
rect 10013 3238 10025 3290
rect 10077 3238 10089 3290
rect 10141 3238 10153 3290
rect 10205 3238 11408 3290
rect 552 3216 11408 3238
rect 7837 3179 7895 3185
rect 7837 3145 7849 3179
rect 7883 3176 7895 3179
rect 8110 3176 8116 3188
rect 7883 3148 8116 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 10594 3136 10600 3188
rect 10652 3136 10658 3188
rect 4065 2975 4123 2981
rect 4065 2972 4077 2975
rect 3712 2944 4077 2972
rect 3712 2848 3740 2944
rect 4065 2941 4077 2944
rect 4111 2941 4123 2975
rect 4065 2935 4123 2941
rect 4338 2932 4344 2984
rect 4396 2932 4402 2984
rect 5534 2932 5540 2984
rect 5592 2972 5598 2984
rect 5813 2975 5871 2981
rect 5813 2972 5825 2975
rect 5592 2944 5825 2972
rect 5592 2932 5598 2944
rect 5813 2941 5825 2944
rect 5859 2941 5871 2975
rect 5813 2935 5871 2941
rect 6178 2932 6184 2984
rect 6236 2972 6242 2984
rect 7653 2975 7711 2981
rect 7653 2972 7665 2975
rect 6236 2944 7665 2972
rect 6236 2932 6242 2944
rect 7653 2941 7665 2944
rect 7699 2941 7711 2975
rect 7653 2935 7711 2941
rect 9033 2975 9091 2981
rect 9033 2941 9045 2975
rect 9079 2972 9091 2975
rect 10612 2972 10640 3136
rect 9079 2944 10640 2972
rect 9079 2941 9091 2944
rect 9033 2935 9091 2941
rect 3694 2796 3700 2848
rect 3752 2796 3758 2848
rect 5534 2796 5540 2848
rect 5592 2836 5598 2848
rect 5629 2839 5687 2845
rect 5629 2836 5641 2839
rect 5592 2808 5641 2836
rect 5592 2796 5598 2808
rect 5629 2805 5641 2808
rect 5675 2836 5687 2839
rect 5718 2836 5724 2848
rect 5675 2808 5724 2836
rect 5675 2805 5687 2808
rect 5629 2799 5687 2805
rect 5718 2796 5724 2808
rect 5776 2836 5782 2848
rect 6730 2836 6736 2848
rect 5776 2808 6736 2836
rect 5776 2796 5782 2808
rect 6730 2796 6736 2808
rect 6788 2796 6794 2848
rect 7098 2796 7104 2848
rect 7156 2796 7162 2848
rect 8113 2839 8171 2845
rect 8113 2805 8125 2839
rect 8159 2836 8171 2839
rect 8294 2836 8300 2848
rect 8159 2808 8300 2836
rect 8159 2805 8171 2808
rect 8113 2799 8171 2805
rect 8294 2796 8300 2808
rect 8352 2796 8358 2848
rect 8386 2796 8392 2848
rect 8444 2836 8450 2848
rect 8941 2839 8999 2845
rect 8941 2836 8953 2839
rect 8444 2808 8953 2836
rect 8444 2796 8450 2808
rect 8941 2805 8953 2808
rect 8987 2805 8999 2839
rect 8941 2799 8999 2805
rect 552 2746 11568 2768
rect 552 2694 3112 2746
rect 3164 2694 3176 2746
rect 3228 2694 3240 2746
rect 3292 2694 3304 2746
rect 3356 2694 3368 2746
rect 3420 2694 5826 2746
rect 5878 2694 5890 2746
rect 5942 2694 5954 2746
rect 6006 2694 6018 2746
rect 6070 2694 6082 2746
rect 6134 2694 8540 2746
rect 8592 2694 8604 2746
rect 8656 2694 8668 2746
rect 8720 2694 8732 2746
rect 8784 2694 8796 2746
rect 8848 2694 11254 2746
rect 11306 2694 11318 2746
rect 11370 2694 11382 2746
rect 11434 2694 11446 2746
rect 11498 2694 11510 2746
rect 11562 2694 11568 2746
rect 552 2672 11568 2694
rect 4709 2635 4767 2641
rect 4709 2601 4721 2635
rect 4755 2632 4767 2635
rect 5626 2632 5632 2644
rect 4755 2604 5632 2632
rect 4755 2601 4767 2604
rect 4709 2595 4767 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 6730 2592 6736 2644
rect 6788 2592 6794 2644
rect 7101 2635 7159 2641
rect 7101 2601 7113 2635
rect 7147 2601 7159 2635
rect 8386 2632 8392 2644
rect 7101 2595 7159 2601
rect 8220 2604 8392 2632
rect 7006 2564 7012 2576
rect 3896 2536 4200 2564
rect 3896 2505 3924 2536
rect 3881 2499 3939 2505
rect 3881 2465 3893 2499
rect 3927 2465 3939 2499
rect 3881 2459 3939 2465
rect 4062 2456 4068 2508
rect 4120 2456 4126 2508
rect 3786 2388 3792 2440
rect 3844 2388 3850 2440
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2428 4031 2431
rect 4019 2400 4108 2428
rect 4019 2397 4031 2400
rect 3973 2391 4031 2397
rect 4080 2304 4108 2400
rect 4172 2304 4200 2536
rect 4356 2536 7012 2564
rect 4356 2437 4384 2536
rect 7006 2524 7012 2536
rect 7064 2564 7070 2576
rect 7116 2564 7144 2595
rect 8220 2564 8248 2604
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 7064 2536 7144 2564
rect 8142 2536 8248 2564
rect 7064 2524 7070 2536
rect 8294 2524 8300 2576
rect 8352 2564 8358 2576
rect 8573 2567 8631 2573
rect 8573 2564 8585 2567
rect 8352 2536 8585 2564
rect 8352 2524 8358 2536
rect 8573 2533 8585 2536
rect 8619 2533 8631 2567
rect 8573 2527 8631 2533
rect 4890 2456 4896 2508
rect 4948 2496 4954 2508
rect 4985 2499 5043 2505
rect 4985 2496 4997 2499
rect 4948 2468 4997 2496
rect 4948 2456 4954 2468
rect 4985 2465 4997 2468
rect 5031 2465 5043 2499
rect 4985 2459 5043 2465
rect 5534 2456 5540 2508
rect 5592 2456 5598 2508
rect 6178 2456 6184 2508
rect 6236 2456 6242 2508
rect 6638 2456 6644 2508
rect 6696 2456 6702 2508
rect 6844 2499 6902 2505
rect 6844 2496 6856 2499
rect 6840 2465 6856 2496
rect 6890 2465 6902 2499
rect 6840 2459 6902 2465
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2397 4399 2431
rect 6196 2428 6224 2456
rect 4341 2391 4399 2397
rect 4908 2400 6224 2428
rect 4908 2369 4936 2400
rect 6270 2388 6276 2440
rect 6328 2428 6334 2440
rect 6457 2431 6515 2437
rect 6457 2428 6469 2431
rect 6328 2400 6469 2428
rect 6328 2388 6334 2400
rect 6457 2397 6469 2400
rect 6503 2428 6515 2431
rect 6840 2428 6868 2459
rect 6503 2400 6868 2428
rect 7009 2431 7067 2437
rect 6503 2397 6515 2400
rect 6457 2391 6515 2397
rect 7009 2397 7021 2431
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 8849 2431 8907 2437
rect 8849 2397 8861 2431
rect 8895 2428 8907 2431
rect 8938 2428 8944 2440
rect 8895 2400 8944 2428
rect 8895 2397 8907 2400
rect 8849 2391 8907 2397
rect 4893 2363 4951 2369
rect 4893 2329 4905 2363
rect 4939 2329 4951 2363
rect 6733 2363 6791 2369
rect 6733 2360 6745 2363
rect 4893 2323 4951 2329
rect 5460 2332 6745 2360
rect 4062 2252 4068 2304
rect 4120 2252 4126 2304
rect 4154 2252 4160 2304
rect 4212 2252 4218 2304
rect 4246 2252 4252 2304
rect 4304 2252 4310 2304
rect 4709 2295 4767 2301
rect 4709 2261 4721 2295
rect 4755 2292 4767 2295
rect 5460 2292 5488 2332
rect 6733 2329 6745 2332
rect 6779 2329 6791 2363
rect 7024 2360 7052 2391
rect 8938 2388 8944 2400
rect 8996 2388 9002 2440
rect 6733 2323 6791 2329
rect 6840 2332 7052 2360
rect 6840 2304 6868 2332
rect 4755 2264 5488 2292
rect 4755 2261 4767 2264
rect 4709 2255 4767 2261
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 5905 2295 5963 2301
rect 5905 2292 5917 2295
rect 5592 2264 5917 2292
rect 5592 2252 5598 2264
rect 5905 2261 5917 2264
rect 5951 2261 5963 2295
rect 5905 2255 5963 2261
rect 6362 2252 6368 2304
rect 6420 2292 6426 2304
rect 6822 2292 6828 2304
rect 6420 2264 6828 2292
rect 6420 2252 6426 2264
rect 6822 2252 6828 2264
rect 6880 2252 6886 2304
rect 552 2202 11408 2224
rect 552 2150 1755 2202
rect 1807 2150 1819 2202
rect 1871 2150 1883 2202
rect 1935 2150 1947 2202
rect 1999 2150 2011 2202
rect 2063 2150 4469 2202
rect 4521 2150 4533 2202
rect 4585 2150 4597 2202
rect 4649 2150 4661 2202
rect 4713 2150 4725 2202
rect 4777 2150 7183 2202
rect 7235 2150 7247 2202
rect 7299 2150 7311 2202
rect 7363 2150 7375 2202
rect 7427 2150 7439 2202
rect 7491 2150 9897 2202
rect 9949 2150 9961 2202
rect 10013 2150 10025 2202
rect 10077 2150 10089 2202
rect 10141 2150 10153 2202
rect 10205 2150 11408 2202
rect 552 2128 11408 2150
rect 3712 2060 4752 2088
rect 3712 2032 3740 2060
rect 3694 1980 3700 2032
rect 3752 1980 3758 2032
rect 4341 2023 4399 2029
rect 4341 1989 4353 2023
rect 4387 2020 4399 2023
rect 4387 1992 4660 2020
rect 4387 1989 4399 1992
rect 4341 1983 4399 1989
rect 4522 1912 4528 1964
rect 4580 1912 4586 1964
rect 4062 1844 4068 1896
rect 4120 1844 4126 1896
rect 4246 1844 4252 1896
rect 4304 1884 4310 1896
rect 4632 1893 4660 1992
rect 4724 1961 4752 2060
rect 7006 2048 7012 2100
rect 7064 2048 7070 2100
rect 4709 1955 4767 1961
rect 4709 1921 4721 1955
rect 4755 1921 4767 1955
rect 4709 1915 4767 1921
rect 4890 1912 4896 1964
rect 4948 1912 4954 1964
rect 4433 1887 4491 1893
rect 4433 1884 4445 1887
rect 4304 1856 4445 1884
rect 4304 1844 4310 1856
rect 4433 1853 4445 1856
rect 4479 1853 4491 1887
rect 4433 1847 4491 1853
rect 4617 1887 4675 1893
rect 4617 1853 4629 1887
rect 4663 1853 4675 1887
rect 4908 1884 4936 1912
rect 4617 1847 4675 1853
rect 4724 1856 4936 1884
rect 14 1776 20 1828
rect 72 1816 78 1828
rect 4080 1816 4108 1844
rect 4341 1819 4399 1825
rect 72 1788 4292 1816
rect 72 1776 78 1788
rect 4154 1708 4160 1760
rect 4212 1708 4218 1760
rect 4264 1748 4292 1788
rect 4341 1785 4353 1819
rect 4387 1816 4399 1819
rect 4724 1816 4752 1856
rect 4982 1844 4988 1896
rect 5040 1844 5046 1896
rect 7024 1884 7052 2048
rect 7469 1887 7527 1893
rect 7469 1884 7481 1887
rect 7024 1856 7481 1884
rect 7469 1853 7481 1856
rect 7515 1853 7527 1887
rect 7469 1847 7527 1853
rect 4387 1788 4752 1816
rect 4387 1785 4399 1788
rect 4341 1779 4399 1785
rect 6089 1751 6147 1757
rect 6089 1748 6101 1751
rect 4264 1720 6101 1748
rect 6089 1717 6101 1720
rect 6135 1748 6147 1751
rect 6178 1748 6184 1760
rect 6135 1720 6184 1748
rect 6135 1717 6147 1720
rect 6089 1711 6147 1717
rect 6178 1708 6184 1720
rect 6236 1708 6242 1760
rect 6914 1708 6920 1760
rect 6972 1748 6978 1760
rect 7285 1751 7343 1757
rect 7285 1748 7297 1751
rect 6972 1720 7297 1748
rect 6972 1708 6978 1720
rect 7285 1717 7297 1720
rect 7331 1717 7343 1751
rect 7285 1711 7343 1717
rect 552 1658 11568 1680
rect 552 1606 3112 1658
rect 3164 1606 3176 1658
rect 3228 1606 3240 1658
rect 3292 1606 3304 1658
rect 3356 1606 3368 1658
rect 3420 1606 5826 1658
rect 5878 1606 5890 1658
rect 5942 1606 5954 1658
rect 6006 1606 6018 1658
rect 6070 1606 6082 1658
rect 6134 1606 8540 1658
rect 8592 1606 8604 1658
rect 8656 1606 8668 1658
rect 8720 1606 8732 1658
rect 8784 1606 8796 1658
rect 8848 1606 11254 1658
rect 11306 1606 11318 1658
rect 11370 1606 11382 1658
rect 11434 1606 11446 1658
rect 11498 1606 11510 1658
rect 11562 1606 11568 1658
rect 552 1584 11568 1606
rect 3786 1504 3792 1556
rect 3844 1504 3850 1556
rect 4982 1504 4988 1556
rect 5040 1544 5046 1556
rect 5169 1547 5227 1553
rect 5169 1544 5181 1547
rect 5040 1516 5181 1544
rect 5040 1504 5046 1516
rect 5169 1513 5181 1516
rect 5215 1513 5227 1547
rect 5169 1507 5227 1513
rect 3804 1476 3832 1504
rect 5813 1479 5871 1485
rect 5813 1476 5825 1479
rect 3804 1448 5825 1476
rect 5813 1445 5825 1448
rect 5859 1476 5871 1479
rect 6914 1476 6920 1488
rect 5859 1448 6920 1476
rect 5859 1445 5871 1448
rect 5813 1439 5871 1445
rect 6914 1436 6920 1448
rect 6972 1436 6978 1488
rect 4154 1368 4160 1420
rect 4212 1408 4218 1420
rect 5353 1411 5411 1417
rect 4212 1380 5304 1408
rect 4212 1368 4218 1380
rect 5276 1340 5304 1380
rect 5353 1377 5365 1411
rect 5399 1408 5411 1411
rect 5997 1411 6055 1417
rect 5399 1380 5948 1408
rect 5399 1377 5411 1380
rect 5353 1371 5411 1377
rect 5276 1312 5488 1340
rect 5460 1272 5488 1312
rect 5534 1300 5540 1352
rect 5592 1300 5598 1352
rect 5629 1343 5687 1349
rect 5629 1309 5641 1343
rect 5675 1309 5687 1343
rect 5629 1303 5687 1309
rect 5644 1272 5672 1303
rect 5460 1244 5672 1272
rect 5644 1204 5672 1244
rect 5813 1275 5871 1281
rect 5813 1241 5825 1275
rect 5859 1272 5871 1275
rect 5920 1272 5948 1380
rect 5997 1377 6009 1411
rect 6043 1377 6055 1411
rect 5997 1371 6055 1377
rect 6089 1411 6147 1417
rect 6089 1377 6101 1411
rect 6135 1408 6147 1411
rect 6178 1408 6184 1420
rect 6135 1380 6184 1408
rect 6135 1377 6147 1380
rect 6089 1371 6147 1377
rect 5859 1244 5948 1272
rect 6012 1340 6040 1371
rect 6178 1368 6184 1380
rect 6236 1368 6242 1420
rect 6012 1312 6592 1340
rect 5859 1241 5871 1244
rect 5813 1235 5871 1241
rect 6012 1204 6040 1312
rect 6564 1213 6592 1312
rect 7650 1300 7656 1352
rect 7708 1300 7714 1352
rect 7929 1343 7987 1349
rect 7929 1309 7941 1343
rect 7975 1340 7987 1343
rect 8846 1340 8852 1352
rect 7975 1312 8852 1340
rect 7975 1309 7987 1312
rect 7929 1303 7987 1309
rect 8846 1300 8852 1312
rect 8904 1300 8910 1352
rect 5644 1176 6040 1204
rect 6549 1207 6607 1213
rect 6549 1173 6561 1207
rect 6595 1204 6607 1207
rect 6822 1204 6828 1216
rect 6595 1176 6828 1204
rect 6595 1173 6607 1176
rect 6549 1167 6607 1173
rect 6822 1164 6828 1176
rect 6880 1204 6886 1216
rect 7742 1204 7748 1216
rect 6880 1176 7748 1204
rect 6880 1164 6886 1176
rect 7742 1164 7748 1176
rect 7800 1164 7806 1216
rect 552 1114 11408 1136
rect 552 1062 1755 1114
rect 1807 1062 1819 1114
rect 1871 1062 1883 1114
rect 1935 1062 1947 1114
rect 1999 1062 2011 1114
rect 2063 1062 4469 1114
rect 4521 1062 4533 1114
rect 4585 1062 4597 1114
rect 4649 1062 4661 1114
rect 4713 1062 4725 1114
rect 4777 1062 7183 1114
rect 7235 1062 7247 1114
rect 7299 1062 7311 1114
rect 7363 1062 7375 1114
rect 7427 1062 7439 1114
rect 7491 1062 9897 1114
rect 9949 1062 9961 1114
rect 10013 1062 10025 1114
rect 10077 1062 10089 1114
rect 10141 1062 10153 1114
rect 10205 1062 11408 1114
rect 552 1040 11408 1062
rect 3694 960 3700 1012
rect 3752 960 3758 1012
rect 7193 1003 7251 1009
rect 7193 969 7205 1003
rect 7239 1000 7251 1003
rect 7650 1000 7656 1012
rect 7239 972 7656 1000
rect 7239 969 7251 972
rect 7193 963 7251 969
rect 7650 960 7656 972
rect 7708 960 7714 1012
rect 8846 960 8852 1012
rect 8904 1000 8910 1012
rect 9677 1003 9735 1009
rect 9677 1000 9689 1003
rect 8904 972 9689 1000
rect 8904 960 8910 972
rect 9677 969 9689 972
rect 9723 969 9735 1003
rect 9677 963 9735 969
rect 6641 867 6699 873
rect 6641 833 6653 867
rect 6687 864 6699 867
rect 7377 867 7435 873
rect 7377 864 7389 867
rect 6687 836 7389 864
rect 6687 833 6699 836
rect 6641 827 6699 833
rect 7377 833 7389 836
rect 7423 833 7435 867
rect 7377 827 7435 833
rect 6914 756 6920 808
rect 6972 796 6978 808
rect 7285 799 7343 805
rect 7285 796 7297 799
rect 6972 768 7297 796
rect 6972 756 6978 768
rect 7285 765 7297 768
rect 7331 765 7343 799
rect 7285 759 7343 765
rect 7469 799 7527 805
rect 7469 765 7481 799
rect 7515 796 7527 799
rect 7742 796 7748 808
rect 7515 768 7748 796
rect 7515 765 7527 768
rect 7469 759 7527 765
rect 7742 756 7748 768
rect 7800 756 7806 808
rect 4985 731 5043 737
rect 4985 697 4997 731
rect 5031 728 5043 731
rect 7098 728 7104 740
rect 5031 700 7104 728
rect 5031 697 5043 700
rect 4985 691 5043 697
rect 7098 688 7104 700
rect 7156 728 7162 740
rect 8389 731 8447 737
rect 8389 728 8401 731
rect 7156 700 8401 728
rect 7156 688 7162 700
rect 8389 697 8401 700
rect 8435 697 8447 731
rect 8389 691 8447 697
rect 552 570 11568 592
rect 552 518 3112 570
rect 3164 518 3176 570
rect 3228 518 3240 570
rect 3292 518 3304 570
rect 3356 518 3368 570
rect 3420 518 5826 570
rect 5878 518 5890 570
rect 5942 518 5954 570
rect 6006 518 6018 570
rect 6070 518 6082 570
rect 6134 518 8540 570
rect 8592 518 8604 570
rect 8656 518 8668 570
rect 8720 518 8732 570
rect 8784 518 8796 570
rect 8848 518 11254 570
rect 11306 518 11318 570
rect 11370 518 11382 570
rect 11434 518 11446 570
rect 11498 518 11510 570
rect 11562 518 11568 570
rect 552 496 11568 518
<< via1 >>
rect 3112 11398 3164 11450
rect 3176 11398 3228 11450
rect 3240 11398 3292 11450
rect 3304 11398 3356 11450
rect 3368 11398 3420 11450
rect 5826 11398 5878 11450
rect 5890 11398 5942 11450
rect 5954 11398 6006 11450
rect 6018 11398 6070 11450
rect 6082 11398 6134 11450
rect 8540 11398 8592 11450
rect 8604 11398 8656 11450
rect 8668 11398 8720 11450
rect 8732 11398 8784 11450
rect 8796 11398 8848 11450
rect 11254 11398 11306 11450
rect 11318 11398 11370 11450
rect 11382 11398 11434 11450
rect 11446 11398 11498 11450
rect 11510 11398 11562 11450
rect 1755 10854 1807 10906
rect 1819 10854 1871 10906
rect 1883 10854 1935 10906
rect 1947 10854 1999 10906
rect 2011 10854 2063 10906
rect 4469 10854 4521 10906
rect 4533 10854 4585 10906
rect 4597 10854 4649 10906
rect 4661 10854 4713 10906
rect 4725 10854 4777 10906
rect 7183 10854 7235 10906
rect 7247 10854 7299 10906
rect 7311 10854 7363 10906
rect 7375 10854 7427 10906
rect 7439 10854 7491 10906
rect 9897 10854 9949 10906
rect 9961 10854 10013 10906
rect 10025 10854 10077 10906
rect 10089 10854 10141 10906
rect 10153 10854 10205 10906
rect 3112 10310 3164 10362
rect 3176 10310 3228 10362
rect 3240 10310 3292 10362
rect 3304 10310 3356 10362
rect 3368 10310 3420 10362
rect 5826 10310 5878 10362
rect 5890 10310 5942 10362
rect 5954 10310 6006 10362
rect 6018 10310 6070 10362
rect 6082 10310 6134 10362
rect 8540 10310 8592 10362
rect 8604 10310 8656 10362
rect 8668 10310 8720 10362
rect 8732 10310 8784 10362
rect 8796 10310 8848 10362
rect 11254 10310 11306 10362
rect 11318 10310 11370 10362
rect 11382 10310 11434 10362
rect 11446 10310 11498 10362
rect 11510 10310 11562 10362
rect 1755 9766 1807 9818
rect 1819 9766 1871 9818
rect 1883 9766 1935 9818
rect 1947 9766 1999 9818
rect 2011 9766 2063 9818
rect 4469 9766 4521 9818
rect 4533 9766 4585 9818
rect 4597 9766 4649 9818
rect 4661 9766 4713 9818
rect 4725 9766 4777 9818
rect 7183 9766 7235 9818
rect 7247 9766 7299 9818
rect 7311 9766 7363 9818
rect 7375 9766 7427 9818
rect 7439 9766 7491 9818
rect 9897 9766 9949 9818
rect 9961 9766 10013 9818
rect 10025 9766 10077 9818
rect 10089 9766 10141 9818
rect 10153 9766 10205 9818
rect 3112 9222 3164 9274
rect 3176 9222 3228 9274
rect 3240 9222 3292 9274
rect 3304 9222 3356 9274
rect 3368 9222 3420 9274
rect 5826 9222 5878 9274
rect 5890 9222 5942 9274
rect 5954 9222 6006 9274
rect 6018 9222 6070 9274
rect 6082 9222 6134 9274
rect 8540 9222 8592 9274
rect 8604 9222 8656 9274
rect 8668 9222 8720 9274
rect 8732 9222 8784 9274
rect 8796 9222 8848 9274
rect 11254 9222 11306 9274
rect 11318 9222 11370 9274
rect 11382 9222 11434 9274
rect 11446 9222 11498 9274
rect 11510 9222 11562 9274
rect 1755 8678 1807 8730
rect 1819 8678 1871 8730
rect 1883 8678 1935 8730
rect 1947 8678 1999 8730
rect 2011 8678 2063 8730
rect 4469 8678 4521 8730
rect 4533 8678 4585 8730
rect 4597 8678 4649 8730
rect 4661 8678 4713 8730
rect 4725 8678 4777 8730
rect 7183 8678 7235 8730
rect 7247 8678 7299 8730
rect 7311 8678 7363 8730
rect 7375 8678 7427 8730
rect 7439 8678 7491 8730
rect 9897 8678 9949 8730
rect 9961 8678 10013 8730
rect 10025 8678 10077 8730
rect 10089 8678 10141 8730
rect 10153 8678 10205 8730
rect 3112 8134 3164 8186
rect 3176 8134 3228 8186
rect 3240 8134 3292 8186
rect 3304 8134 3356 8186
rect 3368 8134 3420 8186
rect 5826 8134 5878 8186
rect 5890 8134 5942 8186
rect 5954 8134 6006 8186
rect 6018 8134 6070 8186
rect 6082 8134 6134 8186
rect 8540 8134 8592 8186
rect 8604 8134 8656 8186
rect 8668 8134 8720 8186
rect 8732 8134 8784 8186
rect 8796 8134 8848 8186
rect 11254 8134 11306 8186
rect 11318 8134 11370 8186
rect 11382 8134 11434 8186
rect 11446 8134 11498 8186
rect 11510 8134 11562 8186
rect 1755 7590 1807 7642
rect 1819 7590 1871 7642
rect 1883 7590 1935 7642
rect 1947 7590 1999 7642
rect 2011 7590 2063 7642
rect 4469 7590 4521 7642
rect 4533 7590 4585 7642
rect 4597 7590 4649 7642
rect 4661 7590 4713 7642
rect 4725 7590 4777 7642
rect 7183 7590 7235 7642
rect 7247 7590 7299 7642
rect 7311 7590 7363 7642
rect 7375 7590 7427 7642
rect 7439 7590 7491 7642
rect 9897 7590 9949 7642
rect 9961 7590 10013 7642
rect 10025 7590 10077 7642
rect 10089 7590 10141 7642
rect 10153 7590 10205 7642
rect 2780 7488 2832 7540
rect 5540 7488 5592 7540
rect 3112 7046 3164 7098
rect 3176 7046 3228 7098
rect 3240 7046 3292 7098
rect 3304 7046 3356 7098
rect 3368 7046 3420 7098
rect 5826 7046 5878 7098
rect 5890 7046 5942 7098
rect 5954 7046 6006 7098
rect 6018 7046 6070 7098
rect 6082 7046 6134 7098
rect 8540 7046 8592 7098
rect 8604 7046 8656 7098
rect 8668 7046 8720 7098
rect 8732 7046 8784 7098
rect 8796 7046 8848 7098
rect 11254 7046 11306 7098
rect 11318 7046 11370 7098
rect 11382 7046 11434 7098
rect 11446 7046 11498 7098
rect 11510 7046 11562 7098
rect 1755 6502 1807 6554
rect 1819 6502 1871 6554
rect 1883 6502 1935 6554
rect 1947 6502 1999 6554
rect 2011 6502 2063 6554
rect 4469 6502 4521 6554
rect 4533 6502 4585 6554
rect 4597 6502 4649 6554
rect 4661 6502 4713 6554
rect 4725 6502 4777 6554
rect 7183 6502 7235 6554
rect 7247 6502 7299 6554
rect 7311 6502 7363 6554
rect 7375 6502 7427 6554
rect 7439 6502 7491 6554
rect 9897 6502 9949 6554
rect 9961 6502 10013 6554
rect 10025 6502 10077 6554
rect 10089 6502 10141 6554
rect 10153 6502 10205 6554
rect 3112 5958 3164 6010
rect 3176 5958 3228 6010
rect 3240 5958 3292 6010
rect 3304 5958 3356 6010
rect 3368 5958 3420 6010
rect 5826 5958 5878 6010
rect 5890 5958 5942 6010
rect 5954 5958 6006 6010
rect 6018 5958 6070 6010
rect 6082 5958 6134 6010
rect 8540 5958 8592 6010
rect 8604 5958 8656 6010
rect 8668 5958 8720 6010
rect 8732 5958 8784 6010
rect 8796 5958 8848 6010
rect 11254 5958 11306 6010
rect 11318 5958 11370 6010
rect 11382 5958 11434 6010
rect 11446 5958 11498 6010
rect 11510 5958 11562 6010
rect 1755 5414 1807 5466
rect 1819 5414 1871 5466
rect 1883 5414 1935 5466
rect 1947 5414 1999 5466
rect 2011 5414 2063 5466
rect 4469 5414 4521 5466
rect 4533 5414 4585 5466
rect 4597 5414 4649 5466
rect 4661 5414 4713 5466
rect 4725 5414 4777 5466
rect 7183 5414 7235 5466
rect 7247 5414 7299 5466
rect 7311 5414 7363 5466
rect 7375 5414 7427 5466
rect 7439 5414 7491 5466
rect 9897 5414 9949 5466
rect 9961 5414 10013 5466
rect 10025 5414 10077 5466
rect 10089 5414 10141 5466
rect 10153 5414 10205 5466
rect 3112 4870 3164 4922
rect 3176 4870 3228 4922
rect 3240 4870 3292 4922
rect 3304 4870 3356 4922
rect 3368 4870 3420 4922
rect 5826 4870 5878 4922
rect 5890 4870 5942 4922
rect 5954 4870 6006 4922
rect 6018 4870 6070 4922
rect 6082 4870 6134 4922
rect 8540 4870 8592 4922
rect 8604 4870 8656 4922
rect 8668 4870 8720 4922
rect 8732 4870 8784 4922
rect 8796 4870 8848 4922
rect 11254 4870 11306 4922
rect 11318 4870 11370 4922
rect 11382 4870 11434 4922
rect 11446 4870 11498 4922
rect 11510 4870 11562 4922
rect 1755 4326 1807 4378
rect 1819 4326 1871 4378
rect 1883 4326 1935 4378
rect 1947 4326 1999 4378
rect 2011 4326 2063 4378
rect 4469 4326 4521 4378
rect 4533 4326 4585 4378
rect 4597 4326 4649 4378
rect 4661 4326 4713 4378
rect 4725 4326 4777 4378
rect 7183 4326 7235 4378
rect 7247 4326 7299 4378
rect 7311 4326 7363 4378
rect 7375 4326 7427 4378
rect 7439 4326 7491 4378
rect 9897 4326 9949 4378
rect 9961 4326 10013 4378
rect 10025 4326 10077 4378
rect 10089 4326 10141 4378
rect 10153 4326 10205 4378
rect 6828 4088 6880 4140
rect 11612 4088 11664 4140
rect 3112 3782 3164 3834
rect 3176 3782 3228 3834
rect 3240 3782 3292 3834
rect 3304 3782 3356 3834
rect 3368 3782 3420 3834
rect 5826 3782 5878 3834
rect 5890 3782 5942 3834
rect 5954 3782 6006 3834
rect 6018 3782 6070 3834
rect 6082 3782 6134 3834
rect 8540 3782 8592 3834
rect 8604 3782 8656 3834
rect 8668 3782 8720 3834
rect 8732 3782 8784 3834
rect 8796 3782 8848 3834
rect 11254 3782 11306 3834
rect 11318 3782 11370 3834
rect 11382 3782 11434 3834
rect 11446 3782 11498 3834
rect 11510 3782 11562 3834
rect 6828 3723 6880 3732
rect 6828 3689 6837 3723
rect 6837 3689 6871 3723
rect 6871 3689 6880 3723
rect 6828 3680 6880 3689
rect 6276 3612 6328 3664
rect 5724 3476 5776 3528
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 8944 3476 8996 3528
rect 11244 3476 11296 3528
rect 5632 3340 5684 3392
rect 6368 3340 6420 3392
rect 10600 3383 10652 3392
rect 10600 3349 10609 3383
rect 10609 3349 10643 3383
rect 10643 3349 10652 3383
rect 10600 3340 10652 3349
rect 1755 3238 1807 3290
rect 1819 3238 1871 3290
rect 1883 3238 1935 3290
rect 1947 3238 1999 3290
rect 2011 3238 2063 3290
rect 4469 3238 4521 3290
rect 4533 3238 4585 3290
rect 4597 3238 4649 3290
rect 4661 3238 4713 3290
rect 4725 3238 4777 3290
rect 7183 3238 7235 3290
rect 7247 3238 7299 3290
rect 7311 3238 7363 3290
rect 7375 3238 7427 3290
rect 7439 3238 7491 3290
rect 9897 3238 9949 3290
rect 9961 3238 10013 3290
rect 10025 3238 10077 3290
rect 10089 3238 10141 3290
rect 10153 3238 10205 3290
rect 8116 3136 8168 3188
rect 10600 3136 10652 3188
rect 4344 2975 4396 2984
rect 4344 2941 4353 2975
rect 4353 2941 4387 2975
rect 4387 2941 4396 2975
rect 4344 2932 4396 2941
rect 5540 2932 5592 2984
rect 6184 2932 6236 2984
rect 3700 2796 3752 2848
rect 5540 2796 5592 2848
rect 5724 2796 5776 2848
rect 6736 2796 6788 2848
rect 7104 2839 7156 2848
rect 7104 2805 7113 2839
rect 7113 2805 7147 2839
rect 7147 2805 7156 2839
rect 7104 2796 7156 2805
rect 8300 2796 8352 2848
rect 8392 2796 8444 2848
rect 3112 2694 3164 2746
rect 3176 2694 3228 2746
rect 3240 2694 3292 2746
rect 3304 2694 3356 2746
rect 3368 2694 3420 2746
rect 5826 2694 5878 2746
rect 5890 2694 5942 2746
rect 5954 2694 6006 2746
rect 6018 2694 6070 2746
rect 6082 2694 6134 2746
rect 8540 2694 8592 2746
rect 8604 2694 8656 2746
rect 8668 2694 8720 2746
rect 8732 2694 8784 2746
rect 8796 2694 8848 2746
rect 11254 2694 11306 2746
rect 11318 2694 11370 2746
rect 11382 2694 11434 2746
rect 11446 2694 11498 2746
rect 11510 2694 11562 2746
rect 5632 2592 5684 2644
rect 6736 2635 6788 2644
rect 6736 2601 6745 2635
rect 6745 2601 6779 2635
rect 6779 2601 6788 2635
rect 6736 2592 6788 2601
rect 4068 2499 4120 2508
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 7012 2524 7064 2576
rect 8392 2592 8444 2644
rect 8300 2524 8352 2576
rect 4896 2456 4948 2508
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 6184 2456 6236 2508
rect 6644 2499 6696 2508
rect 6644 2465 6653 2499
rect 6653 2465 6687 2499
rect 6687 2465 6696 2499
rect 6644 2456 6696 2465
rect 6276 2388 6328 2440
rect 4068 2252 4120 2304
rect 4160 2252 4212 2304
rect 4252 2295 4304 2304
rect 4252 2261 4261 2295
rect 4261 2261 4295 2295
rect 4295 2261 4304 2295
rect 4252 2252 4304 2261
rect 8944 2388 8996 2440
rect 5540 2252 5592 2304
rect 6368 2252 6420 2304
rect 6828 2252 6880 2304
rect 1755 2150 1807 2202
rect 1819 2150 1871 2202
rect 1883 2150 1935 2202
rect 1947 2150 1999 2202
rect 2011 2150 2063 2202
rect 4469 2150 4521 2202
rect 4533 2150 4585 2202
rect 4597 2150 4649 2202
rect 4661 2150 4713 2202
rect 4725 2150 4777 2202
rect 7183 2150 7235 2202
rect 7247 2150 7299 2202
rect 7311 2150 7363 2202
rect 7375 2150 7427 2202
rect 7439 2150 7491 2202
rect 9897 2150 9949 2202
rect 9961 2150 10013 2202
rect 10025 2150 10077 2202
rect 10089 2150 10141 2202
rect 10153 2150 10205 2202
rect 3700 1980 3752 2032
rect 4528 1955 4580 1964
rect 4528 1921 4537 1955
rect 4537 1921 4571 1955
rect 4571 1921 4580 1955
rect 4528 1912 4580 1921
rect 4068 1887 4120 1896
rect 4068 1853 4077 1887
rect 4077 1853 4111 1887
rect 4111 1853 4120 1887
rect 4068 1844 4120 1853
rect 4252 1844 4304 1896
rect 7012 2048 7064 2100
rect 4896 1912 4948 1964
rect 20 1776 72 1828
rect 4160 1751 4212 1760
rect 4160 1717 4169 1751
rect 4169 1717 4203 1751
rect 4203 1717 4212 1751
rect 4160 1708 4212 1717
rect 4988 1887 5040 1896
rect 4988 1853 4997 1887
rect 4997 1853 5031 1887
rect 5031 1853 5040 1887
rect 4988 1844 5040 1853
rect 6184 1708 6236 1760
rect 6920 1708 6972 1760
rect 3112 1606 3164 1658
rect 3176 1606 3228 1658
rect 3240 1606 3292 1658
rect 3304 1606 3356 1658
rect 3368 1606 3420 1658
rect 5826 1606 5878 1658
rect 5890 1606 5942 1658
rect 5954 1606 6006 1658
rect 6018 1606 6070 1658
rect 6082 1606 6134 1658
rect 8540 1606 8592 1658
rect 8604 1606 8656 1658
rect 8668 1606 8720 1658
rect 8732 1606 8784 1658
rect 8796 1606 8848 1658
rect 11254 1606 11306 1658
rect 11318 1606 11370 1658
rect 11382 1606 11434 1658
rect 11446 1606 11498 1658
rect 11510 1606 11562 1658
rect 3792 1504 3844 1556
rect 4988 1504 5040 1556
rect 6920 1436 6972 1488
rect 4160 1368 4212 1420
rect 5540 1343 5592 1352
rect 5540 1309 5549 1343
rect 5549 1309 5583 1343
rect 5583 1309 5592 1343
rect 5540 1300 5592 1309
rect 6184 1368 6236 1420
rect 7656 1343 7708 1352
rect 7656 1309 7665 1343
rect 7665 1309 7699 1343
rect 7699 1309 7708 1343
rect 7656 1300 7708 1309
rect 8852 1300 8904 1352
rect 6828 1164 6880 1216
rect 7748 1164 7800 1216
rect 1755 1062 1807 1114
rect 1819 1062 1871 1114
rect 1883 1062 1935 1114
rect 1947 1062 1999 1114
rect 2011 1062 2063 1114
rect 4469 1062 4521 1114
rect 4533 1062 4585 1114
rect 4597 1062 4649 1114
rect 4661 1062 4713 1114
rect 4725 1062 4777 1114
rect 7183 1062 7235 1114
rect 7247 1062 7299 1114
rect 7311 1062 7363 1114
rect 7375 1062 7427 1114
rect 7439 1062 7491 1114
rect 9897 1062 9949 1114
rect 9961 1062 10013 1114
rect 10025 1062 10077 1114
rect 10089 1062 10141 1114
rect 10153 1062 10205 1114
rect 3700 1003 3752 1012
rect 3700 969 3709 1003
rect 3709 969 3743 1003
rect 3743 969 3752 1003
rect 3700 960 3752 969
rect 7656 960 7708 1012
rect 8852 960 8904 1012
rect 6920 756 6972 808
rect 7748 756 7800 808
rect 7104 688 7156 740
rect 3112 518 3164 570
rect 3176 518 3228 570
rect 3240 518 3292 570
rect 3304 518 3356 570
rect 3368 518 3420 570
rect 5826 518 5878 570
rect 5890 518 5942 570
rect 5954 518 6006 570
rect 6018 518 6070 570
rect 6082 518 6134 570
rect 8540 518 8592 570
rect 8604 518 8656 570
rect 8668 518 8720 570
rect 8732 518 8784 570
rect 8796 518 8848 570
rect 11254 518 11306 570
rect 11318 518 11370 570
rect 11382 518 11434 570
rect 11446 518 11498 570
rect 11510 518 11562 570
<< metal2 >>
rect 3882 11600 3938 12000
rect 11610 11600 11666 12000
rect 3112 11452 3420 11461
rect 3112 11450 3118 11452
rect 3174 11450 3198 11452
rect 3254 11450 3278 11452
rect 3334 11450 3358 11452
rect 3414 11450 3420 11452
rect 3174 11398 3176 11450
rect 3356 11398 3358 11450
rect 3112 11396 3118 11398
rect 3174 11396 3198 11398
rect 3254 11396 3278 11398
rect 3334 11396 3358 11398
rect 3414 11396 3420 11398
rect 3112 11387 3420 11396
rect 1755 10908 2063 10917
rect 1755 10906 1761 10908
rect 1817 10906 1841 10908
rect 1897 10906 1921 10908
rect 1977 10906 2001 10908
rect 2057 10906 2063 10908
rect 1817 10854 1819 10906
rect 1999 10854 2001 10906
rect 1755 10852 1761 10854
rect 1817 10852 1841 10854
rect 1897 10852 1921 10854
rect 1977 10852 2001 10854
rect 2057 10852 2063 10854
rect 1755 10843 2063 10852
rect 3112 10364 3420 10373
rect 3112 10362 3118 10364
rect 3174 10362 3198 10364
rect 3254 10362 3278 10364
rect 3334 10362 3358 10364
rect 3414 10362 3420 10364
rect 3174 10310 3176 10362
rect 3356 10310 3358 10362
rect 3112 10308 3118 10310
rect 3174 10308 3198 10310
rect 3254 10308 3278 10310
rect 3334 10308 3358 10310
rect 3414 10308 3420 10310
rect 3112 10299 3420 10308
rect 1755 9820 2063 9829
rect 1755 9818 1761 9820
rect 1817 9818 1841 9820
rect 1897 9818 1921 9820
rect 1977 9818 2001 9820
rect 2057 9818 2063 9820
rect 1817 9766 1819 9818
rect 1999 9766 2001 9818
rect 1755 9764 1761 9766
rect 1817 9764 1841 9766
rect 1897 9764 1921 9766
rect 1977 9764 2001 9766
rect 2057 9764 2063 9766
rect 1755 9755 2063 9764
rect 3112 9276 3420 9285
rect 3112 9274 3118 9276
rect 3174 9274 3198 9276
rect 3254 9274 3278 9276
rect 3334 9274 3358 9276
rect 3414 9274 3420 9276
rect 3174 9222 3176 9274
rect 3356 9222 3358 9274
rect 3112 9220 3118 9222
rect 3174 9220 3198 9222
rect 3254 9220 3278 9222
rect 3334 9220 3358 9222
rect 3414 9220 3420 9222
rect 3112 9211 3420 9220
rect 1755 8732 2063 8741
rect 1755 8730 1761 8732
rect 1817 8730 1841 8732
rect 1897 8730 1921 8732
rect 1977 8730 2001 8732
rect 2057 8730 2063 8732
rect 1817 8678 1819 8730
rect 1999 8678 2001 8730
rect 1755 8676 1761 8678
rect 1817 8676 1841 8678
rect 1897 8676 1921 8678
rect 1977 8676 2001 8678
rect 2057 8676 2063 8678
rect 1755 8667 2063 8676
rect 2778 8256 2834 8265
rect 2778 8191 2834 8200
rect 1755 7644 2063 7653
rect 1755 7642 1761 7644
rect 1817 7642 1841 7644
rect 1897 7642 1921 7644
rect 1977 7642 2001 7644
rect 2057 7642 2063 7644
rect 1817 7590 1819 7642
rect 1999 7590 2001 7642
rect 1755 7588 1761 7590
rect 1817 7588 1841 7590
rect 1897 7588 1921 7590
rect 1977 7588 2001 7590
rect 2057 7588 2063 7590
rect 1755 7579 2063 7588
rect 2792 7546 2820 8191
rect 3112 8188 3420 8197
rect 3112 8186 3118 8188
rect 3174 8186 3198 8188
rect 3254 8186 3278 8188
rect 3334 8186 3358 8188
rect 3414 8186 3420 8188
rect 3174 8134 3176 8186
rect 3356 8134 3358 8186
rect 3112 8132 3118 8134
rect 3174 8132 3198 8134
rect 3254 8132 3278 8134
rect 3334 8132 3358 8134
rect 3414 8132 3420 8134
rect 3112 8123 3420 8132
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 3112 7100 3420 7109
rect 3112 7098 3118 7100
rect 3174 7098 3198 7100
rect 3254 7098 3278 7100
rect 3334 7098 3358 7100
rect 3414 7098 3420 7100
rect 3174 7046 3176 7098
rect 3356 7046 3358 7098
rect 3112 7044 3118 7046
rect 3174 7044 3198 7046
rect 3254 7044 3278 7046
rect 3334 7044 3358 7046
rect 3414 7044 3420 7046
rect 3112 7035 3420 7044
rect 3896 6914 3924 11600
rect 5826 11452 6134 11461
rect 5826 11450 5832 11452
rect 5888 11450 5912 11452
rect 5968 11450 5992 11452
rect 6048 11450 6072 11452
rect 6128 11450 6134 11452
rect 5888 11398 5890 11450
rect 6070 11398 6072 11450
rect 5826 11396 5832 11398
rect 5888 11396 5912 11398
rect 5968 11396 5992 11398
rect 6048 11396 6072 11398
rect 6128 11396 6134 11398
rect 5826 11387 6134 11396
rect 8540 11452 8848 11461
rect 8540 11450 8546 11452
rect 8602 11450 8626 11452
rect 8682 11450 8706 11452
rect 8762 11450 8786 11452
rect 8842 11450 8848 11452
rect 8602 11398 8604 11450
rect 8784 11398 8786 11450
rect 8540 11396 8546 11398
rect 8602 11396 8626 11398
rect 8682 11396 8706 11398
rect 8762 11396 8786 11398
rect 8842 11396 8848 11398
rect 8540 11387 8848 11396
rect 11254 11452 11562 11461
rect 11254 11450 11260 11452
rect 11316 11450 11340 11452
rect 11396 11450 11420 11452
rect 11476 11450 11500 11452
rect 11556 11450 11562 11452
rect 11316 11398 11318 11450
rect 11498 11398 11500 11450
rect 11254 11396 11260 11398
rect 11316 11396 11340 11398
rect 11396 11396 11420 11398
rect 11476 11396 11500 11398
rect 11556 11396 11562 11398
rect 11254 11387 11562 11396
rect 4469 10908 4777 10917
rect 4469 10906 4475 10908
rect 4531 10906 4555 10908
rect 4611 10906 4635 10908
rect 4691 10906 4715 10908
rect 4771 10906 4777 10908
rect 4531 10854 4533 10906
rect 4713 10854 4715 10906
rect 4469 10852 4475 10854
rect 4531 10852 4555 10854
rect 4611 10852 4635 10854
rect 4691 10852 4715 10854
rect 4771 10852 4777 10854
rect 4469 10843 4777 10852
rect 7183 10908 7491 10917
rect 7183 10906 7189 10908
rect 7245 10906 7269 10908
rect 7325 10906 7349 10908
rect 7405 10906 7429 10908
rect 7485 10906 7491 10908
rect 7245 10854 7247 10906
rect 7427 10854 7429 10906
rect 7183 10852 7189 10854
rect 7245 10852 7269 10854
rect 7325 10852 7349 10854
rect 7405 10852 7429 10854
rect 7485 10852 7491 10854
rect 7183 10843 7491 10852
rect 9897 10908 10205 10917
rect 9897 10906 9903 10908
rect 9959 10906 9983 10908
rect 10039 10906 10063 10908
rect 10119 10906 10143 10908
rect 10199 10906 10205 10908
rect 9959 10854 9961 10906
rect 10141 10854 10143 10906
rect 9897 10852 9903 10854
rect 9959 10852 9983 10854
rect 10039 10852 10063 10854
rect 10119 10852 10143 10854
rect 10199 10852 10205 10854
rect 9897 10843 10205 10852
rect 5826 10364 6134 10373
rect 5826 10362 5832 10364
rect 5888 10362 5912 10364
rect 5968 10362 5992 10364
rect 6048 10362 6072 10364
rect 6128 10362 6134 10364
rect 5888 10310 5890 10362
rect 6070 10310 6072 10362
rect 5826 10308 5832 10310
rect 5888 10308 5912 10310
rect 5968 10308 5992 10310
rect 6048 10308 6072 10310
rect 6128 10308 6134 10310
rect 5826 10299 6134 10308
rect 8540 10364 8848 10373
rect 8540 10362 8546 10364
rect 8602 10362 8626 10364
rect 8682 10362 8706 10364
rect 8762 10362 8786 10364
rect 8842 10362 8848 10364
rect 8602 10310 8604 10362
rect 8784 10310 8786 10362
rect 8540 10308 8546 10310
rect 8602 10308 8626 10310
rect 8682 10308 8706 10310
rect 8762 10308 8786 10310
rect 8842 10308 8848 10310
rect 8540 10299 8848 10308
rect 11254 10364 11562 10373
rect 11254 10362 11260 10364
rect 11316 10362 11340 10364
rect 11396 10362 11420 10364
rect 11476 10362 11500 10364
rect 11556 10362 11562 10364
rect 11316 10310 11318 10362
rect 11498 10310 11500 10362
rect 11254 10308 11260 10310
rect 11316 10308 11340 10310
rect 11396 10308 11420 10310
rect 11476 10308 11500 10310
rect 11556 10308 11562 10310
rect 11254 10299 11562 10308
rect 4469 9820 4777 9829
rect 4469 9818 4475 9820
rect 4531 9818 4555 9820
rect 4611 9818 4635 9820
rect 4691 9818 4715 9820
rect 4771 9818 4777 9820
rect 4531 9766 4533 9818
rect 4713 9766 4715 9818
rect 4469 9764 4475 9766
rect 4531 9764 4555 9766
rect 4611 9764 4635 9766
rect 4691 9764 4715 9766
rect 4771 9764 4777 9766
rect 4469 9755 4777 9764
rect 7183 9820 7491 9829
rect 7183 9818 7189 9820
rect 7245 9818 7269 9820
rect 7325 9818 7349 9820
rect 7405 9818 7429 9820
rect 7485 9818 7491 9820
rect 7245 9766 7247 9818
rect 7427 9766 7429 9818
rect 7183 9764 7189 9766
rect 7245 9764 7269 9766
rect 7325 9764 7349 9766
rect 7405 9764 7429 9766
rect 7485 9764 7491 9766
rect 7183 9755 7491 9764
rect 9897 9820 10205 9829
rect 9897 9818 9903 9820
rect 9959 9818 9983 9820
rect 10039 9818 10063 9820
rect 10119 9818 10143 9820
rect 10199 9818 10205 9820
rect 9959 9766 9961 9818
rect 10141 9766 10143 9818
rect 9897 9764 9903 9766
rect 9959 9764 9983 9766
rect 10039 9764 10063 9766
rect 10119 9764 10143 9766
rect 10199 9764 10205 9766
rect 9897 9755 10205 9764
rect 5826 9276 6134 9285
rect 5826 9274 5832 9276
rect 5888 9274 5912 9276
rect 5968 9274 5992 9276
rect 6048 9274 6072 9276
rect 6128 9274 6134 9276
rect 5888 9222 5890 9274
rect 6070 9222 6072 9274
rect 5826 9220 5832 9222
rect 5888 9220 5912 9222
rect 5968 9220 5992 9222
rect 6048 9220 6072 9222
rect 6128 9220 6134 9222
rect 5826 9211 6134 9220
rect 8540 9276 8848 9285
rect 8540 9274 8546 9276
rect 8602 9274 8626 9276
rect 8682 9274 8706 9276
rect 8762 9274 8786 9276
rect 8842 9274 8848 9276
rect 8602 9222 8604 9274
rect 8784 9222 8786 9274
rect 8540 9220 8546 9222
rect 8602 9220 8626 9222
rect 8682 9220 8706 9222
rect 8762 9220 8786 9222
rect 8842 9220 8848 9222
rect 8540 9211 8848 9220
rect 11254 9276 11562 9285
rect 11254 9274 11260 9276
rect 11316 9274 11340 9276
rect 11396 9274 11420 9276
rect 11476 9274 11500 9276
rect 11556 9274 11562 9276
rect 11316 9222 11318 9274
rect 11498 9222 11500 9274
rect 11254 9220 11260 9222
rect 11316 9220 11340 9222
rect 11396 9220 11420 9222
rect 11476 9220 11500 9222
rect 11556 9220 11562 9222
rect 11254 9211 11562 9220
rect 4469 8732 4777 8741
rect 4469 8730 4475 8732
rect 4531 8730 4555 8732
rect 4611 8730 4635 8732
rect 4691 8730 4715 8732
rect 4771 8730 4777 8732
rect 4531 8678 4533 8730
rect 4713 8678 4715 8730
rect 4469 8676 4475 8678
rect 4531 8676 4555 8678
rect 4611 8676 4635 8678
rect 4691 8676 4715 8678
rect 4771 8676 4777 8678
rect 4469 8667 4777 8676
rect 7183 8732 7491 8741
rect 7183 8730 7189 8732
rect 7245 8730 7269 8732
rect 7325 8730 7349 8732
rect 7405 8730 7429 8732
rect 7485 8730 7491 8732
rect 7245 8678 7247 8730
rect 7427 8678 7429 8730
rect 7183 8676 7189 8678
rect 7245 8676 7269 8678
rect 7325 8676 7349 8678
rect 7405 8676 7429 8678
rect 7485 8676 7491 8678
rect 7183 8667 7491 8676
rect 9897 8732 10205 8741
rect 9897 8730 9903 8732
rect 9959 8730 9983 8732
rect 10039 8730 10063 8732
rect 10119 8730 10143 8732
rect 10199 8730 10205 8732
rect 9959 8678 9961 8730
rect 10141 8678 10143 8730
rect 9897 8676 9903 8678
rect 9959 8676 9983 8678
rect 10039 8676 10063 8678
rect 10119 8676 10143 8678
rect 10199 8676 10205 8678
rect 9897 8667 10205 8676
rect 5826 8188 6134 8197
rect 5826 8186 5832 8188
rect 5888 8186 5912 8188
rect 5968 8186 5992 8188
rect 6048 8186 6072 8188
rect 6128 8186 6134 8188
rect 5888 8134 5890 8186
rect 6070 8134 6072 8186
rect 5826 8132 5832 8134
rect 5888 8132 5912 8134
rect 5968 8132 5992 8134
rect 6048 8132 6072 8134
rect 6128 8132 6134 8134
rect 5826 8123 6134 8132
rect 8540 8188 8848 8197
rect 8540 8186 8546 8188
rect 8602 8186 8626 8188
rect 8682 8186 8706 8188
rect 8762 8186 8786 8188
rect 8842 8186 8848 8188
rect 8602 8134 8604 8186
rect 8784 8134 8786 8186
rect 8540 8132 8546 8134
rect 8602 8132 8626 8134
rect 8682 8132 8706 8134
rect 8762 8132 8786 8134
rect 8842 8132 8848 8134
rect 8540 8123 8848 8132
rect 11254 8188 11562 8197
rect 11254 8186 11260 8188
rect 11316 8186 11340 8188
rect 11396 8186 11420 8188
rect 11476 8186 11500 8188
rect 11556 8186 11562 8188
rect 11316 8134 11318 8186
rect 11498 8134 11500 8186
rect 11254 8132 11260 8134
rect 11316 8132 11340 8134
rect 11396 8132 11420 8134
rect 11476 8132 11500 8134
rect 11556 8132 11562 8134
rect 11254 8123 11562 8132
rect 4469 7644 4777 7653
rect 4469 7642 4475 7644
rect 4531 7642 4555 7644
rect 4611 7642 4635 7644
rect 4691 7642 4715 7644
rect 4771 7642 4777 7644
rect 4531 7590 4533 7642
rect 4713 7590 4715 7642
rect 4469 7588 4475 7590
rect 4531 7588 4555 7590
rect 4611 7588 4635 7590
rect 4691 7588 4715 7590
rect 4771 7588 4777 7590
rect 4469 7579 4777 7588
rect 7183 7644 7491 7653
rect 7183 7642 7189 7644
rect 7245 7642 7269 7644
rect 7325 7642 7349 7644
rect 7405 7642 7429 7644
rect 7485 7642 7491 7644
rect 7245 7590 7247 7642
rect 7427 7590 7429 7642
rect 7183 7588 7189 7590
rect 7245 7588 7269 7590
rect 7325 7588 7349 7590
rect 7405 7588 7429 7590
rect 7485 7588 7491 7590
rect 7183 7579 7491 7588
rect 9897 7644 10205 7653
rect 9897 7642 9903 7644
rect 9959 7642 9983 7644
rect 10039 7642 10063 7644
rect 10119 7642 10143 7644
rect 10199 7642 10205 7644
rect 9959 7590 9961 7642
rect 10141 7590 10143 7642
rect 9897 7588 9903 7590
rect 9959 7588 9983 7590
rect 10039 7588 10063 7590
rect 10119 7588 10143 7590
rect 10199 7588 10205 7590
rect 9897 7579 10205 7588
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 3896 6886 4016 6914
rect 1755 6556 2063 6565
rect 1755 6554 1761 6556
rect 1817 6554 1841 6556
rect 1897 6554 1921 6556
rect 1977 6554 2001 6556
rect 2057 6554 2063 6556
rect 1817 6502 1819 6554
rect 1999 6502 2001 6554
rect 1755 6500 1761 6502
rect 1817 6500 1841 6502
rect 1897 6500 1921 6502
rect 1977 6500 2001 6502
rect 2057 6500 2063 6502
rect 1755 6491 2063 6500
rect 3112 6012 3420 6021
rect 3112 6010 3118 6012
rect 3174 6010 3198 6012
rect 3254 6010 3278 6012
rect 3334 6010 3358 6012
rect 3414 6010 3420 6012
rect 3174 5958 3176 6010
rect 3356 5958 3358 6010
rect 3112 5956 3118 5958
rect 3174 5956 3198 5958
rect 3254 5956 3278 5958
rect 3334 5956 3358 5958
rect 3414 5956 3420 5958
rect 3112 5947 3420 5956
rect 1755 5468 2063 5477
rect 1755 5466 1761 5468
rect 1817 5466 1841 5468
rect 1897 5466 1921 5468
rect 1977 5466 2001 5468
rect 2057 5466 2063 5468
rect 1817 5414 1819 5466
rect 1999 5414 2001 5466
rect 1755 5412 1761 5414
rect 1817 5412 1841 5414
rect 1897 5412 1921 5414
rect 1977 5412 2001 5414
rect 2057 5412 2063 5414
rect 1755 5403 2063 5412
rect 3112 4924 3420 4933
rect 3112 4922 3118 4924
rect 3174 4922 3198 4924
rect 3254 4922 3278 4924
rect 3334 4922 3358 4924
rect 3414 4922 3420 4924
rect 3174 4870 3176 4922
rect 3356 4870 3358 4922
rect 3112 4868 3118 4870
rect 3174 4868 3198 4870
rect 3254 4868 3278 4870
rect 3334 4868 3358 4870
rect 3414 4868 3420 4870
rect 3112 4859 3420 4868
rect 1755 4380 2063 4389
rect 1755 4378 1761 4380
rect 1817 4378 1841 4380
rect 1897 4378 1921 4380
rect 1977 4378 2001 4380
rect 2057 4378 2063 4380
rect 1817 4326 1819 4378
rect 1999 4326 2001 4378
rect 1755 4324 1761 4326
rect 1817 4324 1841 4326
rect 1897 4324 1921 4326
rect 1977 4324 2001 4326
rect 2057 4324 2063 4326
rect 1755 4315 2063 4324
rect 3112 3836 3420 3845
rect 3112 3834 3118 3836
rect 3174 3834 3198 3836
rect 3254 3834 3278 3836
rect 3334 3834 3358 3836
rect 3414 3834 3420 3836
rect 3174 3782 3176 3834
rect 3356 3782 3358 3834
rect 3112 3780 3118 3782
rect 3174 3780 3198 3782
rect 3254 3780 3278 3782
rect 3334 3780 3358 3782
rect 3414 3780 3420 3782
rect 3112 3771 3420 3780
rect 1755 3292 2063 3301
rect 1755 3290 1761 3292
rect 1817 3290 1841 3292
rect 1897 3290 1921 3292
rect 1977 3290 2001 3292
rect 2057 3290 2063 3292
rect 1817 3238 1819 3290
rect 1999 3238 2001 3290
rect 1755 3236 1761 3238
rect 1817 3236 1841 3238
rect 1897 3236 1921 3238
rect 1977 3236 2001 3238
rect 2057 3236 2063 3238
rect 1755 3227 2063 3236
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3112 2748 3420 2757
rect 3112 2746 3118 2748
rect 3174 2746 3198 2748
rect 3254 2746 3278 2748
rect 3334 2746 3358 2748
rect 3414 2746 3420 2748
rect 3174 2694 3176 2746
rect 3356 2694 3358 2746
rect 3112 2692 3118 2694
rect 3174 2692 3198 2694
rect 3254 2692 3278 2694
rect 3334 2692 3358 2694
rect 3414 2692 3420 2694
rect 3112 2683 3420 2692
rect 1755 2204 2063 2213
rect 1755 2202 1761 2204
rect 1817 2202 1841 2204
rect 1897 2202 1921 2204
rect 1977 2202 2001 2204
rect 2057 2202 2063 2204
rect 1817 2150 1819 2202
rect 1999 2150 2001 2202
rect 1755 2148 1761 2150
rect 1817 2148 1841 2150
rect 1897 2148 1921 2150
rect 1977 2148 2001 2150
rect 2057 2148 2063 2150
rect 1755 2139 2063 2148
rect 3712 2038 3740 2790
rect 3988 2774 4016 6886
rect 4469 6556 4777 6565
rect 4469 6554 4475 6556
rect 4531 6554 4555 6556
rect 4611 6554 4635 6556
rect 4691 6554 4715 6556
rect 4771 6554 4777 6556
rect 4531 6502 4533 6554
rect 4713 6502 4715 6554
rect 4469 6500 4475 6502
rect 4531 6500 4555 6502
rect 4611 6500 4635 6502
rect 4691 6500 4715 6502
rect 4771 6500 4777 6502
rect 4469 6491 4777 6500
rect 4469 5468 4777 5477
rect 4469 5466 4475 5468
rect 4531 5466 4555 5468
rect 4611 5466 4635 5468
rect 4691 5466 4715 5468
rect 4771 5466 4777 5468
rect 4531 5414 4533 5466
rect 4713 5414 4715 5466
rect 4469 5412 4475 5414
rect 4531 5412 4555 5414
rect 4611 5412 4635 5414
rect 4691 5412 4715 5414
rect 4771 5412 4777 5414
rect 4469 5403 4777 5412
rect 4469 4380 4777 4389
rect 4469 4378 4475 4380
rect 4531 4378 4555 4380
rect 4611 4378 4635 4380
rect 4691 4378 4715 4380
rect 4771 4378 4777 4380
rect 4531 4326 4533 4378
rect 4713 4326 4715 4378
rect 4469 4324 4475 4326
rect 4531 4324 4555 4326
rect 4611 4324 4635 4326
rect 4691 4324 4715 4326
rect 4771 4324 4777 4326
rect 4469 4315 4777 4324
rect 4469 3292 4777 3301
rect 4469 3290 4475 3292
rect 4531 3290 4555 3292
rect 4611 3290 4635 3292
rect 4691 3290 4715 3292
rect 4771 3290 4777 3292
rect 4531 3238 4533 3290
rect 4713 3238 4715 3290
rect 4469 3236 4475 3238
rect 4531 3236 4555 3238
rect 4611 3236 4635 3238
rect 4691 3236 4715 3238
rect 4771 3236 4777 3238
rect 4469 3227 4777 3236
rect 5552 2990 5580 7482
rect 5826 7100 6134 7109
rect 5826 7098 5832 7100
rect 5888 7098 5912 7100
rect 5968 7098 5992 7100
rect 6048 7098 6072 7100
rect 6128 7098 6134 7100
rect 5888 7046 5890 7098
rect 6070 7046 6072 7098
rect 5826 7044 5832 7046
rect 5888 7044 5912 7046
rect 5968 7044 5992 7046
rect 6048 7044 6072 7046
rect 6128 7044 6134 7046
rect 5826 7035 6134 7044
rect 8540 7100 8848 7109
rect 8540 7098 8546 7100
rect 8602 7098 8626 7100
rect 8682 7098 8706 7100
rect 8762 7098 8786 7100
rect 8842 7098 8848 7100
rect 8602 7046 8604 7098
rect 8784 7046 8786 7098
rect 8540 7044 8546 7046
rect 8602 7044 8626 7046
rect 8682 7044 8706 7046
rect 8762 7044 8786 7046
rect 8842 7044 8848 7046
rect 8540 7035 8848 7044
rect 11254 7100 11562 7109
rect 11254 7098 11260 7100
rect 11316 7098 11340 7100
rect 11396 7098 11420 7100
rect 11476 7098 11500 7100
rect 11556 7098 11562 7100
rect 11316 7046 11318 7098
rect 11498 7046 11500 7098
rect 11254 7044 11260 7046
rect 11316 7044 11340 7046
rect 11396 7044 11420 7046
rect 11476 7044 11500 7046
rect 11556 7044 11562 7046
rect 11254 7035 11562 7044
rect 7183 6556 7491 6565
rect 7183 6554 7189 6556
rect 7245 6554 7269 6556
rect 7325 6554 7349 6556
rect 7405 6554 7429 6556
rect 7485 6554 7491 6556
rect 7245 6502 7247 6554
rect 7427 6502 7429 6554
rect 7183 6500 7189 6502
rect 7245 6500 7269 6502
rect 7325 6500 7349 6502
rect 7405 6500 7429 6502
rect 7485 6500 7491 6502
rect 7183 6491 7491 6500
rect 9897 6556 10205 6565
rect 9897 6554 9903 6556
rect 9959 6554 9983 6556
rect 10039 6554 10063 6556
rect 10119 6554 10143 6556
rect 10199 6554 10205 6556
rect 9959 6502 9961 6554
rect 10141 6502 10143 6554
rect 9897 6500 9903 6502
rect 9959 6500 9983 6502
rect 10039 6500 10063 6502
rect 10119 6500 10143 6502
rect 10199 6500 10205 6502
rect 9897 6491 10205 6500
rect 5826 6012 6134 6021
rect 5826 6010 5832 6012
rect 5888 6010 5912 6012
rect 5968 6010 5992 6012
rect 6048 6010 6072 6012
rect 6128 6010 6134 6012
rect 5888 5958 5890 6010
rect 6070 5958 6072 6010
rect 5826 5956 5832 5958
rect 5888 5956 5912 5958
rect 5968 5956 5992 5958
rect 6048 5956 6072 5958
rect 6128 5956 6134 5958
rect 5826 5947 6134 5956
rect 8540 6012 8848 6021
rect 8540 6010 8546 6012
rect 8602 6010 8626 6012
rect 8682 6010 8706 6012
rect 8762 6010 8786 6012
rect 8842 6010 8848 6012
rect 8602 5958 8604 6010
rect 8784 5958 8786 6010
rect 8540 5956 8546 5958
rect 8602 5956 8626 5958
rect 8682 5956 8706 5958
rect 8762 5956 8786 5958
rect 8842 5956 8848 5958
rect 8540 5947 8848 5956
rect 11254 6012 11562 6021
rect 11254 6010 11260 6012
rect 11316 6010 11340 6012
rect 11396 6010 11420 6012
rect 11476 6010 11500 6012
rect 11556 6010 11562 6012
rect 11316 5958 11318 6010
rect 11498 5958 11500 6010
rect 11254 5956 11260 5958
rect 11316 5956 11340 5958
rect 11396 5956 11420 5958
rect 11476 5956 11500 5958
rect 11556 5956 11562 5958
rect 11254 5947 11562 5956
rect 7183 5468 7491 5477
rect 7183 5466 7189 5468
rect 7245 5466 7269 5468
rect 7325 5466 7349 5468
rect 7405 5466 7429 5468
rect 7485 5466 7491 5468
rect 7245 5414 7247 5466
rect 7427 5414 7429 5466
rect 7183 5412 7189 5414
rect 7245 5412 7269 5414
rect 7325 5412 7349 5414
rect 7405 5412 7429 5414
rect 7485 5412 7491 5414
rect 7183 5403 7491 5412
rect 9897 5468 10205 5477
rect 9897 5466 9903 5468
rect 9959 5466 9983 5468
rect 10039 5466 10063 5468
rect 10119 5466 10143 5468
rect 10199 5466 10205 5468
rect 9959 5414 9961 5466
rect 10141 5414 10143 5466
rect 9897 5412 9903 5414
rect 9959 5412 9983 5414
rect 10039 5412 10063 5414
rect 10119 5412 10143 5414
rect 10199 5412 10205 5414
rect 9897 5403 10205 5412
rect 5826 4924 6134 4933
rect 5826 4922 5832 4924
rect 5888 4922 5912 4924
rect 5968 4922 5992 4924
rect 6048 4922 6072 4924
rect 6128 4922 6134 4924
rect 5888 4870 5890 4922
rect 6070 4870 6072 4922
rect 5826 4868 5832 4870
rect 5888 4868 5912 4870
rect 5968 4868 5992 4870
rect 6048 4868 6072 4870
rect 6128 4868 6134 4870
rect 5826 4859 6134 4868
rect 8540 4924 8848 4933
rect 8540 4922 8546 4924
rect 8602 4922 8626 4924
rect 8682 4922 8706 4924
rect 8762 4922 8786 4924
rect 8842 4922 8848 4924
rect 8602 4870 8604 4922
rect 8784 4870 8786 4922
rect 8540 4868 8546 4870
rect 8602 4868 8626 4870
rect 8682 4868 8706 4870
rect 8762 4868 8786 4870
rect 8842 4868 8848 4870
rect 8540 4859 8848 4868
rect 11254 4924 11562 4933
rect 11254 4922 11260 4924
rect 11316 4922 11340 4924
rect 11396 4922 11420 4924
rect 11476 4922 11500 4924
rect 11556 4922 11562 4924
rect 11316 4870 11318 4922
rect 11498 4870 11500 4922
rect 11254 4868 11260 4870
rect 11316 4868 11340 4870
rect 11396 4868 11420 4870
rect 11476 4868 11500 4870
rect 11556 4868 11562 4870
rect 11254 4859 11562 4868
rect 7183 4380 7491 4389
rect 7183 4378 7189 4380
rect 7245 4378 7269 4380
rect 7325 4378 7349 4380
rect 7405 4378 7429 4380
rect 7485 4378 7491 4380
rect 7245 4326 7247 4378
rect 7427 4326 7429 4378
rect 7183 4324 7189 4326
rect 7245 4324 7269 4326
rect 7325 4324 7349 4326
rect 7405 4324 7429 4326
rect 7485 4324 7491 4326
rect 7183 4315 7491 4324
rect 9897 4380 10205 4389
rect 9897 4378 9903 4380
rect 9959 4378 9983 4380
rect 10039 4378 10063 4380
rect 10119 4378 10143 4380
rect 10199 4378 10205 4380
rect 9959 4326 9961 4378
rect 10141 4326 10143 4378
rect 9897 4324 9903 4326
rect 9959 4324 9983 4326
rect 10039 4324 10063 4326
rect 10119 4324 10143 4326
rect 10199 4324 10205 4326
rect 9897 4315 10205 4324
rect 11624 4146 11652 11600
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 5826 3836 6134 3845
rect 5826 3834 5832 3836
rect 5888 3834 5912 3836
rect 5968 3834 5992 3836
rect 6048 3834 6072 3836
rect 6128 3834 6134 3836
rect 5888 3782 5890 3834
rect 6070 3782 6072 3834
rect 5826 3780 5832 3782
rect 5888 3780 5912 3782
rect 5968 3780 5992 3782
rect 6048 3780 6072 3782
rect 6128 3780 6134 3782
rect 5826 3771 6134 3780
rect 6840 3738 6868 4082
rect 8540 3836 8848 3845
rect 8540 3834 8546 3836
rect 8602 3834 8626 3836
rect 8682 3834 8706 3836
rect 8762 3834 8786 3836
rect 8842 3834 8848 3836
rect 8602 3782 8604 3834
rect 8784 3782 8786 3834
rect 8540 3780 8546 3782
rect 8602 3780 8626 3782
rect 8682 3780 8706 3782
rect 8762 3780 8786 3782
rect 8842 3780 8848 3782
rect 8540 3771 8848 3780
rect 11254 3836 11562 3845
rect 11254 3834 11260 3836
rect 11316 3834 11340 3836
rect 11396 3834 11420 3836
rect 11476 3834 11500 3836
rect 11556 3834 11562 3836
rect 11316 3782 11318 3834
rect 11498 3782 11500 3834
rect 11254 3780 11260 3782
rect 11316 3780 11340 3782
rect 11396 3780 11420 3782
rect 11476 3780 11500 3782
rect 11556 3780 11562 3782
rect 11254 3771 11562 3780
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6276 3664 6328 3670
rect 6276 3606 6328 3612
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 3988 2746 4108 2774
rect 4080 2553 4108 2746
rect 4066 2544 4122 2553
rect 4066 2479 4068 2488
rect 4120 2479 4122 2488
rect 4068 2450 4120 2456
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3700 2032 3752 2038
rect 3700 1974 3752 1980
rect 20 1828 72 1834
rect 20 1770 72 1776
rect 32 400 60 1770
rect 3112 1660 3420 1669
rect 3112 1658 3118 1660
rect 3174 1658 3198 1660
rect 3254 1658 3278 1660
rect 3334 1658 3358 1660
rect 3414 1658 3420 1660
rect 3174 1606 3176 1658
rect 3356 1606 3358 1658
rect 3112 1604 3118 1606
rect 3174 1604 3198 1606
rect 3254 1604 3278 1606
rect 3334 1604 3358 1606
rect 3414 1604 3420 1606
rect 3112 1595 3420 1604
rect 1755 1116 2063 1125
rect 1755 1114 1761 1116
rect 1817 1114 1841 1116
rect 1897 1114 1921 1116
rect 1977 1114 2001 1116
rect 2057 1114 2063 1116
rect 1817 1062 1819 1114
rect 1999 1062 2001 1114
rect 1755 1060 1761 1062
rect 1817 1060 1841 1062
rect 1897 1060 1921 1062
rect 1977 1060 2001 1062
rect 2057 1060 2063 1062
rect 1755 1051 2063 1060
rect 3712 1018 3740 1974
rect 3804 1562 3832 2382
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4252 2304 4304 2310
rect 4252 2246 4304 2252
rect 4080 1902 4108 2246
rect 4068 1896 4120 1902
rect 4068 1838 4120 1844
rect 4172 1766 4200 2246
rect 4264 1902 4292 2246
rect 4356 1986 4384 2926
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5552 2553 5580 2790
rect 5644 2650 5672 3334
rect 5736 2854 5764 3470
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5826 2748 6134 2757
rect 5826 2746 5832 2748
rect 5888 2746 5912 2748
rect 5968 2746 5992 2748
rect 6048 2746 6072 2748
rect 6128 2746 6134 2748
rect 5888 2694 5890 2746
rect 6070 2694 6072 2746
rect 5826 2692 5832 2694
rect 5888 2692 5912 2694
rect 5968 2692 5992 2694
rect 6048 2692 6072 2694
rect 6128 2692 6134 2694
rect 5826 2683 6134 2692
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5538 2544 5594 2553
rect 4896 2508 4948 2514
rect 6196 2514 6224 2926
rect 5538 2479 5540 2488
rect 4896 2450 4948 2456
rect 5592 2479 5594 2488
rect 6184 2508 6236 2514
rect 5540 2450 5592 2456
rect 6184 2450 6236 2456
rect 4469 2204 4777 2213
rect 4469 2202 4475 2204
rect 4531 2202 4555 2204
rect 4611 2202 4635 2204
rect 4691 2202 4715 2204
rect 4771 2202 4777 2204
rect 4531 2150 4533 2202
rect 4713 2150 4715 2202
rect 4469 2148 4475 2150
rect 4531 2148 4555 2150
rect 4611 2148 4635 2150
rect 4691 2148 4715 2150
rect 4771 2148 4777 2150
rect 4469 2139 4777 2148
rect 4356 1970 4568 1986
rect 4908 1970 4936 2450
rect 6288 2446 6316 3606
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 5540 2304 5592 2310
rect 6288 2258 6316 2382
rect 6380 2310 6408 3334
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 6748 2650 6776 2790
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6840 2530 6868 3674
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8944 3528 8996 3534
rect 11244 3528 11296 3534
rect 8944 3470 8996 3476
rect 11242 3496 11244 3505
rect 11296 3496 11298 3505
rect 7183 3292 7491 3301
rect 7183 3290 7189 3292
rect 7245 3290 7269 3292
rect 7325 3290 7349 3292
rect 7405 3290 7429 3292
rect 7485 3290 7491 3292
rect 7245 3238 7247 3290
rect 7427 3238 7429 3290
rect 7183 3236 7189 3238
rect 7245 3236 7269 3238
rect 7325 3236 7349 3238
rect 7405 3236 7429 3238
rect 7485 3236 7491 3238
rect 7183 3227 7491 3236
rect 8128 3194 8156 3470
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 6656 2514 6868 2530
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 6644 2508 6868 2514
rect 6696 2502 6868 2508
rect 6644 2450 6696 2456
rect 5540 2246 5592 2252
rect 4356 1964 4580 1970
rect 4356 1958 4528 1964
rect 4528 1906 4580 1912
rect 4896 1964 4948 1970
rect 4896 1906 4948 1912
rect 4252 1896 4304 1902
rect 4252 1838 4304 1844
rect 4988 1896 5040 1902
rect 4988 1838 5040 1844
rect 4160 1760 4212 1766
rect 4160 1702 4212 1708
rect 3792 1556 3844 1562
rect 3792 1498 3844 1504
rect 4172 1426 4200 1702
rect 5000 1562 5028 1838
rect 4988 1556 5040 1562
rect 4988 1498 5040 1504
rect 4160 1420 4212 1426
rect 4160 1362 4212 1368
rect 5552 1358 5580 2246
rect 6196 2230 6316 2258
rect 6368 2304 6420 2310
rect 6368 2246 6420 2252
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6196 1766 6224 2230
rect 6184 1760 6236 1766
rect 6184 1702 6236 1708
rect 5826 1660 6134 1669
rect 5826 1658 5832 1660
rect 5888 1658 5912 1660
rect 5968 1658 5992 1660
rect 6048 1658 6072 1660
rect 6128 1658 6134 1660
rect 5888 1606 5890 1658
rect 6070 1606 6072 1658
rect 5826 1604 5832 1606
rect 5888 1604 5912 1606
rect 5968 1604 5992 1606
rect 6048 1604 6072 1606
rect 6128 1604 6134 1606
rect 5826 1595 6134 1604
rect 6196 1426 6224 1702
rect 6184 1420 6236 1426
rect 6184 1362 6236 1368
rect 5540 1352 5592 1358
rect 5540 1294 5592 1300
rect 6840 1222 6868 2246
rect 7024 2106 7052 2518
rect 7012 2100 7064 2106
rect 7012 2042 7064 2048
rect 6920 1760 6972 1766
rect 6920 1702 6972 1708
rect 6932 1494 6960 1702
rect 6920 1488 6972 1494
rect 6920 1430 6972 1436
rect 6828 1216 6880 1222
rect 6828 1158 6880 1164
rect 4469 1116 4777 1125
rect 4469 1114 4475 1116
rect 4531 1114 4555 1116
rect 4611 1114 4635 1116
rect 4691 1114 4715 1116
rect 4771 1114 4777 1116
rect 4531 1062 4533 1114
rect 4713 1062 4715 1114
rect 4469 1060 4475 1062
rect 4531 1060 4555 1062
rect 4611 1060 4635 1062
rect 4691 1060 4715 1062
rect 4771 1060 4777 1062
rect 4469 1051 4777 1060
rect 3700 1012 3752 1018
rect 3700 954 3752 960
rect 6932 814 6960 1430
rect 6920 808 6972 814
rect 6920 750 6972 756
rect 7116 746 7144 2790
rect 8312 2582 8340 2790
rect 8404 2650 8432 2790
rect 8540 2748 8848 2757
rect 8540 2746 8546 2748
rect 8602 2746 8626 2748
rect 8682 2746 8706 2748
rect 8762 2746 8786 2748
rect 8842 2746 8848 2748
rect 8602 2694 8604 2746
rect 8784 2694 8786 2746
rect 8540 2692 8546 2694
rect 8602 2692 8626 2694
rect 8682 2692 8706 2694
rect 8762 2692 8786 2694
rect 8842 2692 8848 2694
rect 8540 2683 8848 2692
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8956 2446 8984 3470
rect 11242 3431 11298 3440
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 9897 3292 10205 3301
rect 9897 3290 9903 3292
rect 9959 3290 9983 3292
rect 10039 3290 10063 3292
rect 10119 3290 10143 3292
rect 10199 3290 10205 3292
rect 9959 3238 9961 3290
rect 10141 3238 10143 3290
rect 9897 3236 9903 3238
rect 9959 3236 9983 3238
rect 10039 3236 10063 3238
rect 10119 3236 10143 3238
rect 10199 3236 10205 3238
rect 9897 3227 10205 3236
rect 10612 3194 10640 3334
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 11254 2748 11562 2757
rect 11254 2746 11260 2748
rect 11316 2746 11340 2748
rect 11396 2746 11420 2748
rect 11476 2746 11500 2748
rect 11556 2746 11562 2748
rect 11316 2694 11318 2746
rect 11498 2694 11500 2746
rect 11254 2692 11260 2694
rect 11316 2692 11340 2694
rect 11396 2692 11420 2694
rect 11476 2692 11500 2694
rect 11556 2692 11562 2694
rect 11254 2683 11562 2692
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 7183 2204 7491 2213
rect 7183 2202 7189 2204
rect 7245 2202 7269 2204
rect 7325 2202 7349 2204
rect 7405 2202 7429 2204
rect 7485 2202 7491 2204
rect 7245 2150 7247 2202
rect 7427 2150 7429 2202
rect 7183 2148 7189 2150
rect 7245 2148 7269 2150
rect 7325 2148 7349 2150
rect 7405 2148 7429 2150
rect 7485 2148 7491 2150
rect 7183 2139 7491 2148
rect 8540 1660 8848 1669
rect 8540 1658 8546 1660
rect 8602 1658 8626 1660
rect 8682 1658 8706 1660
rect 8762 1658 8786 1660
rect 8842 1658 8848 1660
rect 8602 1606 8604 1658
rect 8784 1606 8786 1658
rect 8540 1604 8546 1606
rect 8602 1604 8626 1606
rect 8682 1604 8706 1606
rect 8762 1604 8786 1606
rect 8842 1604 8848 1606
rect 8540 1595 8848 1604
rect 8956 1442 8984 2382
rect 9897 2204 10205 2213
rect 9897 2202 9903 2204
rect 9959 2202 9983 2204
rect 10039 2202 10063 2204
rect 10119 2202 10143 2204
rect 10199 2202 10205 2204
rect 9959 2150 9961 2202
rect 10141 2150 10143 2202
rect 9897 2148 9903 2150
rect 9959 2148 9983 2150
rect 10039 2148 10063 2150
rect 10119 2148 10143 2150
rect 10199 2148 10205 2150
rect 9897 2139 10205 2148
rect 11254 1660 11562 1669
rect 11254 1658 11260 1660
rect 11316 1658 11340 1660
rect 11396 1658 11420 1660
rect 11476 1658 11500 1660
rect 11556 1658 11562 1660
rect 11316 1606 11318 1658
rect 11498 1606 11500 1658
rect 11254 1604 11260 1606
rect 11316 1604 11340 1606
rect 11396 1604 11420 1606
rect 11476 1604 11500 1606
rect 11556 1604 11562 1606
rect 11254 1595 11562 1604
rect 8864 1414 8984 1442
rect 8864 1358 8892 1414
rect 7656 1352 7708 1358
rect 7656 1294 7708 1300
rect 8852 1352 8904 1358
rect 8852 1294 8904 1300
rect 7183 1116 7491 1125
rect 7183 1114 7189 1116
rect 7245 1114 7269 1116
rect 7325 1114 7349 1116
rect 7405 1114 7429 1116
rect 7485 1114 7491 1116
rect 7245 1062 7247 1114
rect 7427 1062 7429 1114
rect 7183 1060 7189 1062
rect 7245 1060 7269 1062
rect 7325 1060 7349 1062
rect 7405 1060 7429 1062
rect 7485 1060 7491 1062
rect 7183 1051 7491 1060
rect 7668 1018 7696 1294
rect 7748 1216 7800 1222
rect 7748 1158 7800 1164
rect 7656 1012 7708 1018
rect 7656 954 7708 960
rect 7760 814 7788 1158
rect 8864 1018 8892 1294
rect 9897 1116 10205 1125
rect 9897 1114 9903 1116
rect 9959 1114 9983 1116
rect 10039 1114 10063 1116
rect 10119 1114 10143 1116
rect 10199 1114 10205 1116
rect 9959 1062 9961 1114
rect 10141 1062 10143 1114
rect 9897 1060 9903 1062
rect 9959 1060 9983 1062
rect 10039 1060 10063 1062
rect 10119 1060 10143 1062
rect 10199 1060 10205 1062
rect 9897 1051 10205 1060
rect 8852 1012 8904 1018
rect 8852 954 8904 960
rect 7748 808 7800 814
rect 7748 750 7800 756
rect 7104 740 7156 746
rect 7104 682 7156 688
rect 3112 572 3420 581
rect 3112 570 3118 572
rect 3174 570 3198 572
rect 3254 570 3278 572
rect 3334 570 3358 572
rect 3414 570 3420 572
rect 3174 518 3176 570
rect 3356 518 3358 570
rect 3112 516 3118 518
rect 3174 516 3198 518
rect 3254 516 3278 518
rect 3334 516 3358 518
rect 3414 516 3420 518
rect 3112 507 3420 516
rect 5826 572 6134 581
rect 5826 570 5832 572
rect 5888 570 5912 572
rect 5968 570 5992 572
rect 6048 570 6072 572
rect 6128 570 6134 572
rect 5888 518 5890 570
rect 6070 518 6072 570
rect 5826 516 5832 518
rect 5888 516 5912 518
rect 5968 516 5992 518
rect 6048 516 6072 518
rect 6128 516 6134 518
rect 5826 507 6134 516
rect 7760 400 7788 750
rect 8540 572 8848 581
rect 8540 570 8546 572
rect 8602 570 8626 572
rect 8682 570 8706 572
rect 8762 570 8786 572
rect 8842 570 8848 572
rect 8602 518 8604 570
rect 8784 518 8786 570
rect 8540 516 8546 518
rect 8602 516 8626 518
rect 8682 516 8706 518
rect 8762 516 8786 518
rect 8842 516 8848 518
rect 8540 507 8848 516
rect 11254 572 11562 581
rect 11254 570 11260 572
rect 11316 570 11340 572
rect 11396 570 11420 572
rect 11476 570 11500 572
rect 11556 570 11562 572
rect 11316 518 11318 570
rect 11498 518 11500 570
rect 11254 516 11260 518
rect 11316 516 11340 518
rect 11396 516 11420 518
rect 11476 516 11500 518
rect 11556 516 11562 518
rect 11254 507 11562 516
rect 18 0 74 400
rect 7746 0 7802 400
<< via2 >>
rect 3118 11450 3174 11452
rect 3198 11450 3254 11452
rect 3278 11450 3334 11452
rect 3358 11450 3414 11452
rect 3118 11398 3164 11450
rect 3164 11398 3174 11450
rect 3198 11398 3228 11450
rect 3228 11398 3240 11450
rect 3240 11398 3254 11450
rect 3278 11398 3292 11450
rect 3292 11398 3304 11450
rect 3304 11398 3334 11450
rect 3358 11398 3368 11450
rect 3368 11398 3414 11450
rect 3118 11396 3174 11398
rect 3198 11396 3254 11398
rect 3278 11396 3334 11398
rect 3358 11396 3414 11398
rect 1761 10906 1817 10908
rect 1841 10906 1897 10908
rect 1921 10906 1977 10908
rect 2001 10906 2057 10908
rect 1761 10854 1807 10906
rect 1807 10854 1817 10906
rect 1841 10854 1871 10906
rect 1871 10854 1883 10906
rect 1883 10854 1897 10906
rect 1921 10854 1935 10906
rect 1935 10854 1947 10906
rect 1947 10854 1977 10906
rect 2001 10854 2011 10906
rect 2011 10854 2057 10906
rect 1761 10852 1817 10854
rect 1841 10852 1897 10854
rect 1921 10852 1977 10854
rect 2001 10852 2057 10854
rect 3118 10362 3174 10364
rect 3198 10362 3254 10364
rect 3278 10362 3334 10364
rect 3358 10362 3414 10364
rect 3118 10310 3164 10362
rect 3164 10310 3174 10362
rect 3198 10310 3228 10362
rect 3228 10310 3240 10362
rect 3240 10310 3254 10362
rect 3278 10310 3292 10362
rect 3292 10310 3304 10362
rect 3304 10310 3334 10362
rect 3358 10310 3368 10362
rect 3368 10310 3414 10362
rect 3118 10308 3174 10310
rect 3198 10308 3254 10310
rect 3278 10308 3334 10310
rect 3358 10308 3414 10310
rect 1761 9818 1817 9820
rect 1841 9818 1897 9820
rect 1921 9818 1977 9820
rect 2001 9818 2057 9820
rect 1761 9766 1807 9818
rect 1807 9766 1817 9818
rect 1841 9766 1871 9818
rect 1871 9766 1883 9818
rect 1883 9766 1897 9818
rect 1921 9766 1935 9818
rect 1935 9766 1947 9818
rect 1947 9766 1977 9818
rect 2001 9766 2011 9818
rect 2011 9766 2057 9818
rect 1761 9764 1817 9766
rect 1841 9764 1897 9766
rect 1921 9764 1977 9766
rect 2001 9764 2057 9766
rect 3118 9274 3174 9276
rect 3198 9274 3254 9276
rect 3278 9274 3334 9276
rect 3358 9274 3414 9276
rect 3118 9222 3164 9274
rect 3164 9222 3174 9274
rect 3198 9222 3228 9274
rect 3228 9222 3240 9274
rect 3240 9222 3254 9274
rect 3278 9222 3292 9274
rect 3292 9222 3304 9274
rect 3304 9222 3334 9274
rect 3358 9222 3368 9274
rect 3368 9222 3414 9274
rect 3118 9220 3174 9222
rect 3198 9220 3254 9222
rect 3278 9220 3334 9222
rect 3358 9220 3414 9222
rect 1761 8730 1817 8732
rect 1841 8730 1897 8732
rect 1921 8730 1977 8732
rect 2001 8730 2057 8732
rect 1761 8678 1807 8730
rect 1807 8678 1817 8730
rect 1841 8678 1871 8730
rect 1871 8678 1883 8730
rect 1883 8678 1897 8730
rect 1921 8678 1935 8730
rect 1935 8678 1947 8730
rect 1947 8678 1977 8730
rect 2001 8678 2011 8730
rect 2011 8678 2057 8730
rect 1761 8676 1817 8678
rect 1841 8676 1897 8678
rect 1921 8676 1977 8678
rect 2001 8676 2057 8678
rect 2778 8200 2834 8256
rect 1761 7642 1817 7644
rect 1841 7642 1897 7644
rect 1921 7642 1977 7644
rect 2001 7642 2057 7644
rect 1761 7590 1807 7642
rect 1807 7590 1817 7642
rect 1841 7590 1871 7642
rect 1871 7590 1883 7642
rect 1883 7590 1897 7642
rect 1921 7590 1935 7642
rect 1935 7590 1947 7642
rect 1947 7590 1977 7642
rect 2001 7590 2011 7642
rect 2011 7590 2057 7642
rect 1761 7588 1817 7590
rect 1841 7588 1897 7590
rect 1921 7588 1977 7590
rect 2001 7588 2057 7590
rect 3118 8186 3174 8188
rect 3198 8186 3254 8188
rect 3278 8186 3334 8188
rect 3358 8186 3414 8188
rect 3118 8134 3164 8186
rect 3164 8134 3174 8186
rect 3198 8134 3228 8186
rect 3228 8134 3240 8186
rect 3240 8134 3254 8186
rect 3278 8134 3292 8186
rect 3292 8134 3304 8186
rect 3304 8134 3334 8186
rect 3358 8134 3368 8186
rect 3368 8134 3414 8186
rect 3118 8132 3174 8134
rect 3198 8132 3254 8134
rect 3278 8132 3334 8134
rect 3358 8132 3414 8134
rect 3118 7098 3174 7100
rect 3198 7098 3254 7100
rect 3278 7098 3334 7100
rect 3358 7098 3414 7100
rect 3118 7046 3164 7098
rect 3164 7046 3174 7098
rect 3198 7046 3228 7098
rect 3228 7046 3240 7098
rect 3240 7046 3254 7098
rect 3278 7046 3292 7098
rect 3292 7046 3304 7098
rect 3304 7046 3334 7098
rect 3358 7046 3368 7098
rect 3368 7046 3414 7098
rect 3118 7044 3174 7046
rect 3198 7044 3254 7046
rect 3278 7044 3334 7046
rect 3358 7044 3414 7046
rect 5832 11450 5888 11452
rect 5912 11450 5968 11452
rect 5992 11450 6048 11452
rect 6072 11450 6128 11452
rect 5832 11398 5878 11450
rect 5878 11398 5888 11450
rect 5912 11398 5942 11450
rect 5942 11398 5954 11450
rect 5954 11398 5968 11450
rect 5992 11398 6006 11450
rect 6006 11398 6018 11450
rect 6018 11398 6048 11450
rect 6072 11398 6082 11450
rect 6082 11398 6128 11450
rect 5832 11396 5888 11398
rect 5912 11396 5968 11398
rect 5992 11396 6048 11398
rect 6072 11396 6128 11398
rect 8546 11450 8602 11452
rect 8626 11450 8682 11452
rect 8706 11450 8762 11452
rect 8786 11450 8842 11452
rect 8546 11398 8592 11450
rect 8592 11398 8602 11450
rect 8626 11398 8656 11450
rect 8656 11398 8668 11450
rect 8668 11398 8682 11450
rect 8706 11398 8720 11450
rect 8720 11398 8732 11450
rect 8732 11398 8762 11450
rect 8786 11398 8796 11450
rect 8796 11398 8842 11450
rect 8546 11396 8602 11398
rect 8626 11396 8682 11398
rect 8706 11396 8762 11398
rect 8786 11396 8842 11398
rect 11260 11450 11316 11452
rect 11340 11450 11396 11452
rect 11420 11450 11476 11452
rect 11500 11450 11556 11452
rect 11260 11398 11306 11450
rect 11306 11398 11316 11450
rect 11340 11398 11370 11450
rect 11370 11398 11382 11450
rect 11382 11398 11396 11450
rect 11420 11398 11434 11450
rect 11434 11398 11446 11450
rect 11446 11398 11476 11450
rect 11500 11398 11510 11450
rect 11510 11398 11556 11450
rect 11260 11396 11316 11398
rect 11340 11396 11396 11398
rect 11420 11396 11476 11398
rect 11500 11396 11556 11398
rect 4475 10906 4531 10908
rect 4555 10906 4611 10908
rect 4635 10906 4691 10908
rect 4715 10906 4771 10908
rect 4475 10854 4521 10906
rect 4521 10854 4531 10906
rect 4555 10854 4585 10906
rect 4585 10854 4597 10906
rect 4597 10854 4611 10906
rect 4635 10854 4649 10906
rect 4649 10854 4661 10906
rect 4661 10854 4691 10906
rect 4715 10854 4725 10906
rect 4725 10854 4771 10906
rect 4475 10852 4531 10854
rect 4555 10852 4611 10854
rect 4635 10852 4691 10854
rect 4715 10852 4771 10854
rect 7189 10906 7245 10908
rect 7269 10906 7325 10908
rect 7349 10906 7405 10908
rect 7429 10906 7485 10908
rect 7189 10854 7235 10906
rect 7235 10854 7245 10906
rect 7269 10854 7299 10906
rect 7299 10854 7311 10906
rect 7311 10854 7325 10906
rect 7349 10854 7363 10906
rect 7363 10854 7375 10906
rect 7375 10854 7405 10906
rect 7429 10854 7439 10906
rect 7439 10854 7485 10906
rect 7189 10852 7245 10854
rect 7269 10852 7325 10854
rect 7349 10852 7405 10854
rect 7429 10852 7485 10854
rect 9903 10906 9959 10908
rect 9983 10906 10039 10908
rect 10063 10906 10119 10908
rect 10143 10906 10199 10908
rect 9903 10854 9949 10906
rect 9949 10854 9959 10906
rect 9983 10854 10013 10906
rect 10013 10854 10025 10906
rect 10025 10854 10039 10906
rect 10063 10854 10077 10906
rect 10077 10854 10089 10906
rect 10089 10854 10119 10906
rect 10143 10854 10153 10906
rect 10153 10854 10199 10906
rect 9903 10852 9959 10854
rect 9983 10852 10039 10854
rect 10063 10852 10119 10854
rect 10143 10852 10199 10854
rect 5832 10362 5888 10364
rect 5912 10362 5968 10364
rect 5992 10362 6048 10364
rect 6072 10362 6128 10364
rect 5832 10310 5878 10362
rect 5878 10310 5888 10362
rect 5912 10310 5942 10362
rect 5942 10310 5954 10362
rect 5954 10310 5968 10362
rect 5992 10310 6006 10362
rect 6006 10310 6018 10362
rect 6018 10310 6048 10362
rect 6072 10310 6082 10362
rect 6082 10310 6128 10362
rect 5832 10308 5888 10310
rect 5912 10308 5968 10310
rect 5992 10308 6048 10310
rect 6072 10308 6128 10310
rect 8546 10362 8602 10364
rect 8626 10362 8682 10364
rect 8706 10362 8762 10364
rect 8786 10362 8842 10364
rect 8546 10310 8592 10362
rect 8592 10310 8602 10362
rect 8626 10310 8656 10362
rect 8656 10310 8668 10362
rect 8668 10310 8682 10362
rect 8706 10310 8720 10362
rect 8720 10310 8732 10362
rect 8732 10310 8762 10362
rect 8786 10310 8796 10362
rect 8796 10310 8842 10362
rect 8546 10308 8602 10310
rect 8626 10308 8682 10310
rect 8706 10308 8762 10310
rect 8786 10308 8842 10310
rect 11260 10362 11316 10364
rect 11340 10362 11396 10364
rect 11420 10362 11476 10364
rect 11500 10362 11556 10364
rect 11260 10310 11306 10362
rect 11306 10310 11316 10362
rect 11340 10310 11370 10362
rect 11370 10310 11382 10362
rect 11382 10310 11396 10362
rect 11420 10310 11434 10362
rect 11434 10310 11446 10362
rect 11446 10310 11476 10362
rect 11500 10310 11510 10362
rect 11510 10310 11556 10362
rect 11260 10308 11316 10310
rect 11340 10308 11396 10310
rect 11420 10308 11476 10310
rect 11500 10308 11556 10310
rect 4475 9818 4531 9820
rect 4555 9818 4611 9820
rect 4635 9818 4691 9820
rect 4715 9818 4771 9820
rect 4475 9766 4521 9818
rect 4521 9766 4531 9818
rect 4555 9766 4585 9818
rect 4585 9766 4597 9818
rect 4597 9766 4611 9818
rect 4635 9766 4649 9818
rect 4649 9766 4661 9818
rect 4661 9766 4691 9818
rect 4715 9766 4725 9818
rect 4725 9766 4771 9818
rect 4475 9764 4531 9766
rect 4555 9764 4611 9766
rect 4635 9764 4691 9766
rect 4715 9764 4771 9766
rect 7189 9818 7245 9820
rect 7269 9818 7325 9820
rect 7349 9818 7405 9820
rect 7429 9818 7485 9820
rect 7189 9766 7235 9818
rect 7235 9766 7245 9818
rect 7269 9766 7299 9818
rect 7299 9766 7311 9818
rect 7311 9766 7325 9818
rect 7349 9766 7363 9818
rect 7363 9766 7375 9818
rect 7375 9766 7405 9818
rect 7429 9766 7439 9818
rect 7439 9766 7485 9818
rect 7189 9764 7245 9766
rect 7269 9764 7325 9766
rect 7349 9764 7405 9766
rect 7429 9764 7485 9766
rect 9903 9818 9959 9820
rect 9983 9818 10039 9820
rect 10063 9818 10119 9820
rect 10143 9818 10199 9820
rect 9903 9766 9949 9818
rect 9949 9766 9959 9818
rect 9983 9766 10013 9818
rect 10013 9766 10025 9818
rect 10025 9766 10039 9818
rect 10063 9766 10077 9818
rect 10077 9766 10089 9818
rect 10089 9766 10119 9818
rect 10143 9766 10153 9818
rect 10153 9766 10199 9818
rect 9903 9764 9959 9766
rect 9983 9764 10039 9766
rect 10063 9764 10119 9766
rect 10143 9764 10199 9766
rect 5832 9274 5888 9276
rect 5912 9274 5968 9276
rect 5992 9274 6048 9276
rect 6072 9274 6128 9276
rect 5832 9222 5878 9274
rect 5878 9222 5888 9274
rect 5912 9222 5942 9274
rect 5942 9222 5954 9274
rect 5954 9222 5968 9274
rect 5992 9222 6006 9274
rect 6006 9222 6018 9274
rect 6018 9222 6048 9274
rect 6072 9222 6082 9274
rect 6082 9222 6128 9274
rect 5832 9220 5888 9222
rect 5912 9220 5968 9222
rect 5992 9220 6048 9222
rect 6072 9220 6128 9222
rect 8546 9274 8602 9276
rect 8626 9274 8682 9276
rect 8706 9274 8762 9276
rect 8786 9274 8842 9276
rect 8546 9222 8592 9274
rect 8592 9222 8602 9274
rect 8626 9222 8656 9274
rect 8656 9222 8668 9274
rect 8668 9222 8682 9274
rect 8706 9222 8720 9274
rect 8720 9222 8732 9274
rect 8732 9222 8762 9274
rect 8786 9222 8796 9274
rect 8796 9222 8842 9274
rect 8546 9220 8602 9222
rect 8626 9220 8682 9222
rect 8706 9220 8762 9222
rect 8786 9220 8842 9222
rect 11260 9274 11316 9276
rect 11340 9274 11396 9276
rect 11420 9274 11476 9276
rect 11500 9274 11556 9276
rect 11260 9222 11306 9274
rect 11306 9222 11316 9274
rect 11340 9222 11370 9274
rect 11370 9222 11382 9274
rect 11382 9222 11396 9274
rect 11420 9222 11434 9274
rect 11434 9222 11446 9274
rect 11446 9222 11476 9274
rect 11500 9222 11510 9274
rect 11510 9222 11556 9274
rect 11260 9220 11316 9222
rect 11340 9220 11396 9222
rect 11420 9220 11476 9222
rect 11500 9220 11556 9222
rect 4475 8730 4531 8732
rect 4555 8730 4611 8732
rect 4635 8730 4691 8732
rect 4715 8730 4771 8732
rect 4475 8678 4521 8730
rect 4521 8678 4531 8730
rect 4555 8678 4585 8730
rect 4585 8678 4597 8730
rect 4597 8678 4611 8730
rect 4635 8678 4649 8730
rect 4649 8678 4661 8730
rect 4661 8678 4691 8730
rect 4715 8678 4725 8730
rect 4725 8678 4771 8730
rect 4475 8676 4531 8678
rect 4555 8676 4611 8678
rect 4635 8676 4691 8678
rect 4715 8676 4771 8678
rect 7189 8730 7245 8732
rect 7269 8730 7325 8732
rect 7349 8730 7405 8732
rect 7429 8730 7485 8732
rect 7189 8678 7235 8730
rect 7235 8678 7245 8730
rect 7269 8678 7299 8730
rect 7299 8678 7311 8730
rect 7311 8678 7325 8730
rect 7349 8678 7363 8730
rect 7363 8678 7375 8730
rect 7375 8678 7405 8730
rect 7429 8678 7439 8730
rect 7439 8678 7485 8730
rect 7189 8676 7245 8678
rect 7269 8676 7325 8678
rect 7349 8676 7405 8678
rect 7429 8676 7485 8678
rect 9903 8730 9959 8732
rect 9983 8730 10039 8732
rect 10063 8730 10119 8732
rect 10143 8730 10199 8732
rect 9903 8678 9949 8730
rect 9949 8678 9959 8730
rect 9983 8678 10013 8730
rect 10013 8678 10025 8730
rect 10025 8678 10039 8730
rect 10063 8678 10077 8730
rect 10077 8678 10089 8730
rect 10089 8678 10119 8730
rect 10143 8678 10153 8730
rect 10153 8678 10199 8730
rect 9903 8676 9959 8678
rect 9983 8676 10039 8678
rect 10063 8676 10119 8678
rect 10143 8676 10199 8678
rect 5832 8186 5888 8188
rect 5912 8186 5968 8188
rect 5992 8186 6048 8188
rect 6072 8186 6128 8188
rect 5832 8134 5878 8186
rect 5878 8134 5888 8186
rect 5912 8134 5942 8186
rect 5942 8134 5954 8186
rect 5954 8134 5968 8186
rect 5992 8134 6006 8186
rect 6006 8134 6018 8186
rect 6018 8134 6048 8186
rect 6072 8134 6082 8186
rect 6082 8134 6128 8186
rect 5832 8132 5888 8134
rect 5912 8132 5968 8134
rect 5992 8132 6048 8134
rect 6072 8132 6128 8134
rect 8546 8186 8602 8188
rect 8626 8186 8682 8188
rect 8706 8186 8762 8188
rect 8786 8186 8842 8188
rect 8546 8134 8592 8186
rect 8592 8134 8602 8186
rect 8626 8134 8656 8186
rect 8656 8134 8668 8186
rect 8668 8134 8682 8186
rect 8706 8134 8720 8186
rect 8720 8134 8732 8186
rect 8732 8134 8762 8186
rect 8786 8134 8796 8186
rect 8796 8134 8842 8186
rect 8546 8132 8602 8134
rect 8626 8132 8682 8134
rect 8706 8132 8762 8134
rect 8786 8132 8842 8134
rect 11260 8186 11316 8188
rect 11340 8186 11396 8188
rect 11420 8186 11476 8188
rect 11500 8186 11556 8188
rect 11260 8134 11306 8186
rect 11306 8134 11316 8186
rect 11340 8134 11370 8186
rect 11370 8134 11382 8186
rect 11382 8134 11396 8186
rect 11420 8134 11434 8186
rect 11434 8134 11446 8186
rect 11446 8134 11476 8186
rect 11500 8134 11510 8186
rect 11510 8134 11556 8186
rect 11260 8132 11316 8134
rect 11340 8132 11396 8134
rect 11420 8132 11476 8134
rect 11500 8132 11556 8134
rect 4475 7642 4531 7644
rect 4555 7642 4611 7644
rect 4635 7642 4691 7644
rect 4715 7642 4771 7644
rect 4475 7590 4521 7642
rect 4521 7590 4531 7642
rect 4555 7590 4585 7642
rect 4585 7590 4597 7642
rect 4597 7590 4611 7642
rect 4635 7590 4649 7642
rect 4649 7590 4661 7642
rect 4661 7590 4691 7642
rect 4715 7590 4725 7642
rect 4725 7590 4771 7642
rect 4475 7588 4531 7590
rect 4555 7588 4611 7590
rect 4635 7588 4691 7590
rect 4715 7588 4771 7590
rect 7189 7642 7245 7644
rect 7269 7642 7325 7644
rect 7349 7642 7405 7644
rect 7429 7642 7485 7644
rect 7189 7590 7235 7642
rect 7235 7590 7245 7642
rect 7269 7590 7299 7642
rect 7299 7590 7311 7642
rect 7311 7590 7325 7642
rect 7349 7590 7363 7642
rect 7363 7590 7375 7642
rect 7375 7590 7405 7642
rect 7429 7590 7439 7642
rect 7439 7590 7485 7642
rect 7189 7588 7245 7590
rect 7269 7588 7325 7590
rect 7349 7588 7405 7590
rect 7429 7588 7485 7590
rect 9903 7642 9959 7644
rect 9983 7642 10039 7644
rect 10063 7642 10119 7644
rect 10143 7642 10199 7644
rect 9903 7590 9949 7642
rect 9949 7590 9959 7642
rect 9983 7590 10013 7642
rect 10013 7590 10025 7642
rect 10025 7590 10039 7642
rect 10063 7590 10077 7642
rect 10077 7590 10089 7642
rect 10089 7590 10119 7642
rect 10143 7590 10153 7642
rect 10153 7590 10199 7642
rect 9903 7588 9959 7590
rect 9983 7588 10039 7590
rect 10063 7588 10119 7590
rect 10143 7588 10199 7590
rect 1761 6554 1817 6556
rect 1841 6554 1897 6556
rect 1921 6554 1977 6556
rect 2001 6554 2057 6556
rect 1761 6502 1807 6554
rect 1807 6502 1817 6554
rect 1841 6502 1871 6554
rect 1871 6502 1883 6554
rect 1883 6502 1897 6554
rect 1921 6502 1935 6554
rect 1935 6502 1947 6554
rect 1947 6502 1977 6554
rect 2001 6502 2011 6554
rect 2011 6502 2057 6554
rect 1761 6500 1817 6502
rect 1841 6500 1897 6502
rect 1921 6500 1977 6502
rect 2001 6500 2057 6502
rect 3118 6010 3174 6012
rect 3198 6010 3254 6012
rect 3278 6010 3334 6012
rect 3358 6010 3414 6012
rect 3118 5958 3164 6010
rect 3164 5958 3174 6010
rect 3198 5958 3228 6010
rect 3228 5958 3240 6010
rect 3240 5958 3254 6010
rect 3278 5958 3292 6010
rect 3292 5958 3304 6010
rect 3304 5958 3334 6010
rect 3358 5958 3368 6010
rect 3368 5958 3414 6010
rect 3118 5956 3174 5958
rect 3198 5956 3254 5958
rect 3278 5956 3334 5958
rect 3358 5956 3414 5958
rect 1761 5466 1817 5468
rect 1841 5466 1897 5468
rect 1921 5466 1977 5468
rect 2001 5466 2057 5468
rect 1761 5414 1807 5466
rect 1807 5414 1817 5466
rect 1841 5414 1871 5466
rect 1871 5414 1883 5466
rect 1883 5414 1897 5466
rect 1921 5414 1935 5466
rect 1935 5414 1947 5466
rect 1947 5414 1977 5466
rect 2001 5414 2011 5466
rect 2011 5414 2057 5466
rect 1761 5412 1817 5414
rect 1841 5412 1897 5414
rect 1921 5412 1977 5414
rect 2001 5412 2057 5414
rect 3118 4922 3174 4924
rect 3198 4922 3254 4924
rect 3278 4922 3334 4924
rect 3358 4922 3414 4924
rect 3118 4870 3164 4922
rect 3164 4870 3174 4922
rect 3198 4870 3228 4922
rect 3228 4870 3240 4922
rect 3240 4870 3254 4922
rect 3278 4870 3292 4922
rect 3292 4870 3304 4922
rect 3304 4870 3334 4922
rect 3358 4870 3368 4922
rect 3368 4870 3414 4922
rect 3118 4868 3174 4870
rect 3198 4868 3254 4870
rect 3278 4868 3334 4870
rect 3358 4868 3414 4870
rect 1761 4378 1817 4380
rect 1841 4378 1897 4380
rect 1921 4378 1977 4380
rect 2001 4378 2057 4380
rect 1761 4326 1807 4378
rect 1807 4326 1817 4378
rect 1841 4326 1871 4378
rect 1871 4326 1883 4378
rect 1883 4326 1897 4378
rect 1921 4326 1935 4378
rect 1935 4326 1947 4378
rect 1947 4326 1977 4378
rect 2001 4326 2011 4378
rect 2011 4326 2057 4378
rect 1761 4324 1817 4326
rect 1841 4324 1897 4326
rect 1921 4324 1977 4326
rect 2001 4324 2057 4326
rect 3118 3834 3174 3836
rect 3198 3834 3254 3836
rect 3278 3834 3334 3836
rect 3358 3834 3414 3836
rect 3118 3782 3164 3834
rect 3164 3782 3174 3834
rect 3198 3782 3228 3834
rect 3228 3782 3240 3834
rect 3240 3782 3254 3834
rect 3278 3782 3292 3834
rect 3292 3782 3304 3834
rect 3304 3782 3334 3834
rect 3358 3782 3368 3834
rect 3368 3782 3414 3834
rect 3118 3780 3174 3782
rect 3198 3780 3254 3782
rect 3278 3780 3334 3782
rect 3358 3780 3414 3782
rect 1761 3290 1817 3292
rect 1841 3290 1897 3292
rect 1921 3290 1977 3292
rect 2001 3290 2057 3292
rect 1761 3238 1807 3290
rect 1807 3238 1817 3290
rect 1841 3238 1871 3290
rect 1871 3238 1883 3290
rect 1883 3238 1897 3290
rect 1921 3238 1935 3290
rect 1935 3238 1947 3290
rect 1947 3238 1977 3290
rect 2001 3238 2011 3290
rect 2011 3238 2057 3290
rect 1761 3236 1817 3238
rect 1841 3236 1897 3238
rect 1921 3236 1977 3238
rect 2001 3236 2057 3238
rect 3118 2746 3174 2748
rect 3198 2746 3254 2748
rect 3278 2746 3334 2748
rect 3358 2746 3414 2748
rect 3118 2694 3164 2746
rect 3164 2694 3174 2746
rect 3198 2694 3228 2746
rect 3228 2694 3240 2746
rect 3240 2694 3254 2746
rect 3278 2694 3292 2746
rect 3292 2694 3304 2746
rect 3304 2694 3334 2746
rect 3358 2694 3368 2746
rect 3368 2694 3414 2746
rect 3118 2692 3174 2694
rect 3198 2692 3254 2694
rect 3278 2692 3334 2694
rect 3358 2692 3414 2694
rect 1761 2202 1817 2204
rect 1841 2202 1897 2204
rect 1921 2202 1977 2204
rect 2001 2202 2057 2204
rect 1761 2150 1807 2202
rect 1807 2150 1817 2202
rect 1841 2150 1871 2202
rect 1871 2150 1883 2202
rect 1883 2150 1897 2202
rect 1921 2150 1935 2202
rect 1935 2150 1947 2202
rect 1947 2150 1977 2202
rect 2001 2150 2011 2202
rect 2011 2150 2057 2202
rect 1761 2148 1817 2150
rect 1841 2148 1897 2150
rect 1921 2148 1977 2150
rect 2001 2148 2057 2150
rect 4475 6554 4531 6556
rect 4555 6554 4611 6556
rect 4635 6554 4691 6556
rect 4715 6554 4771 6556
rect 4475 6502 4521 6554
rect 4521 6502 4531 6554
rect 4555 6502 4585 6554
rect 4585 6502 4597 6554
rect 4597 6502 4611 6554
rect 4635 6502 4649 6554
rect 4649 6502 4661 6554
rect 4661 6502 4691 6554
rect 4715 6502 4725 6554
rect 4725 6502 4771 6554
rect 4475 6500 4531 6502
rect 4555 6500 4611 6502
rect 4635 6500 4691 6502
rect 4715 6500 4771 6502
rect 4475 5466 4531 5468
rect 4555 5466 4611 5468
rect 4635 5466 4691 5468
rect 4715 5466 4771 5468
rect 4475 5414 4521 5466
rect 4521 5414 4531 5466
rect 4555 5414 4585 5466
rect 4585 5414 4597 5466
rect 4597 5414 4611 5466
rect 4635 5414 4649 5466
rect 4649 5414 4661 5466
rect 4661 5414 4691 5466
rect 4715 5414 4725 5466
rect 4725 5414 4771 5466
rect 4475 5412 4531 5414
rect 4555 5412 4611 5414
rect 4635 5412 4691 5414
rect 4715 5412 4771 5414
rect 4475 4378 4531 4380
rect 4555 4378 4611 4380
rect 4635 4378 4691 4380
rect 4715 4378 4771 4380
rect 4475 4326 4521 4378
rect 4521 4326 4531 4378
rect 4555 4326 4585 4378
rect 4585 4326 4597 4378
rect 4597 4326 4611 4378
rect 4635 4326 4649 4378
rect 4649 4326 4661 4378
rect 4661 4326 4691 4378
rect 4715 4326 4725 4378
rect 4725 4326 4771 4378
rect 4475 4324 4531 4326
rect 4555 4324 4611 4326
rect 4635 4324 4691 4326
rect 4715 4324 4771 4326
rect 4475 3290 4531 3292
rect 4555 3290 4611 3292
rect 4635 3290 4691 3292
rect 4715 3290 4771 3292
rect 4475 3238 4521 3290
rect 4521 3238 4531 3290
rect 4555 3238 4585 3290
rect 4585 3238 4597 3290
rect 4597 3238 4611 3290
rect 4635 3238 4649 3290
rect 4649 3238 4661 3290
rect 4661 3238 4691 3290
rect 4715 3238 4725 3290
rect 4725 3238 4771 3290
rect 4475 3236 4531 3238
rect 4555 3236 4611 3238
rect 4635 3236 4691 3238
rect 4715 3236 4771 3238
rect 5832 7098 5888 7100
rect 5912 7098 5968 7100
rect 5992 7098 6048 7100
rect 6072 7098 6128 7100
rect 5832 7046 5878 7098
rect 5878 7046 5888 7098
rect 5912 7046 5942 7098
rect 5942 7046 5954 7098
rect 5954 7046 5968 7098
rect 5992 7046 6006 7098
rect 6006 7046 6018 7098
rect 6018 7046 6048 7098
rect 6072 7046 6082 7098
rect 6082 7046 6128 7098
rect 5832 7044 5888 7046
rect 5912 7044 5968 7046
rect 5992 7044 6048 7046
rect 6072 7044 6128 7046
rect 8546 7098 8602 7100
rect 8626 7098 8682 7100
rect 8706 7098 8762 7100
rect 8786 7098 8842 7100
rect 8546 7046 8592 7098
rect 8592 7046 8602 7098
rect 8626 7046 8656 7098
rect 8656 7046 8668 7098
rect 8668 7046 8682 7098
rect 8706 7046 8720 7098
rect 8720 7046 8732 7098
rect 8732 7046 8762 7098
rect 8786 7046 8796 7098
rect 8796 7046 8842 7098
rect 8546 7044 8602 7046
rect 8626 7044 8682 7046
rect 8706 7044 8762 7046
rect 8786 7044 8842 7046
rect 11260 7098 11316 7100
rect 11340 7098 11396 7100
rect 11420 7098 11476 7100
rect 11500 7098 11556 7100
rect 11260 7046 11306 7098
rect 11306 7046 11316 7098
rect 11340 7046 11370 7098
rect 11370 7046 11382 7098
rect 11382 7046 11396 7098
rect 11420 7046 11434 7098
rect 11434 7046 11446 7098
rect 11446 7046 11476 7098
rect 11500 7046 11510 7098
rect 11510 7046 11556 7098
rect 11260 7044 11316 7046
rect 11340 7044 11396 7046
rect 11420 7044 11476 7046
rect 11500 7044 11556 7046
rect 7189 6554 7245 6556
rect 7269 6554 7325 6556
rect 7349 6554 7405 6556
rect 7429 6554 7485 6556
rect 7189 6502 7235 6554
rect 7235 6502 7245 6554
rect 7269 6502 7299 6554
rect 7299 6502 7311 6554
rect 7311 6502 7325 6554
rect 7349 6502 7363 6554
rect 7363 6502 7375 6554
rect 7375 6502 7405 6554
rect 7429 6502 7439 6554
rect 7439 6502 7485 6554
rect 7189 6500 7245 6502
rect 7269 6500 7325 6502
rect 7349 6500 7405 6502
rect 7429 6500 7485 6502
rect 9903 6554 9959 6556
rect 9983 6554 10039 6556
rect 10063 6554 10119 6556
rect 10143 6554 10199 6556
rect 9903 6502 9949 6554
rect 9949 6502 9959 6554
rect 9983 6502 10013 6554
rect 10013 6502 10025 6554
rect 10025 6502 10039 6554
rect 10063 6502 10077 6554
rect 10077 6502 10089 6554
rect 10089 6502 10119 6554
rect 10143 6502 10153 6554
rect 10153 6502 10199 6554
rect 9903 6500 9959 6502
rect 9983 6500 10039 6502
rect 10063 6500 10119 6502
rect 10143 6500 10199 6502
rect 5832 6010 5888 6012
rect 5912 6010 5968 6012
rect 5992 6010 6048 6012
rect 6072 6010 6128 6012
rect 5832 5958 5878 6010
rect 5878 5958 5888 6010
rect 5912 5958 5942 6010
rect 5942 5958 5954 6010
rect 5954 5958 5968 6010
rect 5992 5958 6006 6010
rect 6006 5958 6018 6010
rect 6018 5958 6048 6010
rect 6072 5958 6082 6010
rect 6082 5958 6128 6010
rect 5832 5956 5888 5958
rect 5912 5956 5968 5958
rect 5992 5956 6048 5958
rect 6072 5956 6128 5958
rect 8546 6010 8602 6012
rect 8626 6010 8682 6012
rect 8706 6010 8762 6012
rect 8786 6010 8842 6012
rect 8546 5958 8592 6010
rect 8592 5958 8602 6010
rect 8626 5958 8656 6010
rect 8656 5958 8668 6010
rect 8668 5958 8682 6010
rect 8706 5958 8720 6010
rect 8720 5958 8732 6010
rect 8732 5958 8762 6010
rect 8786 5958 8796 6010
rect 8796 5958 8842 6010
rect 8546 5956 8602 5958
rect 8626 5956 8682 5958
rect 8706 5956 8762 5958
rect 8786 5956 8842 5958
rect 11260 6010 11316 6012
rect 11340 6010 11396 6012
rect 11420 6010 11476 6012
rect 11500 6010 11556 6012
rect 11260 5958 11306 6010
rect 11306 5958 11316 6010
rect 11340 5958 11370 6010
rect 11370 5958 11382 6010
rect 11382 5958 11396 6010
rect 11420 5958 11434 6010
rect 11434 5958 11446 6010
rect 11446 5958 11476 6010
rect 11500 5958 11510 6010
rect 11510 5958 11556 6010
rect 11260 5956 11316 5958
rect 11340 5956 11396 5958
rect 11420 5956 11476 5958
rect 11500 5956 11556 5958
rect 7189 5466 7245 5468
rect 7269 5466 7325 5468
rect 7349 5466 7405 5468
rect 7429 5466 7485 5468
rect 7189 5414 7235 5466
rect 7235 5414 7245 5466
rect 7269 5414 7299 5466
rect 7299 5414 7311 5466
rect 7311 5414 7325 5466
rect 7349 5414 7363 5466
rect 7363 5414 7375 5466
rect 7375 5414 7405 5466
rect 7429 5414 7439 5466
rect 7439 5414 7485 5466
rect 7189 5412 7245 5414
rect 7269 5412 7325 5414
rect 7349 5412 7405 5414
rect 7429 5412 7485 5414
rect 9903 5466 9959 5468
rect 9983 5466 10039 5468
rect 10063 5466 10119 5468
rect 10143 5466 10199 5468
rect 9903 5414 9949 5466
rect 9949 5414 9959 5466
rect 9983 5414 10013 5466
rect 10013 5414 10025 5466
rect 10025 5414 10039 5466
rect 10063 5414 10077 5466
rect 10077 5414 10089 5466
rect 10089 5414 10119 5466
rect 10143 5414 10153 5466
rect 10153 5414 10199 5466
rect 9903 5412 9959 5414
rect 9983 5412 10039 5414
rect 10063 5412 10119 5414
rect 10143 5412 10199 5414
rect 5832 4922 5888 4924
rect 5912 4922 5968 4924
rect 5992 4922 6048 4924
rect 6072 4922 6128 4924
rect 5832 4870 5878 4922
rect 5878 4870 5888 4922
rect 5912 4870 5942 4922
rect 5942 4870 5954 4922
rect 5954 4870 5968 4922
rect 5992 4870 6006 4922
rect 6006 4870 6018 4922
rect 6018 4870 6048 4922
rect 6072 4870 6082 4922
rect 6082 4870 6128 4922
rect 5832 4868 5888 4870
rect 5912 4868 5968 4870
rect 5992 4868 6048 4870
rect 6072 4868 6128 4870
rect 8546 4922 8602 4924
rect 8626 4922 8682 4924
rect 8706 4922 8762 4924
rect 8786 4922 8842 4924
rect 8546 4870 8592 4922
rect 8592 4870 8602 4922
rect 8626 4870 8656 4922
rect 8656 4870 8668 4922
rect 8668 4870 8682 4922
rect 8706 4870 8720 4922
rect 8720 4870 8732 4922
rect 8732 4870 8762 4922
rect 8786 4870 8796 4922
rect 8796 4870 8842 4922
rect 8546 4868 8602 4870
rect 8626 4868 8682 4870
rect 8706 4868 8762 4870
rect 8786 4868 8842 4870
rect 11260 4922 11316 4924
rect 11340 4922 11396 4924
rect 11420 4922 11476 4924
rect 11500 4922 11556 4924
rect 11260 4870 11306 4922
rect 11306 4870 11316 4922
rect 11340 4870 11370 4922
rect 11370 4870 11382 4922
rect 11382 4870 11396 4922
rect 11420 4870 11434 4922
rect 11434 4870 11446 4922
rect 11446 4870 11476 4922
rect 11500 4870 11510 4922
rect 11510 4870 11556 4922
rect 11260 4868 11316 4870
rect 11340 4868 11396 4870
rect 11420 4868 11476 4870
rect 11500 4868 11556 4870
rect 7189 4378 7245 4380
rect 7269 4378 7325 4380
rect 7349 4378 7405 4380
rect 7429 4378 7485 4380
rect 7189 4326 7235 4378
rect 7235 4326 7245 4378
rect 7269 4326 7299 4378
rect 7299 4326 7311 4378
rect 7311 4326 7325 4378
rect 7349 4326 7363 4378
rect 7363 4326 7375 4378
rect 7375 4326 7405 4378
rect 7429 4326 7439 4378
rect 7439 4326 7485 4378
rect 7189 4324 7245 4326
rect 7269 4324 7325 4326
rect 7349 4324 7405 4326
rect 7429 4324 7485 4326
rect 9903 4378 9959 4380
rect 9983 4378 10039 4380
rect 10063 4378 10119 4380
rect 10143 4378 10199 4380
rect 9903 4326 9949 4378
rect 9949 4326 9959 4378
rect 9983 4326 10013 4378
rect 10013 4326 10025 4378
rect 10025 4326 10039 4378
rect 10063 4326 10077 4378
rect 10077 4326 10089 4378
rect 10089 4326 10119 4378
rect 10143 4326 10153 4378
rect 10153 4326 10199 4378
rect 9903 4324 9959 4326
rect 9983 4324 10039 4326
rect 10063 4324 10119 4326
rect 10143 4324 10199 4326
rect 5832 3834 5888 3836
rect 5912 3834 5968 3836
rect 5992 3834 6048 3836
rect 6072 3834 6128 3836
rect 5832 3782 5878 3834
rect 5878 3782 5888 3834
rect 5912 3782 5942 3834
rect 5942 3782 5954 3834
rect 5954 3782 5968 3834
rect 5992 3782 6006 3834
rect 6006 3782 6018 3834
rect 6018 3782 6048 3834
rect 6072 3782 6082 3834
rect 6082 3782 6128 3834
rect 5832 3780 5888 3782
rect 5912 3780 5968 3782
rect 5992 3780 6048 3782
rect 6072 3780 6128 3782
rect 8546 3834 8602 3836
rect 8626 3834 8682 3836
rect 8706 3834 8762 3836
rect 8786 3834 8842 3836
rect 8546 3782 8592 3834
rect 8592 3782 8602 3834
rect 8626 3782 8656 3834
rect 8656 3782 8668 3834
rect 8668 3782 8682 3834
rect 8706 3782 8720 3834
rect 8720 3782 8732 3834
rect 8732 3782 8762 3834
rect 8786 3782 8796 3834
rect 8796 3782 8842 3834
rect 8546 3780 8602 3782
rect 8626 3780 8682 3782
rect 8706 3780 8762 3782
rect 8786 3780 8842 3782
rect 11260 3834 11316 3836
rect 11340 3834 11396 3836
rect 11420 3834 11476 3836
rect 11500 3834 11556 3836
rect 11260 3782 11306 3834
rect 11306 3782 11316 3834
rect 11340 3782 11370 3834
rect 11370 3782 11382 3834
rect 11382 3782 11396 3834
rect 11420 3782 11434 3834
rect 11434 3782 11446 3834
rect 11446 3782 11476 3834
rect 11500 3782 11510 3834
rect 11510 3782 11556 3834
rect 11260 3780 11316 3782
rect 11340 3780 11396 3782
rect 11420 3780 11476 3782
rect 11500 3780 11556 3782
rect 4066 2508 4122 2544
rect 4066 2488 4068 2508
rect 4068 2488 4120 2508
rect 4120 2488 4122 2508
rect 3118 1658 3174 1660
rect 3198 1658 3254 1660
rect 3278 1658 3334 1660
rect 3358 1658 3414 1660
rect 3118 1606 3164 1658
rect 3164 1606 3174 1658
rect 3198 1606 3228 1658
rect 3228 1606 3240 1658
rect 3240 1606 3254 1658
rect 3278 1606 3292 1658
rect 3292 1606 3304 1658
rect 3304 1606 3334 1658
rect 3358 1606 3368 1658
rect 3368 1606 3414 1658
rect 3118 1604 3174 1606
rect 3198 1604 3254 1606
rect 3278 1604 3334 1606
rect 3358 1604 3414 1606
rect 1761 1114 1817 1116
rect 1841 1114 1897 1116
rect 1921 1114 1977 1116
rect 2001 1114 2057 1116
rect 1761 1062 1807 1114
rect 1807 1062 1817 1114
rect 1841 1062 1871 1114
rect 1871 1062 1883 1114
rect 1883 1062 1897 1114
rect 1921 1062 1935 1114
rect 1935 1062 1947 1114
rect 1947 1062 1977 1114
rect 2001 1062 2011 1114
rect 2011 1062 2057 1114
rect 1761 1060 1817 1062
rect 1841 1060 1897 1062
rect 1921 1060 1977 1062
rect 2001 1060 2057 1062
rect 5832 2746 5888 2748
rect 5912 2746 5968 2748
rect 5992 2746 6048 2748
rect 6072 2746 6128 2748
rect 5832 2694 5878 2746
rect 5878 2694 5888 2746
rect 5912 2694 5942 2746
rect 5942 2694 5954 2746
rect 5954 2694 5968 2746
rect 5992 2694 6006 2746
rect 6006 2694 6018 2746
rect 6018 2694 6048 2746
rect 6072 2694 6082 2746
rect 6082 2694 6128 2746
rect 5832 2692 5888 2694
rect 5912 2692 5968 2694
rect 5992 2692 6048 2694
rect 6072 2692 6128 2694
rect 5538 2508 5594 2544
rect 5538 2488 5540 2508
rect 5540 2488 5592 2508
rect 5592 2488 5594 2508
rect 4475 2202 4531 2204
rect 4555 2202 4611 2204
rect 4635 2202 4691 2204
rect 4715 2202 4771 2204
rect 4475 2150 4521 2202
rect 4521 2150 4531 2202
rect 4555 2150 4585 2202
rect 4585 2150 4597 2202
rect 4597 2150 4611 2202
rect 4635 2150 4649 2202
rect 4649 2150 4661 2202
rect 4661 2150 4691 2202
rect 4715 2150 4725 2202
rect 4725 2150 4771 2202
rect 4475 2148 4531 2150
rect 4555 2148 4611 2150
rect 4635 2148 4691 2150
rect 4715 2148 4771 2150
rect 11242 3476 11244 3496
rect 11244 3476 11296 3496
rect 11296 3476 11298 3496
rect 7189 3290 7245 3292
rect 7269 3290 7325 3292
rect 7349 3290 7405 3292
rect 7429 3290 7485 3292
rect 7189 3238 7235 3290
rect 7235 3238 7245 3290
rect 7269 3238 7299 3290
rect 7299 3238 7311 3290
rect 7311 3238 7325 3290
rect 7349 3238 7363 3290
rect 7363 3238 7375 3290
rect 7375 3238 7405 3290
rect 7429 3238 7439 3290
rect 7439 3238 7485 3290
rect 7189 3236 7245 3238
rect 7269 3236 7325 3238
rect 7349 3236 7405 3238
rect 7429 3236 7485 3238
rect 5832 1658 5888 1660
rect 5912 1658 5968 1660
rect 5992 1658 6048 1660
rect 6072 1658 6128 1660
rect 5832 1606 5878 1658
rect 5878 1606 5888 1658
rect 5912 1606 5942 1658
rect 5942 1606 5954 1658
rect 5954 1606 5968 1658
rect 5992 1606 6006 1658
rect 6006 1606 6018 1658
rect 6018 1606 6048 1658
rect 6072 1606 6082 1658
rect 6082 1606 6128 1658
rect 5832 1604 5888 1606
rect 5912 1604 5968 1606
rect 5992 1604 6048 1606
rect 6072 1604 6128 1606
rect 4475 1114 4531 1116
rect 4555 1114 4611 1116
rect 4635 1114 4691 1116
rect 4715 1114 4771 1116
rect 4475 1062 4521 1114
rect 4521 1062 4531 1114
rect 4555 1062 4585 1114
rect 4585 1062 4597 1114
rect 4597 1062 4611 1114
rect 4635 1062 4649 1114
rect 4649 1062 4661 1114
rect 4661 1062 4691 1114
rect 4715 1062 4725 1114
rect 4725 1062 4771 1114
rect 4475 1060 4531 1062
rect 4555 1060 4611 1062
rect 4635 1060 4691 1062
rect 4715 1060 4771 1062
rect 8546 2746 8602 2748
rect 8626 2746 8682 2748
rect 8706 2746 8762 2748
rect 8786 2746 8842 2748
rect 8546 2694 8592 2746
rect 8592 2694 8602 2746
rect 8626 2694 8656 2746
rect 8656 2694 8668 2746
rect 8668 2694 8682 2746
rect 8706 2694 8720 2746
rect 8720 2694 8732 2746
rect 8732 2694 8762 2746
rect 8786 2694 8796 2746
rect 8796 2694 8842 2746
rect 8546 2692 8602 2694
rect 8626 2692 8682 2694
rect 8706 2692 8762 2694
rect 8786 2692 8842 2694
rect 11242 3440 11298 3476
rect 9903 3290 9959 3292
rect 9983 3290 10039 3292
rect 10063 3290 10119 3292
rect 10143 3290 10199 3292
rect 9903 3238 9949 3290
rect 9949 3238 9959 3290
rect 9983 3238 10013 3290
rect 10013 3238 10025 3290
rect 10025 3238 10039 3290
rect 10063 3238 10077 3290
rect 10077 3238 10089 3290
rect 10089 3238 10119 3290
rect 10143 3238 10153 3290
rect 10153 3238 10199 3290
rect 9903 3236 9959 3238
rect 9983 3236 10039 3238
rect 10063 3236 10119 3238
rect 10143 3236 10199 3238
rect 11260 2746 11316 2748
rect 11340 2746 11396 2748
rect 11420 2746 11476 2748
rect 11500 2746 11556 2748
rect 11260 2694 11306 2746
rect 11306 2694 11316 2746
rect 11340 2694 11370 2746
rect 11370 2694 11382 2746
rect 11382 2694 11396 2746
rect 11420 2694 11434 2746
rect 11434 2694 11446 2746
rect 11446 2694 11476 2746
rect 11500 2694 11510 2746
rect 11510 2694 11556 2746
rect 11260 2692 11316 2694
rect 11340 2692 11396 2694
rect 11420 2692 11476 2694
rect 11500 2692 11556 2694
rect 7189 2202 7245 2204
rect 7269 2202 7325 2204
rect 7349 2202 7405 2204
rect 7429 2202 7485 2204
rect 7189 2150 7235 2202
rect 7235 2150 7245 2202
rect 7269 2150 7299 2202
rect 7299 2150 7311 2202
rect 7311 2150 7325 2202
rect 7349 2150 7363 2202
rect 7363 2150 7375 2202
rect 7375 2150 7405 2202
rect 7429 2150 7439 2202
rect 7439 2150 7485 2202
rect 7189 2148 7245 2150
rect 7269 2148 7325 2150
rect 7349 2148 7405 2150
rect 7429 2148 7485 2150
rect 8546 1658 8602 1660
rect 8626 1658 8682 1660
rect 8706 1658 8762 1660
rect 8786 1658 8842 1660
rect 8546 1606 8592 1658
rect 8592 1606 8602 1658
rect 8626 1606 8656 1658
rect 8656 1606 8668 1658
rect 8668 1606 8682 1658
rect 8706 1606 8720 1658
rect 8720 1606 8732 1658
rect 8732 1606 8762 1658
rect 8786 1606 8796 1658
rect 8796 1606 8842 1658
rect 8546 1604 8602 1606
rect 8626 1604 8682 1606
rect 8706 1604 8762 1606
rect 8786 1604 8842 1606
rect 9903 2202 9959 2204
rect 9983 2202 10039 2204
rect 10063 2202 10119 2204
rect 10143 2202 10199 2204
rect 9903 2150 9949 2202
rect 9949 2150 9959 2202
rect 9983 2150 10013 2202
rect 10013 2150 10025 2202
rect 10025 2150 10039 2202
rect 10063 2150 10077 2202
rect 10077 2150 10089 2202
rect 10089 2150 10119 2202
rect 10143 2150 10153 2202
rect 10153 2150 10199 2202
rect 9903 2148 9959 2150
rect 9983 2148 10039 2150
rect 10063 2148 10119 2150
rect 10143 2148 10199 2150
rect 11260 1658 11316 1660
rect 11340 1658 11396 1660
rect 11420 1658 11476 1660
rect 11500 1658 11556 1660
rect 11260 1606 11306 1658
rect 11306 1606 11316 1658
rect 11340 1606 11370 1658
rect 11370 1606 11382 1658
rect 11382 1606 11396 1658
rect 11420 1606 11434 1658
rect 11434 1606 11446 1658
rect 11446 1606 11476 1658
rect 11500 1606 11510 1658
rect 11510 1606 11556 1658
rect 11260 1604 11316 1606
rect 11340 1604 11396 1606
rect 11420 1604 11476 1606
rect 11500 1604 11556 1606
rect 7189 1114 7245 1116
rect 7269 1114 7325 1116
rect 7349 1114 7405 1116
rect 7429 1114 7485 1116
rect 7189 1062 7235 1114
rect 7235 1062 7245 1114
rect 7269 1062 7299 1114
rect 7299 1062 7311 1114
rect 7311 1062 7325 1114
rect 7349 1062 7363 1114
rect 7363 1062 7375 1114
rect 7375 1062 7405 1114
rect 7429 1062 7439 1114
rect 7439 1062 7485 1114
rect 7189 1060 7245 1062
rect 7269 1060 7325 1062
rect 7349 1060 7405 1062
rect 7429 1060 7485 1062
rect 9903 1114 9959 1116
rect 9983 1114 10039 1116
rect 10063 1114 10119 1116
rect 10143 1114 10199 1116
rect 9903 1062 9949 1114
rect 9949 1062 9959 1114
rect 9983 1062 10013 1114
rect 10013 1062 10025 1114
rect 10025 1062 10039 1114
rect 10063 1062 10077 1114
rect 10077 1062 10089 1114
rect 10089 1062 10119 1114
rect 10143 1062 10153 1114
rect 10153 1062 10199 1114
rect 9903 1060 9959 1062
rect 9983 1060 10039 1062
rect 10063 1060 10119 1062
rect 10143 1060 10199 1062
rect 3118 570 3174 572
rect 3198 570 3254 572
rect 3278 570 3334 572
rect 3358 570 3414 572
rect 3118 518 3164 570
rect 3164 518 3174 570
rect 3198 518 3228 570
rect 3228 518 3240 570
rect 3240 518 3254 570
rect 3278 518 3292 570
rect 3292 518 3304 570
rect 3304 518 3334 570
rect 3358 518 3368 570
rect 3368 518 3414 570
rect 3118 516 3174 518
rect 3198 516 3254 518
rect 3278 516 3334 518
rect 3358 516 3414 518
rect 5832 570 5888 572
rect 5912 570 5968 572
rect 5992 570 6048 572
rect 6072 570 6128 572
rect 5832 518 5878 570
rect 5878 518 5888 570
rect 5912 518 5942 570
rect 5942 518 5954 570
rect 5954 518 5968 570
rect 5992 518 6006 570
rect 6006 518 6018 570
rect 6018 518 6048 570
rect 6072 518 6082 570
rect 6082 518 6128 570
rect 5832 516 5888 518
rect 5912 516 5968 518
rect 5992 516 6048 518
rect 6072 516 6128 518
rect 8546 570 8602 572
rect 8626 570 8682 572
rect 8706 570 8762 572
rect 8786 570 8842 572
rect 8546 518 8592 570
rect 8592 518 8602 570
rect 8626 518 8656 570
rect 8656 518 8668 570
rect 8668 518 8682 570
rect 8706 518 8720 570
rect 8720 518 8732 570
rect 8732 518 8762 570
rect 8786 518 8796 570
rect 8796 518 8842 570
rect 8546 516 8602 518
rect 8626 516 8682 518
rect 8706 516 8762 518
rect 8786 516 8842 518
rect 11260 570 11316 572
rect 11340 570 11396 572
rect 11420 570 11476 572
rect 11500 570 11556 572
rect 11260 518 11306 570
rect 11306 518 11316 570
rect 11340 518 11370 570
rect 11370 518 11382 570
rect 11382 518 11396 570
rect 11420 518 11434 570
rect 11434 518 11446 570
rect 11446 518 11476 570
rect 11500 518 11510 570
rect 11510 518 11556 570
rect 11260 516 11316 518
rect 11340 516 11396 518
rect 11420 516 11476 518
rect 11500 516 11556 518
<< metal3 >>
rect 3108 11456 3424 11457
rect 3108 11392 3114 11456
rect 3178 11392 3194 11456
rect 3258 11392 3274 11456
rect 3338 11392 3354 11456
rect 3418 11392 3424 11456
rect 3108 11391 3424 11392
rect 5822 11456 6138 11457
rect 5822 11392 5828 11456
rect 5892 11392 5908 11456
rect 5972 11392 5988 11456
rect 6052 11392 6068 11456
rect 6132 11392 6138 11456
rect 5822 11391 6138 11392
rect 8536 11456 8852 11457
rect 8536 11392 8542 11456
rect 8606 11392 8622 11456
rect 8686 11392 8702 11456
rect 8766 11392 8782 11456
rect 8846 11392 8852 11456
rect 8536 11391 8852 11392
rect 11250 11456 11566 11457
rect 11250 11392 11256 11456
rect 11320 11392 11336 11456
rect 11400 11392 11416 11456
rect 11480 11392 11496 11456
rect 11560 11392 11566 11456
rect 11250 11391 11566 11392
rect 1751 10912 2067 10913
rect 1751 10848 1757 10912
rect 1821 10848 1837 10912
rect 1901 10848 1917 10912
rect 1981 10848 1997 10912
rect 2061 10848 2067 10912
rect 1751 10847 2067 10848
rect 4465 10912 4781 10913
rect 4465 10848 4471 10912
rect 4535 10848 4551 10912
rect 4615 10848 4631 10912
rect 4695 10848 4711 10912
rect 4775 10848 4781 10912
rect 4465 10847 4781 10848
rect 7179 10912 7495 10913
rect 7179 10848 7185 10912
rect 7249 10848 7265 10912
rect 7329 10848 7345 10912
rect 7409 10848 7425 10912
rect 7489 10848 7495 10912
rect 7179 10847 7495 10848
rect 9893 10912 10209 10913
rect 9893 10848 9899 10912
rect 9963 10848 9979 10912
rect 10043 10848 10059 10912
rect 10123 10848 10139 10912
rect 10203 10848 10209 10912
rect 9893 10847 10209 10848
rect 3108 10368 3424 10369
rect 3108 10304 3114 10368
rect 3178 10304 3194 10368
rect 3258 10304 3274 10368
rect 3338 10304 3354 10368
rect 3418 10304 3424 10368
rect 3108 10303 3424 10304
rect 5822 10368 6138 10369
rect 5822 10304 5828 10368
rect 5892 10304 5908 10368
rect 5972 10304 5988 10368
rect 6052 10304 6068 10368
rect 6132 10304 6138 10368
rect 5822 10303 6138 10304
rect 8536 10368 8852 10369
rect 8536 10304 8542 10368
rect 8606 10304 8622 10368
rect 8686 10304 8702 10368
rect 8766 10304 8782 10368
rect 8846 10304 8852 10368
rect 8536 10303 8852 10304
rect 11250 10368 11566 10369
rect 11250 10304 11256 10368
rect 11320 10304 11336 10368
rect 11400 10304 11416 10368
rect 11480 10304 11496 10368
rect 11560 10304 11566 10368
rect 11250 10303 11566 10304
rect 1751 9824 2067 9825
rect 1751 9760 1757 9824
rect 1821 9760 1837 9824
rect 1901 9760 1917 9824
rect 1981 9760 1997 9824
rect 2061 9760 2067 9824
rect 1751 9759 2067 9760
rect 4465 9824 4781 9825
rect 4465 9760 4471 9824
rect 4535 9760 4551 9824
rect 4615 9760 4631 9824
rect 4695 9760 4711 9824
rect 4775 9760 4781 9824
rect 4465 9759 4781 9760
rect 7179 9824 7495 9825
rect 7179 9760 7185 9824
rect 7249 9760 7265 9824
rect 7329 9760 7345 9824
rect 7409 9760 7425 9824
rect 7489 9760 7495 9824
rect 7179 9759 7495 9760
rect 9893 9824 10209 9825
rect 9893 9760 9899 9824
rect 9963 9760 9979 9824
rect 10043 9760 10059 9824
rect 10123 9760 10139 9824
rect 10203 9760 10209 9824
rect 9893 9759 10209 9760
rect 3108 9280 3424 9281
rect 3108 9216 3114 9280
rect 3178 9216 3194 9280
rect 3258 9216 3274 9280
rect 3338 9216 3354 9280
rect 3418 9216 3424 9280
rect 3108 9215 3424 9216
rect 5822 9280 6138 9281
rect 5822 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5988 9280
rect 6052 9216 6068 9280
rect 6132 9216 6138 9280
rect 5822 9215 6138 9216
rect 8536 9280 8852 9281
rect 8536 9216 8542 9280
rect 8606 9216 8622 9280
rect 8686 9216 8702 9280
rect 8766 9216 8782 9280
rect 8846 9216 8852 9280
rect 8536 9215 8852 9216
rect 11250 9280 11566 9281
rect 11250 9216 11256 9280
rect 11320 9216 11336 9280
rect 11400 9216 11416 9280
rect 11480 9216 11496 9280
rect 11560 9216 11566 9280
rect 11250 9215 11566 9216
rect 1751 8736 2067 8737
rect 1751 8672 1757 8736
rect 1821 8672 1837 8736
rect 1901 8672 1917 8736
rect 1981 8672 1997 8736
rect 2061 8672 2067 8736
rect 1751 8671 2067 8672
rect 4465 8736 4781 8737
rect 4465 8672 4471 8736
rect 4535 8672 4551 8736
rect 4615 8672 4631 8736
rect 4695 8672 4711 8736
rect 4775 8672 4781 8736
rect 4465 8671 4781 8672
rect 7179 8736 7495 8737
rect 7179 8672 7185 8736
rect 7249 8672 7265 8736
rect 7329 8672 7345 8736
rect 7409 8672 7425 8736
rect 7489 8672 7495 8736
rect 7179 8671 7495 8672
rect 9893 8736 10209 8737
rect 9893 8672 9899 8736
rect 9963 8672 9979 8736
rect 10043 8672 10059 8736
rect 10123 8672 10139 8736
rect 10203 8672 10209 8736
rect 9893 8671 10209 8672
rect 0 8258 400 8288
rect 2773 8258 2839 8261
rect 0 8256 2839 8258
rect 0 8200 2778 8256
rect 2834 8200 2839 8256
rect 0 8198 2839 8200
rect 0 8168 400 8198
rect 2773 8195 2839 8198
rect 3108 8192 3424 8193
rect 3108 8128 3114 8192
rect 3178 8128 3194 8192
rect 3258 8128 3274 8192
rect 3338 8128 3354 8192
rect 3418 8128 3424 8192
rect 3108 8127 3424 8128
rect 5822 8192 6138 8193
rect 5822 8128 5828 8192
rect 5892 8128 5908 8192
rect 5972 8128 5988 8192
rect 6052 8128 6068 8192
rect 6132 8128 6138 8192
rect 5822 8127 6138 8128
rect 8536 8192 8852 8193
rect 8536 8128 8542 8192
rect 8606 8128 8622 8192
rect 8686 8128 8702 8192
rect 8766 8128 8782 8192
rect 8846 8128 8852 8192
rect 8536 8127 8852 8128
rect 11250 8192 11566 8193
rect 11250 8128 11256 8192
rect 11320 8128 11336 8192
rect 11400 8128 11416 8192
rect 11480 8128 11496 8192
rect 11560 8128 11566 8192
rect 11250 8127 11566 8128
rect 1751 7648 2067 7649
rect 1751 7584 1757 7648
rect 1821 7584 1837 7648
rect 1901 7584 1917 7648
rect 1981 7584 1997 7648
rect 2061 7584 2067 7648
rect 1751 7583 2067 7584
rect 4465 7648 4781 7649
rect 4465 7584 4471 7648
rect 4535 7584 4551 7648
rect 4615 7584 4631 7648
rect 4695 7584 4711 7648
rect 4775 7584 4781 7648
rect 4465 7583 4781 7584
rect 7179 7648 7495 7649
rect 7179 7584 7185 7648
rect 7249 7584 7265 7648
rect 7329 7584 7345 7648
rect 7409 7584 7425 7648
rect 7489 7584 7495 7648
rect 7179 7583 7495 7584
rect 9893 7648 10209 7649
rect 9893 7584 9899 7648
rect 9963 7584 9979 7648
rect 10043 7584 10059 7648
rect 10123 7584 10139 7648
rect 10203 7584 10209 7648
rect 9893 7583 10209 7584
rect 3108 7104 3424 7105
rect 3108 7040 3114 7104
rect 3178 7040 3194 7104
rect 3258 7040 3274 7104
rect 3338 7040 3354 7104
rect 3418 7040 3424 7104
rect 3108 7039 3424 7040
rect 5822 7104 6138 7105
rect 5822 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5988 7104
rect 6052 7040 6068 7104
rect 6132 7040 6138 7104
rect 5822 7039 6138 7040
rect 8536 7104 8852 7105
rect 8536 7040 8542 7104
rect 8606 7040 8622 7104
rect 8686 7040 8702 7104
rect 8766 7040 8782 7104
rect 8846 7040 8852 7104
rect 8536 7039 8852 7040
rect 11250 7104 11566 7105
rect 11250 7040 11256 7104
rect 11320 7040 11336 7104
rect 11400 7040 11416 7104
rect 11480 7040 11496 7104
rect 11560 7040 11566 7104
rect 11250 7039 11566 7040
rect 1751 6560 2067 6561
rect 1751 6496 1757 6560
rect 1821 6496 1837 6560
rect 1901 6496 1917 6560
rect 1981 6496 1997 6560
rect 2061 6496 2067 6560
rect 1751 6495 2067 6496
rect 4465 6560 4781 6561
rect 4465 6496 4471 6560
rect 4535 6496 4551 6560
rect 4615 6496 4631 6560
rect 4695 6496 4711 6560
rect 4775 6496 4781 6560
rect 4465 6495 4781 6496
rect 7179 6560 7495 6561
rect 7179 6496 7185 6560
rect 7249 6496 7265 6560
rect 7329 6496 7345 6560
rect 7409 6496 7425 6560
rect 7489 6496 7495 6560
rect 7179 6495 7495 6496
rect 9893 6560 10209 6561
rect 9893 6496 9899 6560
rect 9963 6496 9979 6560
rect 10043 6496 10059 6560
rect 10123 6496 10139 6560
rect 10203 6496 10209 6560
rect 9893 6495 10209 6496
rect 3108 6016 3424 6017
rect 3108 5952 3114 6016
rect 3178 5952 3194 6016
rect 3258 5952 3274 6016
rect 3338 5952 3354 6016
rect 3418 5952 3424 6016
rect 3108 5951 3424 5952
rect 5822 6016 6138 6017
rect 5822 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5988 6016
rect 6052 5952 6068 6016
rect 6132 5952 6138 6016
rect 5822 5951 6138 5952
rect 8536 6016 8852 6017
rect 8536 5952 8542 6016
rect 8606 5952 8622 6016
rect 8686 5952 8702 6016
rect 8766 5952 8782 6016
rect 8846 5952 8852 6016
rect 8536 5951 8852 5952
rect 11250 6016 11566 6017
rect 11250 5952 11256 6016
rect 11320 5952 11336 6016
rect 11400 5952 11416 6016
rect 11480 5952 11496 6016
rect 11560 5952 11566 6016
rect 11250 5951 11566 5952
rect 1751 5472 2067 5473
rect 1751 5408 1757 5472
rect 1821 5408 1837 5472
rect 1901 5408 1917 5472
rect 1981 5408 1997 5472
rect 2061 5408 2067 5472
rect 1751 5407 2067 5408
rect 4465 5472 4781 5473
rect 4465 5408 4471 5472
rect 4535 5408 4551 5472
rect 4615 5408 4631 5472
rect 4695 5408 4711 5472
rect 4775 5408 4781 5472
rect 4465 5407 4781 5408
rect 7179 5472 7495 5473
rect 7179 5408 7185 5472
rect 7249 5408 7265 5472
rect 7329 5408 7345 5472
rect 7409 5408 7425 5472
rect 7489 5408 7495 5472
rect 7179 5407 7495 5408
rect 9893 5472 10209 5473
rect 9893 5408 9899 5472
rect 9963 5408 9979 5472
rect 10043 5408 10059 5472
rect 10123 5408 10139 5472
rect 10203 5408 10209 5472
rect 9893 5407 10209 5408
rect 3108 4928 3424 4929
rect 3108 4864 3114 4928
rect 3178 4864 3194 4928
rect 3258 4864 3274 4928
rect 3338 4864 3354 4928
rect 3418 4864 3424 4928
rect 3108 4863 3424 4864
rect 5822 4928 6138 4929
rect 5822 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5988 4928
rect 6052 4864 6068 4928
rect 6132 4864 6138 4928
rect 5822 4863 6138 4864
rect 8536 4928 8852 4929
rect 8536 4864 8542 4928
rect 8606 4864 8622 4928
rect 8686 4864 8702 4928
rect 8766 4864 8782 4928
rect 8846 4864 8852 4928
rect 8536 4863 8852 4864
rect 11250 4928 11566 4929
rect 11250 4864 11256 4928
rect 11320 4864 11336 4928
rect 11400 4864 11416 4928
rect 11480 4864 11496 4928
rect 11560 4864 11566 4928
rect 11250 4863 11566 4864
rect 1751 4384 2067 4385
rect 1751 4320 1757 4384
rect 1821 4320 1837 4384
rect 1901 4320 1917 4384
rect 1981 4320 1997 4384
rect 2061 4320 2067 4384
rect 1751 4319 2067 4320
rect 4465 4384 4781 4385
rect 4465 4320 4471 4384
rect 4535 4320 4551 4384
rect 4615 4320 4631 4384
rect 4695 4320 4711 4384
rect 4775 4320 4781 4384
rect 4465 4319 4781 4320
rect 7179 4384 7495 4385
rect 7179 4320 7185 4384
rect 7249 4320 7265 4384
rect 7329 4320 7345 4384
rect 7409 4320 7425 4384
rect 7489 4320 7495 4384
rect 7179 4319 7495 4320
rect 9893 4384 10209 4385
rect 9893 4320 9899 4384
rect 9963 4320 9979 4384
rect 10043 4320 10059 4384
rect 10123 4320 10139 4384
rect 10203 4320 10209 4384
rect 9893 4319 10209 4320
rect 3108 3840 3424 3841
rect 3108 3776 3114 3840
rect 3178 3776 3194 3840
rect 3258 3776 3274 3840
rect 3338 3776 3354 3840
rect 3418 3776 3424 3840
rect 3108 3775 3424 3776
rect 5822 3840 6138 3841
rect 5822 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5988 3840
rect 6052 3776 6068 3840
rect 6132 3776 6138 3840
rect 5822 3775 6138 3776
rect 8536 3840 8852 3841
rect 8536 3776 8542 3840
rect 8606 3776 8622 3840
rect 8686 3776 8702 3840
rect 8766 3776 8782 3840
rect 8846 3776 8852 3840
rect 8536 3775 8852 3776
rect 11250 3840 11566 3841
rect 11250 3776 11256 3840
rect 11320 3776 11336 3840
rect 11400 3776 11416 3840
rect 11480 3776 11496 3840
rect 11560 3776 11566 3840
rect 11250 3775 11566 3776
rect 11237 3498 11303 3501
rect 11600 3498 12000 3528
rect 11237 3496 12000 3498
rect 11237 3440 11242 3496
rect 11298 3440 12000 3496
rect 11237 3438 12000 3440
rect 11237 3435 11303 3438
rect 11600 3408 12000 3438
rect 1751 3296 2067 3297
rect 1751 3232 1757 3296
rect 1821 3232 1837 3296
rect 1901 3232 1917 3296
rect 1981 3232 1997 3296
rect 2061 3232 2067 3296
rect 1751 3231 2067 3232
rect 4465 3296 4781 3297
rect 4465 3232 4471 3296
rect 4535 3232 4551 3296
rect 4615 3232 4631 3296
rect 4695 3232 4711 3296
rect 4775 3232 4781 3296
rect 4465 3231 4781 3232
rect 7179 3296 7495 3297
rect 7179 3232 7185 3296
rect 7249 3232 7265 3296
rect 7329 3232 7345 3296
rect 7409 3232 7425 3296
rect 7489 3232 7495 3296
rect 7179 3231 7495 3232
rect 9893 3296 10209 3297
rect 9893 3232 9899 3296
rect 9963 3232 9979 3296
rect 10043 3232 10059 3296
rect 10123 3232 10139 3296
rect 10203 3232 10209 3296
rect 9893 3231 10209 3232
rect 3108 2752 3424 2753
rect 3108 2688 3114 2752
rect 3178 2688 3194 2752
rect 3258 2688 3274 2752
rect 3338 2688 3354 2752
rect 3418 2688 3424 2752
rect 3108 2687 3424 2688
rect 5822 2752 6138 2753
rect 5822 2688 5828 2752
rect 5892 2688 5908 2752
rect 5972 2688 5988 2752
rect 6052 2688 6068 2752
rect 6132 2688 6138 2752
rect 5822 2687 6138 2688
rect 8536 2752 8852 2753
rect 8536 2688 8542 2752
rect 8606 2688 8622 2752
rect 8686 2688 8702 2752
rect 8766 2688 8782 2752
rect 8846 2688 8852 2752
rect 8536 2687 8852 2688
rect 11250 2752 11566 2753
rect 11250 2688 11256 2752
rect 11320 2688 11336 2752
rect 11400 2688 11416 2752
rect 11480 2688 11496 2752
rect 11560 2688 11566 2752
rect 11250 2687 11566 2688
rect 4061 2546 4127 2549
rect 5533 2546 5599 2549
rect 4061 2544 5599 2546
rect 4061 2488 4066 2544
rect 4122 2488 5538 2544
rect 5594 2488 5599 2544
rect 4061 2486 5599 2488
rect 4061 2483 4127 2486
rect 5533 2483 5599 2486
rect 1751 2208 2067 2209
rect 1751 2144 1757 2208
rect 1821 2144 1837 2208
rect 1901 2144 1917 2208
rect 1981 2144 1997 2208
rect 2061 2144 2067 2208
rect 1751 2143 2067 2144
rect 4465 2208 4781 2209
rect 4465 2144 4471 2208
rect 4535 2144 4551 2208
rect 4615 2144 4631 2208
rect 4695 2144 4711 2208
rect 4775 2144 4781 2208
rect 4465 2143 4781 2144
rect 7179 2208 7495 2209
rect 7179 2144 7185 2208
rect 7249 2144 7265 2208
rect 7329 2144 7345 2208
rect 7409 2144 7425 2208
rect 7489 2144 7495 2208
rect 7179 2143 7495 2144
rect 9893 2208 10209 2209
rect 9893 2144 9899 2208
rect 9963 2144 9979 2208
rect 10043 2144 10059 2208
rect 10123 2144 10139 2208
rect 10203 2144 10209 2208
rect 9893 2143 10209 2144
rect 3108 1664 3424 1665
rect 3108 1600 3114 1664
rect 3178 1600 3194 1664
rect 3258 1600 3274 1664
rect 3338 1600 3354 1664
rect 3418 1600 3424 1664
rect 3108 1599 3424 1600
rect 5822 1664 6138 1665
rect 5822 1600 5828 1664
rect 5892 1600 5908 1664
rect 5972 1600 5988 1664
rect 6052 1600 6068 1664
rect 6132 1600 6138 1664
rect 5822 1599 6138 1600
rect 8536 1664 8852 1665
rect 8536 1600 8542 1664
rect 8606 1600 8622 1664
rect 8686 1600 8702 1664
rect 8766 1600 8782 1664
rect 8846 1600 8852 1664
rect 8536 1599 8852 1600
rect 11250 1664 11566 1665
rect 11250 1600 11256 1664
rect 11320 1600 11336 1664
rect 11400 1600 11416 1664
rect 11480 1600 11496 1664
rect 11560 1600 11566 1664
rect 11250 1599 11566 1600
rect 1751 1120 2067 1121
rect 1751 1056 1757 1120
rect 1821 1056 1837 1120
rect 1901 1056 1917 1120
rect 1981 1056 1997 1120
rect 2061 1056 2067 1120
rect 1751 1055 2067 1056
rect 4465 1120 4781 1121
rect 4465 1056 4471 1120
rect 4535 1056 4551 1120
rect 4615 1056 4631 1120
rect 4695 1056 4711 1120
rect 4775 1056 4781 1120
rect 4465 1055 4781 1056
rect 7179 1120 7495 1121
rect 7179 1056 7185 1120
rect 7249 1056 7265 1120
rect 7329 1056 7345 1120
rect 7409 1056 7425 1120
rect 7489 1056 7495 1120
rect 7179 1055 7495 1056
rect 9893 1120 10209 1121
rect 9893 1056 9899 1120
rect 9963 1056 9979 1120
rect 10043 1056 10059 1120
rect 10123 1056 10139 1120
rect 10203 1056 10209 1120
rect 9893 1055 10209 1056
rect 3108 576 3424 577
rect 3108 512 3114 576
rect 3178 512 3194 576
rect 3258 512 3274 576
rect 3338 512 3354 576
rect 3418 512 3424 576
rect 3108 511 3424 512
rect 5822 576 6138 577
rect 5822 512 5828 576
rect 5892 512 5908 576
rect 5972 512 5988 576
rect 6052 512 6068 576
rect 6132 512 6138 576
rect 5822 511 6138 512
rect 8536 576 8852 577
rect 8536 512 8542 576
rect 8606 512 8622 576
rect 8686 512 8702 576
rect 8766 512 8782 576
rect 8846 512 8852 576
rect 8536 511 8852 512
rect 11250 576 11566 577
rect 11250 512 11256 576
rect 11320 512 11336 576
rect 11400 512 11416 576
rect 11480 512 11496 576
rect 11560 512 11566 576
rect 11250 511 11566 512
<< via3 >>
rect 3114 11452 3178 11456
rect 3114 11396 3118 11452
rect 3118 11396 3174 11452
rect 3174 11396 3178 11452
rect 3114 11392 3178 11396
rect 3194 11452 3258 11456
rect 3194 11396 3198 11452
rect 3198 11396 3254 11452
rect 3254 11396 3258 11452
rect 3194 11392 3258 11396
rect 3274 11452 3338 11456
rect 3274 11396 3278 11452
rect 3278 11396 3334 11452
rect 3334 11396 3338 11452
rect 3274 11392 3338 11396
rect 3354 11452 3418 11456
rect 3354 11396 3358 11452
rect 3358 11396 3414 11452
rect 3414 11396 3418 11452
rect 3354 11392 3418 11396
rect 5828 11452 5892 11456
rect 5828 11396 5832 11452
rect 5832 11396 5888 11452
rect 5888 11396 5892 11452
rect 5828 11392 5892 11396
rect 5908 11452 5972 11456
rect 5908 11396 5912 11452
rect 5912 11396 5968 11452
rect 5968 11396 5972 11452
rect 5908 11392 5972 11396
rect 5988 11452 6052 11456
rect 5988 11396 5992 11452
rect 5992 11396 6048 11452
rect 6048 11396 6052 11452
rect 5988 11392 6052 11396
rect 6068 11452 6132 11456
rect 6068 11396 6072 11452
rect 6072 11396 6128 11452
rect 6128 11396 6132 11452
rect 6068 11392 6132 11396
rect 8542 11452 8606 11456
rect 8542 11396 8546 11452
rect 8546 11396 8602 11452
rect 8602 11396 8606 11452
rect 8542 11392 8606 11396
rect 8622 11452 8686 11456
rect 8622 11396 8626 11452
rect 8626 11396 8682 11452
rect 8682 11396 8686 11452
rect 8622 11392 8686 11396
rect 8702 11452 8766 11456
rect 8702 11396 8706 11452
rect 8706 11396 8762 11452
rect 8762 11396 8766 11452
rect 8702 11392 8766 11396
rect 8782 11452 8846 11456
rect 8782 11396 8786 11452
rect 8786 11396 8842 11452
rect 8842 11396 8846 11452
rect 8782 11392 8846 11396
rect 11256 11452 11320 11456
rect 11256 11396 11260 11452
rect 11260 11396 11316 11452
rect 11316 11396 11320 11452
rect 11256 11392 11320 11396
rect 11336 11452 11400 11456
rect 11336 11396 11340 11452
rect 11340 11396 11396 11452
rect 11396 11396 11400 11452
rect 11336 11392 11400 11396
rect 11416 11452 11480 11456
rect 11416 11396 11420 11452
rect 11420 11396 11476 11452
rect 11476 11396 11480 11452
rect 11416 11392 11480 11396
rect 11496 11452 11560 11456
rect 11496 11396 11500 11452
rect 11500 11396 11556 11452
rect 11556 11396 11560 11452
rect 11496 11392 11560 11396
rect 1757 10908 1821 10912
rect 1757 10852 1761 10908
rect 1761 10852 1817 10908
rect 1817 10852 1821 10908
rect 1757 10848 1821 10852
rect 1837 10908 1901 10912
rect 1837 10852 1841 10908
rect 1841 10852 1897 10908
rect 1897 10852 1901 10908
rect 1837 10848 1901 10852
rect 1917 10908 1981 10912
rect 1917 10852 1921 10908
rect 1921 10852 1977 10908
rect 1977 10852 1981 10908
rect 1917 10848 1981 10852
rect 1997 10908 2061 10912
rect 1997 10852 2001 10908
rect 2001 10852 2057 10908
rect 2057 10852 2061 10908
rect 1997 10848 2061 10852
rect 4471 10908 4535 10912
rect 4471 10852 4475 10908
rect 4475 10852 4531 10908
rect 4531 10852 4535 10908
rect 4471 10848 4535 10852
rect 4551 10908 4615 10912
rect 4551 10852 4555 10908
rect 4555 10852 4611 10908
rect 4611 10852 4615 10908
rect 4551 10848 4615 10852
rect 4631 10908 4695 10912
rect 4631 10852 4635 10908
rect 4635 10852 4691 10908
rect 4691 10852 4695 10908
rect 4631 10848 4695 10852
rect 4711 10908 4775 10912
rect 4711 10852 4715 10908
rect 4715 10852 4771 10908
rect 4771 10852 4775 10908
rect 4711 10848 4775 10852
rect 7185 10908 7249 10912
rect 7185 10852 7189 10908
rect 7189 10852 7245 10908
rect 7245 10852 7249 10908
rect 7185 10848 7249 10852
rect 7265 10908 7329 10912
rect 7265 10852 7269 10908
rect 7269 10852 7325 10908
rect 7325 10852 7329 10908
rect 7265 10848 7329 10852
rect 7345 10908 7409 10912
rect 7345 10852 7349 10908
rect 7349 10852 7405 10908
rect 7405 10852 7409 10908
rect 7345 10848 7409 10852
rect 7425 10908 7489 10912
rect 7425 10852 7429 10908
rect 7429 10852 7485 10908
rect 7485 10852 7489 10908
rect 7425 10848 7489 10852
rect 9899 10908 9963 10912
rect 9899 10852 9903 10908
rect 9903 10852 9959 10908
rect 9959 10852 9963 10908
rect 9899 10848 9963 10852
rect 9979 10908 10043 10912
rect 9979 10852 9983 10908
rect 9983 10852 10039 10908
rect 10039 10852 10043 10908
rect 9979 10848 10043 10852
rect 10059 10908 10123 10912
rect 10059 10852 10063 10908
rect 10063 10852 10119 10908
rect 10119 10852 10123 10908
rect 10059 10848 10123 10852
rect 10139 10908 10203 10912
rect 10139 10852 10143 10908
rect 10143 10852 10199 10908
rect 10199 10852 10203 10908
rect 10139 10848 10203 10852
rect 3114 10364 3178 10368
rect 3114 10308 3118 10364
rect 3118 10308 3174 10364
rect 3174 10308 3178 10364
rect 3114 10304 3178 10308
rect 3194 10364 3258 10368
rect 3194 10308 3198 10364
rect 3198 10308 3254 10364
rect 3254 10308 3258 10364
rect 3194 10304 3258 10308
rect 3274 10364 3338 10368
rect 3274 10308 3278 10364
rect 3278 10308 3334 10364
rect 3334 10308 3338 10364
rect 3274 10304 3338 10308
rect 3354 10364 3418 10368
rect 3354 10308 3358 10364
rect 3358 10308 3414 10364
rect 3414 10308 3418 10364
rect 3354 10304 3418 10308
rect 5828 10364 5892 10368
rect 5828 10308 5832 10364
rect 5832 10308 5888 10364
rect 5888 10308 5892 10364
rect 5828 10304 5892 10308
rect 5908 10364 5972 10368
rect 5908 10308 5912 10364
rect 5912 10308 5968 10364
rect 5968 10308 5972 10364
rect 5908 10304 5972 10308
rect 5988 10364 6052 10368
rect 5988 10308 5992 10364
rect 5992 10308 6048 10364
rect 6048 10308 6052 10364
rect 5988 10304 6052 10308
rect 6068 10364 6132 10368
rect 6068 10308 6072 10364
rect 6072 10308 6128 10364
rect 6128 10308 6132 10364
rect 6068 10304 6132 10308
rect 8542 10364 8606 10368
rect 8542 10308 8546 10364
rect 8546 10308 8602 10364
rect 8602 10308 8606 10364
rect 8542 10304 8606 10308
rect 8622 10364 8686 10368
rect 8622 10308 8626 10364
rect 8626 10308 8682 10364
rect 8682 10308 8686 10364
rect 8622 10304 8686 10308
rect 8702 10364 8766 10368
rect 8702 10308 8706 10364
rect 8706 10308 8762 10364
rect 8762 10308 8766 10364
rect 8702 10304 8766 10308
rect 8782 10364 8846 10368
rect 8782 10308 8786 10364
rect 8786 10308 8842 10364
rect 8842 10308 8846 10364
rect 8782 10304 8846 10308
rect 11256 10364 11320 10368
rect 11256 10308 11260 10364
rect 11260 10308 11316 10364
rect 11316 10308 11320 10364
rect 11256 10304 11320 10308
rect 11336 10364 11400 10368
rect 11336 10308 11340 10364
rect 11340 10308 11396 10364
rect 11396 10308 11400 10364
rect 11336 10304 11400 10308
rect 11416 10364 11480 10368
rect 11416 10308 11420 10364
rect 11420 10308 11476 10364
rect 11476 10308 11480 10364
rect 11416 10304 11480 10308
rect 11496 10364 11560 10368
rect 11496 10308 11500 10364
rect 11500 10308 11556 10364
rect 11556 10308 11560 10364
rect 11496 10304 11560 10308
rect 1757 9820 1821 9824
rect 1757 9764 1761 9820
rect 1761 9764 1817 9820
rect 1817 9764 1821 9820
rect 1757 9760 1821 9764
rect 1837 9820 1901 9824
rect 1837 9764 1841 9820
rect 1841 9764 1897 9820
rect 1897 9764 1901 9820
rect 1837 9760 1901 9764
rect 1917 9820 1981 9824
rect 1917 9764 1921 9820
rect 1921 9764 1977 9820
rect 1977 9764 1981 9820
rect 1917 9760 1981 9764
rect 1997 9820 2061 9824
rect 1997 9764 2001 9820
rect 2001 9764 2057 9820
rect 2057 9764 2061 9820
rect 1997 9760 2061 9764
rect 4471 9820 4535 9824
rect 4471 9764 4475 9820
rect 4475 9764 4531 9820
rect 4531 9764 4535 9820
rect 4471 9760 4535 9764
rect 4551 9820 4615 9824
rect 4551 9764 4555 9820
rect 4555 9764 4611 9820
rect 4611 9764 4615 9820
rect 4551 9760 4615 9764
rect 4631 9820 4695 9824
rect 4631 9764 4635 9820
rect 4635 9764 4691 9820
rect 4691 9764 4695 9820
rect 4631 9760 4695 9764
rect 4711 9820 4775 9824
rect 4711 9764 4715 9820
rect 4715 9764 4771 9820
rect 4771 9764 4775 9820
rect 4711 9760 4775 9764
rect 7185 9820 7249 9824
rect 7185 9764 7189 9820
rect 7189 9764 7245 9820
rect 7245 9764 7249 9820
rect 7185 9760 7249 9764
rect 7265 9820 7329 9824
rect 7265 9764 7269 9820
rect 7269 9764 7325 9820
rect 7325 9764 7329 9820
rect 7265 9760 7329 9764
rect 7345 9820 7409 9824
rect 7345 9764 7349 9820
rect 7349 9764 7405 9820
rect 7405 9764 7409 9820
rect 7345 9760 7409 9764
rect 7425 9820 7489 9824
rect 7425 9764 7429 9820
rect 7429 9764 7485 9820
rect 7485 9764 7489 9820
rect 7425 9760 7489 9764
rect 9899 9820 9963 9824
rect 9899 9764 9903 9820
rect 9903 9764 9959 9820
rect 9959 9764 9963 9820
rect 9899 9760 9963 9764
rect 9979 9820 10043 9824
rect 9979 9764 9983 9820
rect 9983 9764 10039 9820
rect 10039 9764 10043 9820
rect 9979 9760 10043 9764
rect 10059 9820 10123 9824
rect 10059 9764 10063 9820
rect 10063 9764 10119 9820
rect 10119 9764 10123 9820
rect 10059 9760 10123 9764
rect 10139 9820 10203 9824
rect 10139 9764 10143 9820
rect 10143 9764 10199 9820
rect 10199 9764 10203 9820
rect 10139 9760 10203 9764
rect 3114 9276 3178 9280
rect 3114 9220 3118 9276
rect 3118 9220 3174 9276
rect 3174 9220 3178 9276
rect 3114 9216 3178 9220
rect 3194 9276 3258 9280
rect 3194 9220 3198 9276
rect 3198 9220 3254 9276
rect 3254 9220 3258 9276
rect 3194 9216 3258 9220
rect 3274 9276 3338 9280
rect 3274 9220 3278 9276
rect 3278 9220 3334 9276
rect 3334 9220 3338 9276
rect 3274 9216 3338 9220
rect 3354 9276 3418 9280
rect 3354 9220 3358 9276
rect 3358 9220 3414 9276
rect 3414 9220 3418 9276
rect 3354 9216 3418 9220
rect 5828 9276 5892 9280
rect 5828 9220 5832 9276
rect 5832 9220 5888 9276
rect 5888 9220 5892 9276
rect 5828 9216 5892 9220
rect 5908 9276 5972 9280
rect 5908 9220 5912 9276
rect 5912 9220 5968 9276
rect 5968 9220 5972 9276
rect 5908 9216 5972 9220
rect 5988 9276 6052 9280
rect 5988 9220 5992 9276
rect 5992 9220 6048 9276
rect 6048 9220 6052 9276
rect 5988 9216 6052 9220
rect 6068 9276 6132 9280
rect 6068 9220 6072 9276
rect 6072 9220 6128 9276
rect 6128 9220 6132 9276
rect 6068 9216 6132 9220
rect 8542 9276 8606 9280
rect 8542 9220 8546 9276
rect 8546 9220 8602 9276
rect 8602 9220 8606 9276
rect 8542 9216 8606 9220
rect 8622 9276 8686 9280
rect 8622 9220 8626 9276
rect 8626 9220 8682 9276
rect 8682 9220 8686 9276
rect 8622 9216 8686 9220
rect 8702 9276 8766 9280
rect 8702 9220 8706 9276
rect 8706 9220 8762 9276
rect 8762 9220 8766 9276
rect 8702 9216 8766 9220
rect 8782 9276 8846 9280
rect 8782 9220 8786 9276
rect 8786 9220 8842 9276
rect 8842 9220 8846 9276
rect 8782 9216 8846 9220
rect 11256 9276 11320 9280
rect 11256 9220 11260 9276
rect 11260 9220 11316 9276
rect 11316 9220 11320 9276
rect 11256 9216 11320 9220
rect 11336 9276 11400 9280
rect 11336 9220 11340 9276
rect 11340 9220 11396 9276
rect 11396 9220 11400 9276
rect 11336 9216 11400 9220
rect 11416 9276 11480 9280
rect 11416 9220 11420 9276
rect 11420 9220 11476 9276
rect 11476 9220 11480 9276
rect 11416 9216 11480 9220
rect 11496 9276 11560 9280
rect 11496 9220 11500 9276
rect 11500 9220 11556 9276
rect 11556 9220 11560 9276
rect 11496 9216 11560 9220
rect 1757 8732 1821 8736
rect 1757 8676 1761 8732
rect 1761 8676 1817 8732
rect 1817 8676 1821 8732
rect 1757 8672 1821 8676
rect 1837 8732 1901 8736
rect 1837 8676 1841 8732
rect 1841 8676 1897 8732
rect 1897 8676 1901 8732
rect 1837 8672 1901 8676
rect 1917 8732 1981 8736
rect 1917 8676 1921 8732
rect 1921 8676 1977 8732
rect 1977 8676 1981 8732
rect 1917 8672 1981 8676
rect 1997 8732 2061 8736
rect 1997 8676 2001 8732
rect 2001 8676 2057 8732
rect 2057 8676 2061 8732
rect 1997 8672 2061 8676
rect 4471 8732 4535 8736
rect 4471 8676 4475 8732
rect 4475 8676 4531 8732
rect 4531 8676 4535 8732
rect 4471 8672 4535 8676
rect 4551 8732 4615 8736
rect 4551 8676 4555 8732
rect 4555 8676 4611 8732
rect 4611 8676 4615 8732
rect 4551 8672 4615 8676
rect 4631 8732 4695 8736
rect 4631 8676 4635 8732
rect 4635 8676 4691 8732
rect 4691 8676 4695 8732
rect 4631 8672 4695 8676
rect 4711 8732 4775 8736
rect 4711 8676 4715 8732
rect 4715 8676 4771 8732
rect 4771 8676 4775 8732
rect 4711 8672 4775 8676
rect 7185 8732 7249 8736
rect 7185 8676 7189 8732
rect 7189 8676 7245 8732
rect 7245 8676 7249 8732
rect 7185 8672 7249 8676
rect 7265 8732 7329 8736
rect 7265 8676 7269 8732
rect 7269 8676 7325 8732
rect 7325 8676 7329 8732
rect 7265 8672 7329 8676
rect 7345 8732 7409 8736
rect 7345 8676 7349 8732
rect 7349 8676 7405 8732
rect 7405 8676 7409 8732
rect 7345 8672 7409 8676
rect 7425 8732 7489 8736
rect 7425 8676 7429 8732
rect 7429 8676 7485 8732
rect 7485 8676 7489 8732
rect 7425 8672 7489 8676
rect 9899 8732 9963 8736
rect 9899 8676 9903 8732
rect 9903 8676 9959 8732
rect 9959 8676 9963 8732
rect 9899 8672 9963 8676
rect 9979 8732 10043 8736
rect 9979 8676 9983 8732
rect 9983 8676 10039 8732
rect 10039 8676 10043 8732
rect 9979 8672 10043 8676
rect 10059 8732 10123 8736
rect 10059 8676 10063 8732
rect 10063 8676 10119 8732
rect 10119 8676 10123 8732
rect 10059 8672 10123 8676
rect 10139 8732 10203 8736
rect 10139 8676 10143 8732
rect 10143 8676 10199 8732
rect 10199 8676 10203 8732
rect 10139 8672 10203 8676
rect 3114 8188 3178 8192
rect 3114 8132 3118 8188
rect 3118 8132 3174 8188
rect 3174 8132 3178 8188
rect 3114 8128 3178 8132
rect 3194 8188 3258 8192
rect 3194 8132 3198 8188
rect 3198 8132 3254 8188
rect 3254 8132 3258 8188
rect 3194 8128 3258 8132
rect 3274 8188 3338 8192
rect 3274 8132 3278 8188
rect 3278 8132 3334 8188
rect 3334 8132 3338 8188
rect 3274 8128 3338 8132
rect 3354 8188 3418 8192
rect 3354 8132 3358 8188
rect 3358 8132 3414 8188
rect 3414 8132 3418 8188
rect 3354 8128 3418 8132
rect 5828 8188 5892 8192
rect 5828 8132 5832 8188
rect 5832 8132 5888 8188
rect 5888 8132 5892 8188
rect 5828 8128 5892 8132
rect 5908 8188 5972 8192
rect 5908 8132 5912 8188
rect 5912 8132 5968 8188
rect 5968 8132 5972 8188
rect 5908 8128 5972 8132
rect 5988 8188 6052 8192
rect 5988 8132 5992 8188
rect 5992 8132 6048 8188
rect 6048 8132 6052 8188
rect 5988 8128 6052 8132
rect 6068 8188 6132 8192
rect 6068 8132 6072 8188
rect 6072 8132 6128 8188
rect 6128 8132 6132 8188
rect 6068 8128 6132 8132
rect 8542 8188 8606 8192
rect 8542 8132 8546 8188
rect 8546 8132 8602 8188
rect 8602 8132 8606 8188
rect 8542 8128 8606 8132
rect 8622 8188 8686 8192
rect 8622 8132 8626 8188
rect 8626 8132 8682 8188
rect 8682 8132 8686 8188
rect 8622 8128 8686 8132
rect 8702 8188 8766 8192
rect 8702 8132 8706 8188
rect 8706 8132 8762 8188
rect 8762 8132 8766 8188
rect 8702 8128 8766 8132
rect 8782 8188 8846 8192
rect 8782 8132 8786 8188
rect 8786 8132 8842 8188
rect 8842 8132 8846 8188
rect 8782 8128 8846 8132
rect 11256 8188 11320 8192
rect 11256 8132 11260 8188
rect 11260 8132 11316 8188
rect 11316 8132 11320 8188
rect 11256 8128 11320 8132
rect 11336 8188 11400 8192
rect 11336 8132 11340 8188
rect 11340 8132 11396 8188
rect 11396 8132 11400 8188
rect 11336 8128 11400 8132
rect 11416 8188 11480 8192
rect 11416 8132 11420 8188
rect 11420 8132 11476 8188
rect 11476 8132 11480 8188
rect 11416 8128 11480 8132
rect 11496 8188 11560 8192
rect 11496 8132 11500 8188
rect 11500 8132 11556 8188
rect 11556 8132 11560 8188
rect 11496 8128 11560 8132
rect 1757 7644 1821 7648
rect 1757 7588 1761 7644
rect 1761 7588 1817 7644
rect 1817 7588 1821 7644
rect 1757 7584 1821 7588
rect 1837 7644 1901 7648
rect 1837 7588 1841 7644
rect 1841 7588 1897 7644
rect 1897 7588 1901 7644
rect 1837 7584 1901 7588
rect 1917 7644 1981 7648
rect 1917 7588 1921 7644
rect 1921 7588 1977 7644
rect 1977 7588 1981 7644
rect 1917 7584 1981 7588
rect 1997 7644 2061 7648
rect 1997 7588 2001 7644
rect 2001 7588 2057 7644
rect 2057 7588 2061 7644
rect 1997 7584 2061 7588
rect 4471 7644 4535 7648
rect 4471 7588 4475 7644
rect 4475 7588 4531 7644
rect 4531 7588 4535 7644
rect 4471 7584 4535 7588
rect 4551 7644 4615 7648
rect 4551 7588 4555 7644
rect 4555 7588 4611 7644
rect 4611 7588 4615 7644
rect 4551 7584 4615 7588
rect 4631 7644 4695 7648
rect 4631 7588 4635 7644
rect 4635 7588 4691 7644
rect 4691 7588 4695 7644
rect 4631 7584 4695 7588
rect 4711 7644 4775 7648
rect 4711 7588 4715 7644
rect 4715 7588 4771 7644
rect 4771 7588 4775 7644
rect 4711 7584 4775 7588
rect 7185 7644 7249 7648
rect 7185 7588 7189 7644
rect 7189 7588 7245 7644
rect 7245 7588 7249 7644
rect 7185 7584 7249 7588
rect 7265 7644 7329 7648
rect 7265 7588 7269 7644
rect 7269 7588 7325 7644
rect 7325 7588 7329 7644
rect 7265 7584 7329 7588
rect 7345 7644 7409 7648
rect 7345 7588 7349 7644
rect 7349 7588 7405 7644
rect 7405 7588 7409 7644
rect 7345 7584 7409 7588
rect 7425 7644 7489 7648
rect 7425 7588 7429 7644
rect 7429 7588 7485 7644
rect 7485 7588 7489 7644
rect 7425 7584 7489 7588
rect 9899 7644 9963 7648
rect 9899 7588 9903 7644
rect 9903 7588 9959 7644
rect 9959 7588 9963 7644
rect 9899 7584 9963 7588
rect 9979 7644 10043 7648
rect 9979 7588 9983 7644
rect 9983 7588 10039 7644
rect 10039 7588 10043 7644
rect 9979 7584 10043 7588
rect 10059 7644 10123 7648
rect 10059 7588 10063 7644
rect 10063 7588 10119 7644
rect 10119 7588 10123 7644
rect 10059 7584 10123 7588
rect 10139 7644 10203 7648
rect 10139 7588 10143 7644
rect 10143 7588 10199 7644
rect 10199 7588 10203 7644
rect 10139 7584 10203 7588
rect 3114 7100 3178 7104
rect 3114 7044 3118 7100
rect 3118 7044 3174 7100
rect 3174 7044 3178 7100
rect 3114 7040 3178 7044
rect 3194 7100 3258 7104
rect 3194 7044 3198 7100
rect 3198 7044 3254 7100
rect 3254 7044 3258 7100
rect 3194 7040 3258 7044
rect 3274 7100 3338 7104
rect 3274 7044 3278 7100
rect 3278 7044 3334 7100
rect 3334 7044 3338 7100
rect 3274 7040 3338 7044
rect 3354 7100 3418 7104
rect 3354 7044 3358 7100
rect 3358 7044 3414 7100
rect 3414 7044 3418 7100
rect 3354 7040 3418 7044
rect 5828 7100 5892 7104
rect 5828 7044 5832 7100
rect 5832 7044 5888 7100
rect 5888 7044 5892 7100
rect 5828 7040 5892 7044
rect 5908 7100 5972 7104
rect 5908 7044 5912 7100
rect 5912 7044 5968 7100
rect 5968 7044 5972 7100
rect 5908 7040 5972 7044
rect 5988 7100 6052 7104
rect 5988 7044 5992 7100
rect 5992 7044 6048 7100
rect 6048 7044 6052 7100
rect 5988 7040 6052 7044
rect 6068 7100 6132 7104
rect 6068 7044 6072 7100
rect 6072 7044 6128 7100
rect 6128 7044 6132 7100
rect 6068 7040 6132 7044
rect 8542 7100 8606 7104
rect 8542 7044 8546 7100
rect 8546 7044 8602 7100
rect 8602 7044 8606 7100
rect 8542 7040 8606 7044
rect 8622 7100 8686 7104
rect 8622 7044 8626 7100
rect 8626 7044 8682 7100
rect 8682 7044 8686 7100
rect 8622 7040 8686 7044
rect 8702 7100 8766 7104
rect 8702 7044 8706 7100
rect 8706 7044 8762 7100
rect 8762 7044 8766 7100
rect 8702 7040 8766 7044
rect 8782 7100 8846 7104
rect 8782 7044 8786 7100
rect 8786 7044 8842 7100
rect 8842 7044 8846 7100
rect 8782 7040 8846 7044
rect 11256 7100 11320 7104
rect 11256 7044 11260 7100
rect 11260 7044 11316 7100
rect 11316 7044 11320 7100
rect 11256 7040 11320 7044
rect 11336 7100 11400 7104
rect 11336 7044 11340 7100
rect 11340 7044 11396 7100
rect 11396 7044 11400 7100
rect 11336 7040 11400 7044
rect 11416 7100 11480 7104
rect 11416 7044 11420 7100
rect 11420 7044 11476 7100
rect 11476 7044 11480 7100
rect 11416 7040 11480 7044
rect 11496 7100 11560 7104
rect 11496 7044 11500 7100
rect 11500 7044 11556 7100
rect 11556 7044 11560 7100
rect 11496 7040 11560 7044
rect 1757 6556 1821 6560
rect 1757 6500 1761 6556
rect 1761 6500 1817 6556
rect 1817 6500 1821 6556
rect 1757 6496 1821 6500
rect 1837 6556 1901 6560
rect 1837 6500 1841 6556
rect 1841 6500 1897 6556
rect 1897 6500 1901 6556
rect 1837 6496 1901 6500
rect 1917 6556 1981 6560
rect 1917 6500 1921 6556
rect 1921 6500 1977 6556
rect 1977 6500 1981 6556
rect 1917 6496 1981 6500
rect 1997 6556 2061 6560
rect 1997 6500 2001 6556
rect 2001 6500 2057 6556
rect 2057 6500 2061 6556
rect 1997 6496 2061 6500
rect 4471 6556 4535 6560
rect 4471 6500 4475 6556
rect 4475 6500 4531 6556
rect 4531 6500 4535 6556
rect 4471 6496 4535 6500
rect 4551 6556 4615 6560
rect 4551 6500 4555 6556
rect 4555 6500 4611 6556
rect 4611 6500 4615 6556
rect 4551 6496 4615 6500
rect 4631 6556 4695 6560
rect 4631 6500 4635 6556
rect 4635 6500 4691 6556
rect 4691 6500 4695 6556
rect 4631 6496 4695 6500
rect 4711 6556 4775 6560
rect 4711 6500 4715 6556
rect 4715 6500 4771 6556
rect 4771 6500 4775 6556
rect 4711 6496 4775 6500
rect 7185 6556 7249 6560
rect 7185 6500 7189 6556
rect 7189 6500 7245 6556
rect 7245 6500 7249 6556
rect 7185 6496 7249 6500
rect 7265 6556 7329 6560
rect 7265 6500 7269 6556
rect 7269 6500 7325 6556
rect 7325 6500 7329 6556
rect 7265 6496 7329 6500
rect 7345 6556 7409 6560
rect 7345 6500 7349 6556
rect 7349 6500 7405 6556
rect 7405 6500 7409 6556
rect 7345 6496 7409 6500
rect 7425 6556 7489 6560
rect 7425 6500 7429 6556
rect 7429 6500 7485 6556
rect 7485 6500 7489 6556
rect 7425 6496 7489 6500
rect 9899 6556 9963 6560
rect 9899 6500 9903 6556
rect 9903 6500 9959 6556
rect 9959 6500 9963 6556
rect 9899 6496 9963 6500
rect 9979 6556 10043 6560
rect 9979 6500 9983 6556
rect 9983 6500 10039 6556
rect 10039 6500 10043 6556
rect 9979 6496 10043 6500
rect 10059 6556 10123 6560
rect 10059 6500 10063 6556
rect 10063 6500 10119 6556
rect 10119 6500 10123 6556
rect 10059 6496 10123 6500
rect 10139 6556 10203 6560
rect 10139 6500 10143 6556
rect 10143 6500 10199 6556
rect 10199 6500 10203 6556
rect 10139 6496 10203 6500
rect 3114 6012 3178 6016
rect 3114 5956 3118 6012
rect 3118 5956 3174 6012
rect 3174 5956 3178 6012
rect 3114 5952 3178 5956
rect 3194 6012 3258 6016
rect 3194 5956 3198 6012
rect 3198 5956 3254 6012
rect 3254 5956 3258 6012
rect 3194 5952 3258 5956
rect 3274 6012 3338 6016
rect 3274 5956 3278 6012
rect 3278 5956 3334 6012
rect 3334 5956 3338 6012
rect 3274 5952 3338 5956
rect 3354 6012 3418 6016
rect 3354 5956 3358 6012
rect 3358 5956 3414 6012
rect 3414 5956 3418 6012
rect 3354 5952 3418 5956
rect 5828 6012 5892 6016
rect 5828 5956 5832 6012
rect 5832 5956 5888 6012
rect 5888 5956 5892 6012
rect 5828 5952 5892 5956
rect 5908 6012 5972 6016
rect 5908 5956 5912 6012
rect 5912 5956 5968 6012
rect 5968 5956 5972 6012
rect 5908 5952 5972 5956
rect 5988 6012 6052 6016
rect 5988 5956 5992 6012
rect 5992 5956 6048 6012
rect 6048 5956 6052 6012
rect 5988 5952 6052 5956
rect 6068 6012 6132 6016
rect 6068 5956 6072 6012
rect 6072 5956 6128 6012
rect 6128 5956 6132 6012
rect 6068 5952 6132 5956
rect 8542 6012 8606 6016
rect 8542 5956 8546 6012
rect 8546 5956 8602 6012
rect 8602 5956 8606 6012
rect 8542 5952 8606 5956
rect 8622 6012 8686 6016
rect 8622 5956 8626 6012
rect 8626 5956 8682 6012
rect 8682 5956 8686 6012
rect 8622 5952 8686 5956
rect 8702 6012 8766 6016
rect 8702 5956 8706 6012
rect 8706 5956 8762 6012
rect 8762 5956 8766 6012
rect 8702 5952 8766 5956
rect 8782 6012 8846 6016
rect 8782 5956 8786 6012
rect 8786 5956 8842 6012
rect 8842 5956 8846 6012
rect 8782 5952 8846 5956
rect 11256 6012 11320 6016
rect 11256 5956 11260 6012
rect 11260 5956 11316 6012
rect 11316 5956 11320 6012
rect 11256 5952 11320 5956
rect 11336 6012 11400 6016
rect 11336 5956 11340 6012
rect 11340 5956 11396 6012
rect 11396 5956 11400 6012
rect 11336 5952 11400 5956
rect 11416 6012 11480 6016
rect 11416 5956 11420 6012
rect 11420 5956 11476 6012
rect 11476 5956 11480 6012
rect 11416 5952 11480 5956
rect 11496 6012 11560 6016
rect 11496 5956 11500 6012
rect 11500 5956 11556 6012
rect 11556 5956 11560 6012
rect 11496 5952 11560 5956
rect 1757 5468 1821 5472
rect 1757 5412 1761 5468
rect 1761 5412 1817 5468
rect 1817 5412 1821 5468
rect 1757 5408 1821 5412
rect 1837 5468 1901 5472
rect 1837 5412 1841 5468
rect 1841 5412 1897 5468
rect 1897 5412 1901 5468
rect 1837 5408 1901 5412
rect 1917 5468 1981 5472
rect 1917 5412 1921 5468
rect 1921 5412 1977 5468
rect 1977 5412 1981 5468
rect 1917 5408 1981 5412
rect 1997 5468 2061 5472
rect 1997 5412 2001 5468
rect 2001 5412 2057 5468
rect 2057 5412 2061 5468
rect 1997 5408 2061 5412
rect 4471 5468 4535 5472
rect 4471 5412 4475 5468
rect 4475 5412 4531 5468
rect 4531 5412 4535 5468
rect 4471 5408 4535 5412
rect 4551 5468 4615 5472
rect 4551 5412 4555 5468
rect 4555 5412 4611 5468
rect 4611 5412 4615 5468
rect 4551 5408 4615 5412
rect 4631 5468 4695 5472
rect 4631 5412 4635 5468
rect 4635 5412 4691 5468
rect 4691 5412 4695 5468
rect 4631 5408 4695 5412
rect 4711 5468 4775 5472
rect 4711 5412 4715 5468
rect 4715 5412 4771 5468
rect 4771 5412 4775 5468
rect 4711 5408 4775 5412
rect 7185 5468 7249 5472
rect 7185 5412 7189 5468
rect 7189 5412 7245 5468
rect 7245 5412 7249 5468
rect 7185 5408 7249 5412
rect 7265 5468 7329 5472
rect 7265 5412 7269 5468
rect 7269 5412 7325 5468
rect 7325 5412 7329 5468
rect 7265 5408 7329 5412
rect 7345 5468 7409 5472
rect 7345 5412 7349 5468
rect 7349 5412 7405 5468
rect 7405 5412 7409 5468
rect 7345 5408 7409 5412
rect 7425 5468 7489 5472
rect 7425 5412 7429 5468
rect 7429 5412 7485 5468
rect 7485 5412 7489 5468
rect 7425 5408 7489 5412
rect 9899 5468 9963 5472
rect 9899 5412 9903 5468
rect 9903 5412 9959 5468
rect 9959 5412 9963 5468
rect 9899 5408 9963 5412
rect 9979 5468 10043 5472
rect 9979 5412 9983 5468
rect 9983 5412 10039 5468
rect 10039 5412 10043 5468
rect 9979 5408 10043 5412
rect 10059 5468 10123 5472
rect 10059 5412 10063 5468
rect 10063 5412 10119 5468
rect 10119 5412 10123 5468
rect 10059 5408 10123 5412
rect 10139 5468 10203 5472
rect 10139 5412 10143 5468
rect 10143 5412 10199 5468
rect 10199 5412 10203 5468
rect 10139 5408 10203 5412
rect 3114 4924 3178 4928
rect 3114 4868 3118 4924
rect 3118 4868 3174 4924
rect 3174 4868 3178 4924
rect 3114 4864 3178 4868
rect 3194 4924 3258 4928
rect 3194 4868 3198 4924
rect 3198 4868 3254 4924
rect 3254 4868 3258 4924
rect 3194 4864 3258 4868
rect 3274 4924 3338 4928
rect 3274 4868 3278 4924
rect 3278 4868 3334 4924
rect 3334 4868 3338 4924
rect 3274 4864 3338 4868
rect 3354 4924 3418 4928
rect 3354 4868 3358 4924
rect 3358 4868 3414 4924
rect 3414 4868 3418 4924
rect 3354 4864 3418 4868
rect 5828 4924 5892 4928
rect 5828 4868 5832 4924
rect 5832 4868 5888 4924
rect 5888 4868 5892 4924
rect 5828 4864 5892 4868
rect 5908 4924 5972 4928
rect 5908 4868 5912 4924
rect 5912 4868 5968 4924
rect 5968 4868 5972 4924
rect 5908 4864 5972 4868
rect 5988 4924 6052 4928
rect 5988 4868 5992 4924
rect 5992 4868 6048 4924
rect 6048 4868 6052 4924
rect 5988 4864 6052 4868
rect 6068 4924 6132 4928
rect 6068 4868 6072 4924
rect 6072 4868 6128 4924
rect 6128 4868 6132 4924
rect 6068 4864 6132 4868
rect 8542 4924 8606 4928
rect 8542 4868 8546 4924
rect 8546 4868 8602 4924
rect 8602 4868 8606 4924
rect 8542 4864 8606 4868
rect 8622 4924 8686 4928
rect 8622 4868 8626 4924
rect 8626 4868 8682 4924
rect 8682 4868 8686 4924
rect 8622 4864 8686 4868
rect 8702 4924 8766 4928
rect 8702 4868 8706 4924
rect 8706 4868 8762 4924
rect 8762 4868 8766 4924
rect 8702 4864 8766 4868
rect 8782 4924 8846 4928
rect 8782 4868 8786 4924
rect 8786 4868 8842 4924
rect 8842 4868 8846 4924
rect 8782 4864 8846 4868
rect 11256 4924 11320 4928
rect 11256 4868 11260 4924
rect 11260 4868 11316 4924
rect 11316 4868 11320 4924
rect 11256 4864 11320 4868
rect 11336 4924 11400 4928
rect 11336 4868 11340 4924
rect 11340 4868 11396 4924
rect 11396 4868 11400 4924
rect 11336 4864 11400 4868
rect 11416 4924 11480 4928
rect 11416 4868 11420 4924
rect 11420 4868 11476 4924
rect 11476 4868 11480 4924
rect 11416 4864 11480 4868
rect 11496 4924 11560 4928
rect 11496 4868 11500 4924
rect 11500 4868 11556 4924
rect 11556 4868 11560 4924
rect 11496 4864 11560 4868
rect 1757 4380 1821 4384
rect 1757 4324 1761 4380
rect 1761 4324 1817 4380
rect 1817 4324 1821 4380
rect 1757 4320 1821 4324
rect 1837 4380 1901 4384
rect 1837 4324 1841 4380
rect 1841 4324 1897 4380
rect 1897 4324 1901 4380
rect 1837 4320 1901 4324
rect 1917 4380 1981 4384
rect 1917 4324 1921 4380
rect 1921 4324 1977 4380
rect 1977 4324 1981 4380
rect 1917 4320 1981 4324
rect 1997 4380 2061 4384
rect 1997 4324 2001 4380
rect 2001 4324 2057 4380
rect 2057 4324 2061 4380
rect 1997 4320 2061 4324
rect 4471 4380 4535 4384
rect 4471 4324 4475 4380
rect 4475 4324 4531 4380
rect 4531 4324 4535 4380
rect 4471 4320 4535 4324
rect 4551 4380 4615 4384
rect 4551 4324 4555 4380
rect 4555 4324 4611 4380
rect 4611 4324 4615 4380
rect 4551 4320 4615 4324
rect 4631 4380 4695 4384
rect 4631 4324 4635 4380
rect 4635 4324 4691 4380
rect 4691 4324 4695 4380
rect 4631 4320 4695 4324
rect 4711 4380 4775 4384
rect 4711 4324 4715 4380
rect 4715 4324 4771 4380
rect 4771 4324 4775 4380
rect 4711 4320 4775 4324
rect 7185 4380 7249 4384
rect 7185 4324 7189 4380
rect 7189 4324 7245 4380
rect 7245 4324 7249 4380
rect 7185 4320 7249 4324
rect 7265 4380 7329 4384
rect 7265 4324 7269 4380
rect 7269 4324 7325 4380
rect 7325 4324 7329 4380
rect 7265 4320 7329 4324
rect 7345 4380 7409 4384
rect 7345 4324 7349 4380
rect 7349 4324 7405 4380
rect 7405 4324 7409 4380
rect 7345 4320 7409 4324
rect 7425 4380 7489 4384
rect 7425 4324 7429 4380
rect 7429 4324 7485 4380
rect 7485 4324 7489 4380
rect 7425 4320 7489 4324
rect 9899 4380 9963 4384
rect 9899 4324 9903 4380
rect 9903 4324 9959 4380
rect 9959 4324 9963 4380
rect 9899 4320 9963 4324
rect 9979 4380 10043 4384
rect 9979 4324 9983 4380
rect 9983 4324 10039 4380
rect 10039 4324 10043 4380
rect 9979 4320 10043 4324
rect 10059 4380 10123 4384
rect 10059 4324 10063 4380
rect 10063 4324 10119 4380
rect 10119 4324 10123 4380
rect 10059 4320 10123 4324
rect 10139 4380 10203 4384
rect 10139 4324 10143 4380
rect 10143 4324 10199 4380
rect 10199 4324 10203 4380
rect 10139 4320 10203 4324
rect 3114 3836 3178 3840
rect 3114 3780 3118 3836
rect 3118 3780 3174 3836
rect 3174 3780 3178 3836
rect 3114 3776 3178 3780
rect 3194 3836 3258 3840
rect 3194 3780 3198 3836
rect 3198 3780 3254 3836
rect 3254 3780 3258 3836
rect 3194 3776 3258 3780
rect 3274 3836 3338 3840
rect 3274 3780 3278 3836
rect 3278 3780 3334 3836
rect 3334 3780 3338 3836
rect 3274 3776 3338 3780
rect 3354 3836 3418 3840
rect 3354 3780 3358 3836
rect 3358 3780 3414 3836
rect 3414 3780 3418 3836
rect 3354 3776 3418 3780
rect 5828 3836 5892 3840
rect 5828 3780 5832 3836
rect 5832 3780 5888 3836
rect 5888 3780 5892 3836
rect 5828 3776 5892 3780
rect 5908 3836 5972 3840
rect 5908 3780 5912 3836
rect 5912 3780 5968 3836
rect 5968 3780 5972 3836
rect 5908 3776 5972 3780
rect 5988 3836 6052 3840
rect 5988 3780 5992 3836
rect 5992 3780 6048 3836
rect 6048 3780 6052 3836
rect 5988 3776 6052 3780
rect 6068 3836 6132 3840
rect 6068 3780 6072 3836
rect 6072 3780 6128 3836
rect 6128 3780 6132 3836
rect 6068 3776 6132 3780
rect 8542 3836 8606 3840
rect 8542 3780 8546 3836
rect 8546 3780 8602 3836
rect 8602 3780 8606 3836
rect 8542 3776 8606 3780
rect 8622 3836 8686 3840
rect 8622 3780 8626 3836
rect 8626 3780 8682 3836
rect 8682 3780 8686 3836
rect 8622 3776 8686 3780
rect 8702 3836 8766 3840
rect 8702 3780 8706 3836
rect 8706 3780 8762 3836
rect 8762 3780 8766 3836
rect 8702 3776 8766 3780
rect 8782 3836 8846 3840
rect 8782 3780 8786 3836
rect 8786 3780 8842 3836
rect 8842 3780 8846 3836
rect 8782 3776 8846 3780
rect 11256 3836 11320 3840
rect 11256 3780 11260 3836
rect 11260 3780 11316 3836
rect 11316 3780 11320 3836
rect 11256 3776 11320 3780
rect 11336 3836 11400 3840
rect 11336 3780 11340 3836
rect 11340 3780 11396 3836
rect 11396 3780 11400 3836
rect 11336 3776 11400 3780
rect 11416 3836 11480 3840
rect 11416 3780 11420 3836
rect 11420 3780 11476 3836
rect 11476 3780 11480 3836
rect 11416 3776 11480 3780
rect 11496 3836 11560 3840
rect 11496 3780 11500 3836
rect 11500 3780 11556 3836
rect 11556 3780 11560 3836
rect 11496 3776 11560 3780
rect 1757 3292 1821 3296
rect 1757 3236 1761 3292
rect 1761 3236 1817 3292
rect 1817 3236 1821 3292
rect 1757 3232 1821 3236
rect 1837 3292 1901 3296
rect 1837 3236 1841 3292
rect 1841 3236 1897 3292
rect 1897 3236 1901 3292
rect 1837 3232 1901 3236
rect 1917 3292 1981 3296
rect 1917 3236 1921 3292
rect 1921 3236 1977 3292
rect 1977 3236 1981 3292
rect 1917 3232 1981 3236
rect 1997 3292 2061 3296
rect 1997 3236 2001 3292
rect 2001 3236 2057 3292
rect 2057 3236 2061 3292
rect 1997 3232 2061 3236
rect 4471 3292 4535 3296
rect 4471 3236 4475 3292
rect 4475 3236 4531 3292
rect 4531 3236 4535 3292
rect 4471 3232 4535 3236
rect 4551 3292 4615 3296
rect 4551 3236 4555 3292
rect 4555 3236 4611 3292
rect 4611 3236 4615 3292
rect 4551 3232 4615 3236
rect 4631 3292 4695 3296
rect 4631 3236 4635 3292
rect 4635 3236 4691 3292
rect 4691 3236 4695 3292
rect 4631 3232 4695 3236
rect 4711 3292 4775 3296
rect 4711 3236 4715 3292
rect 4715 3236 4771 3292
rect 4771 3236 4775 3292
rect 4711 3232 4775 3236
rect 7185 3292 7249 3296
rect 7185 3236 7189 3292
rect 7189 3236 7245 3292
rect 7245 3236 7249 3292
rect 7185 3232 7249 3236
rect 7265 3292 7329 3296
rect 7265 3236 7269 3292
rect 7269 3236 7325 3292
rect 7325 3236 7329 3292
rect 7265 3232 7329 3236
rect 7345 3292 7409 3296
rect 7345 3236 7349 3292
rect 7349 3236 7405 3292
rect 7405 3236 7409 3292
rect 7345 3232 7409 3236
rect 7425 3292 7489 3296
rect 7425 3236 7429 3292
rect 7429 3236 7485 3292
rect 7485 3236 7489 3292
rect 7425 3232 7489 3236
rect 9899 3292 9963 3296
rect 9899 3236 9903 3292
rect 9903 3236 9959 3292
rect 9959 3236 9963 3292
rect 9899 3232 9963 3236
rect 9979 3292 10043 3296
rect 9979 3236 9983 3292
rect 9983 3236 10039 3292
rect 10039 3236 10043 3292
rect 9979 3232 10043 3236
rect 10059 3292 10123 3296
rect 10059 3236 10063 3292
rect 10063 3236 10119 3292
rect 10119 3236 10123 3292
rect 10059 3232 10123 3236
rect 10139 3292 10203 3296
rect 10139 3236 10143 3292
rect 10143 3236 10199 3292
rect 10199 3236 10203 3292
rect 10139 3232 10203 3236
rect 3114 2748 3178 2752
rect 3114 2692 3118 2748
rect 3118 2692 3174 2748
rect 3174 2692 3178 2748
rect 3114 2688 3178 2692
rect 3194 2748 3258 2752
rect 3194 2692 3198 2748
rect 3198 2692 3254 2748
rect 3254 2692 3258 2748
rect 3194 2688 3258 2692
rect 3274 2748 3338 2752
rect 3274 2692 3278 2748
rect 3278 2692 3334 2748
rect 3334 2692 3338 2748
rect 3274 2688 3338 2692
rect 3354 2748 3418 2752
rect 3354 2692 3358 2748
rect 3358 2692 3414 2748
rect 3414 2692 3418 2748
rect 3354 2688 3418 2692
rect 5828 2748 5892 2752
rect 5828 2692 5832 2748
rect 5832 2692 5888 2748
rect 5888 2692 5892 2748
rect 5828 2688 5892 2692
rect 5908 2748 5972 2752
rect 5908 2692 5912 2748
rect 5912 2692 5968 2748
rect 5968 2692 5972 2748
rect 5908 2688 5972 2692
rect 5988 2748 6052 2752
rect 5988 2692 5992 2748
rect 5992 2692 6048 2748
rect 6048 2692 6052 2748
rect 5988 2688 6052 2692
rect 6068 2748 6132 2752
rect 6068 2692 6072 2748
rect 6072 2692 6128 2748
rect 6128 2692 6132 2748
rect 6068 2688 6132 2692
rect 8542 2748 8606 2752
rect 8542 2692 8546 2748
rect 8546 2692 8602 2748
rect 8602 2692 8606 2748
rect 8542 2688 8606 2692
rect 8622 2748 8686 2752
rect 8622 2692 8626 2748
rect 8626 2692 8682 2748
rect 8682 2692 8686 2748
rect 8622 2688 8686 2692
rect 8702 2748 8766 2752
rect 8702 2692 8706 2748
rect 8706 2692 8762 2748
rect 8762 2692 8766 2748
rect 8702 2688 8766 2692
rect 8782 2748 8846 2752
rect 8782 2692 8786 2748
rect 8786 2692 8842 2748
rect 8842 2692 8846 2748
rect 8782 2688 8846 2692
rect 11256 2748 11320 2752
rect 11256 2692 11260 2748
rect 11260 2692 11316 2748
rect 11316 2692 11320 2748
rect 11256 2688 11320 2692
rect 11336 2748 11400 2752
rect 11336 2692 11340 2748
rect 11340 2692 11396 2748
rect 11396 2692 11400 2748
rect 11336 2688 11400 2692
rect 11416 2748 11480 2752
rect 11416 2692 11420 2748
rect 11420 2692 11476 2748
rect 11476 2692 11480 2748
rect 11416 2688 11480 2692
rect 11496 2748 11560 2752
rect 11496 2692 11500 2748
rect 11500 2692 11556 2748
rect 11556 2692 11560 2748
rect 11496 2688 11560 2692
rect 1757 2204 1821 2208
rect 1757 2148 1761 2204
rect 1761 2148 1817 2204
rect 1817 2148 1821 2204
rect 1757 2144 1821 2148
rect 1837 2204 1901 2208
rect 1837 2148 1841 2204
rect 1841 2148 1897 2204
rect 1897 2148 1901 2204
rect 1837 2144 1901 2148
rect 1917 2204 1981 2208
rect 1917 2148 1921 2204
rect 1921 2148 1977 2204
rect 1977 2148 1981 2204
rect 1917 2144 1981 2148
rect 1997 2204 2061 2208
rect 1997 2148 2001 2204
rect 2001 2148 2057 2204
rect 2057 2148 2061 2204
rect 1997 2144 2061 2148
rect 4471 2204 4535 2208
rect 4471 2148 4475 2204
rect 4475 2148 4531 2204
rect 4531 2148 4535 2204
rect 4471 2144 4535 2148
rect 4551 2204 4615 2208
rect 4551 2148 4555 2204
rect 4555 2148 4611 2204
rect 4611 2148 4615 2204
rect 4551 2144 4615 2148
rect 4631 2204 4695 2208
rect 4631 2148 4635 2204
rect 4635 2148 4691 2204
rect 4691 2148 4695 2204
rect 4631 2144 4695 2148
rect 4711 2204 4775 2208
rect 4711 2148 4715 2204
rect 4715 2148 4771 2204
rect 4771 2148 4775 2204
rect 4711 2144 4775 2148
rect 7185 2204 7249 2208
rect 7185 2148 7189 2204
rect 7189 2148 7245 2204
rect 7245 2148 7249 2204
rect 7185 2144 7249 2148
rect 7265 2204 7329 2208
rect 7265 2148 7269 2204
rect 7269 2148 7325 2204
rect 7325 2148 7329 2204
rect 7265 2144 7329 2148
rect 7345 2204 7409 2208
rect 7345 2148 7349 2204
rect 7349 2148 7405 2204
rect 7405 2148 7409 2204
rect 7345 2144 7409 2148
rect 7425 2204 7489 2208
rect 7425 2148 7429 2204
rect 7429 2148 7485 2204
rect 7485 2148 7489 2204
rect 7425 2144 7489 2148
rect 9899 2204 9963 2208
rect 9899 2148 9903 2204
rect 9903 2148 9959 2204
rect 9959 2148 9963 2204
rect 9899 2144 9963 2148
rect 9979 2204 10043 2208
rect 9979 2148 9983 2204
rect 9983 2148 10039 2204
rect 10039 2148 10043 2204
rect 9979 2144 10043 2148
rect 10059 2204 10123 2208
rect 10059 2148 10063 2204
rect 10063 2148 10119 2204
rect 10119 2148 10123 2204
rect 10059 2144 10123 2148
rect 10139 2204 10203 2208
rect 10139 2148 10143 2204
rect 10143 2148 10199 2204
rect 10199 2148 10203 2204
rect 10139 2144 10203 2148
rect 3114 1660 3178 1664
rect 3114 1604 3118 1660
rect 3118 1604 3174 1660
rect 3174 1604 3178 1660
rect 3114 1600 3178 1604
rect 3194 1660 3258 1664
rect 3194 1604 3198 1660
rect 3198 1604 3254 1660
rect 3254 1604 3258 1660
rect 3194 1600 3258 1604
rect 3274 1660 3338 1664
rect 3274 1604 3278 1660
rect 3278 1604 3334 1660
rect 3334 1604 3338 1660
rect 3274 1600 3338 1604
rect 3354 1660 3418 1664
rect 3354 1604 3358 1660
rect 3358 1604 3414 1660
rect 3414 1604 3418 1660
rect 3354 1600 3418 1604
rect 5828 1660 5892 1664
rect 5828 1604 5832 1660
rect 5832 1604 5888 1660
rect 5888 1604 5892 1660
rect 5828 1600 5892 1604
rect 5908 1660 5972 1664
rect 5908 1604 5912 1660
rect 5912 1604 5968 1660
rect 5968 1604 5972 1660
rect 5908 1600 5972 1604
rect 5988 1660 6052 1664
rect 5988 1604 5992 1660
rect 5992 1604 6048 1660
rect 6048 1604 6052 1660
rect 5988 1600 6052 1604
rect 6068 1660 6132 1664
rect 6068 1604 6072 1660
rect 6072 1604 6128 1660
rect 6128 1604 6132 1660
rect 6068 1600 6132 1604
rect 8542 1660 8606 1664
rect 8542 1604 8546 1660
rect 8546 1604 8602 1660
rect 8602 1604 8606 1660
rect 8542 1600 8606 1604
rect 8622 1660 8686 1664
rect 8622 1604 8626 1660
rect 8626 1604 8682 1660
rect 8682 1604 8686 1660
rect 8622 1600 8686 1604
rect 8702 1660 8766 1664
rect 8702 1604 8706 1660
rect 8706 1604 8762 1660
rect 8762 1604 8766 1660
rect 8702 1600 8766 1604
rect 8782 1660 8846 1664
rect 8782 1604 8786 1660
rect 8786 1604 8842 1660
rect 8842 1604 8846 1660
rect 8782 1600 8846 1604
rect 11256 1660 11320 1664
rect 11256 1604 11260 1660
rect 11260 1604 11316 1660
rect 11316 1604 11320 1660
rect 11256 1600 11320 1604
rect 11336 1660 11400 1664
rect 11336 1604 11340 1660
rect 11340 1604 11396 1660
rect 11396 1604 11400 1660
rect 11336 1600 11400 1604
rect 11416 1660 11480 1664
rect 11416 1604 11420 1660
rect 11420 1604 11476 1660
rect 11476 1604 11480 1660
rect 11416 1600 11480 1604
rect 11496 1660 11560 1664
rect 11496 1604 11500 1660
rect 11500 1604 11556 1660
rect 11556 1604 11560 1660
rect 11496 1600 11560 1604
rect 1757 1116 1821 1120
rect 1757 1060 1761 1116
rect 1761 1060 1817 1116
rect 1817 1060 1821 1116
rect 1757 1056 1821 1060
rect 1837 1116 1901 1120
rect 1837 1060 1841 1116
rect 1841 1060 1897 1116
rect 1897 1060 1901 1116
rect 1837 1056 1901 1060
rect 1917 1116 1981 1120
rect 1917 1060 1921 1116
rect 1921 1060 1977 1116
rect 1977 1060 1981 1116
rect 1917 1056 1981 1060
rect 1997 1116 2061 1120
rect 1997 1060 2001 1116
rect 2001 1060 2057 1116
rect 2057 1060 2061 1116
rect 1997 1056 2061 1060
rect 4471 1116 4535 1120
rect 4471 1060 4475 1116
rect 4475 1060 4531 1116
rect 4531 1060 4535 1116
rect 4471 1056 4535 1060
rect 4551 1116 4615 1120
rect 4551 1060 4555 1116
rect 4555 1060 4611 1116
rect 4611 1060 4615 1116
rect 4551 1056 4615 1060
rect 4631 1116 4695 1120
rect 4631 1060 4635 1116
rect 4635 1060 4691 1116
rect 4691 1060 4695 1116
rect 4631 1056 4695 1060
rect 4711 1116 4775 1120
rect 4711 1060 4715 1116
rect 4715 1060 4771 1116
rect 4771 1060 4775 1116
rect 4711 1056 4775 1060
rect 7185 1116 7249 1120
rect 7185 1060 7189 1116
rect 7189 1060 7245 1116
rect 7245 1060 7249 1116
rect 7185 1056 7249 1060
rect 7265 1116 7329 1120
rect 7265 1060 7269 1116
rect 7269 1060 7325 1116
rect 7325 1060 7329 1116
rect 7265 1056 7329 1060
rect 7345 1116 7409 1120
rect 7345 1060 7349 1116
rect 7349 1060 7405 1116
rect 7405 1060 7409 1116
rect 7345 1056 7409 1060
rect 7425 1116 7489 1120
rect 7425 1060 7429 1116
rect 7429 1060 7485 1116
rect 7485 1060 7489 1116
rect 7425 1056 7489 1060
rect 9899 1116 9963 1120
rect 9899 1060 9903 1116
rect 9903 1060 9959 1116
rect 9959 1060 9963 1116
rect 9899 1056 9963 1060
rect 9979 1116 10043 1120
rect 9979 1060 9983 1116
rect 9983 1060 10039 1116
rect 10039 1060 10043 1116
rect 9979 1056 10043 1060
rect 10059 1116 10123 1120
rect 10059 1060 10063 1116
rect 10063 1060 10119 1116
rect 10119 1060 10123 1116
rect 10059 1056 10123 1060
rect 10139 1116 10203 1120
rect 10139 1060 10143 1116
rect 10143 1060 10199 1116
rect 10199 1060 10203 1116
rect 10139 1056 10203 1060
rect 3114 572 3178 576
rect 3114 516 3118 572
rect 3118 516 3174 572
rect 3174 516 3178 572
rect 3114 512 3178 516
rect 3194 572 3258 576
rect 3194 516 3198 572
rect 3198 516 3254 572
rect 3254 516 3258 572
rect 3194 512 3258 516
rect 3274 572 3338 576
rect 3274 516 3278 572
rect 3278 516 3334 572
rect 3334 516 3338 572
rect 3274 512 3338 516
rect 3354 572 3418 576
rect 3354 516 3358 572
rect 3358 516 3414 572
rect 3414 516 3418 572
rect 3354 512 3418 516
rect 5828 572 5892 576
rect 5828 516 5832 572
rect 5832 516 5888 572
rect 5888 516 5892 572
rect 5828 512 5892 516
rect 5908 572 5972 576
rect 5908 516 5912 572
rect 5912 516 5968 572
rect 5968 516 5972 572
rect 5908 512 5972 516
rect 5988 572 6052 576
rect 5988 516 5992 572
rect 5992 516 6048 572
rect 6048 516 6052 572
rect 5988 512 6052 516
rect 6068 572 6132 576
rect 6068 516 6072 572
rect 6072 516 6128 572
rect 6128 516 6132 572
rect 6068 512 6132 516
rect 8542 572 8606 576
rect 8542 516 8546 572
rect 8546 516 8602 572
rect 8602 516 8606 572
rect 8542 512 8606 516
rect 8622 572 8686 576
rect 8622 516 8626 572
rect 8626 516 8682 572
rect 8682 516 8686 572
rect 8622 512 8686 516
rect 8702 572 8766 576
rect 8702 516 8706 572
rect 8706 516 8762 572
rect 8762 516 8766 572
rect 8702 512 8766 516
rect 8782 572 8846 576
rect 8782 516 8786 572
rect 8786 516 8842 572
rect 8842 516 8846 572
rect 8782 512 8846 516
rect 11256 572 11320 576
rect 11256 516 11260 572
rect 11260 516 11316 572
rect 11316 516 11320 572
rect 11256 512 11320 516
rect 11336 572 11400 576
rect 11336 516 11340 572
rect 11340 516 11396 572
rect 11396 516 11400 572
rect 11336 512 11400 516
rect 11416 572 11480 576
rect 11416 516 11420 572
rect 11420 516 11476 572
rect 11476 516 11480 572
rect 11416 512 11480 516
rect 11496 572 11560 576
rect 11496 516 11500 572
rect 11500 516 11556 572
rect 11556 516 11560 572
rect 11496 512 11560 516
<< metal4 >>
rect 1749 10912 2069 11472
rect 1749 10848 1757 10912
rect 1821 10848 1837 10912
rect 1901 10848 1917 10912
rect 1981 10848 1997 10912
rect 2061 10848 2069 10912
rect 1749 9824 2069 10848
rect 1749 9760 1757 9824
rect 1821 9760 1837 9824
rect 1901 9760 1917 9824
rect 1981 9760 1997 9824
rect 2061 9760 2069 9824
rect 1749 8736 2069 9760
rect 1749 8672 1757 8736
rect 1821 8672 1837 8736
rect 1901 8672 1917 8736
rect 1981 8672 1997 8736
rect 2061 8672 2069 8736
rect 1749 7648 2069 8672
rect 1749 7584 1757 7648
rect 1821 7584 1837 7648
rect 1901 7584 1917 7648
rect 1981 7584 1997 7648
rect 2061 7584 2069 7648
rect 1749 6560 2069 7584
rect 1749 6496 1757 6560
rect 1821 6496 1837 6560
rect 1901 6496 1917 6560
rect 1981 6496 1997 6560
rect 2061 6496 2069 6560
rect 1749 5472 2069 6496
rect 1749 5408 1757 5472
rect 1821 5408 1837 5472
rect 1901 5408 1917 5472
rect 1981 5408 1997 5472
rect 2061 5408 2069 5472
rect 1749 4384 2069 5408
rect 1749 4320 1757 4384
rect 1821 4320 1837 4384
rect 1901 4320 1917 4384
rect 1981 4320 1997 4384
rect 2061 4320 2069 4384
rect 1749 3296 2069 4320
rect 1749 3232 1757 3296
rect 1821 3232 1837 3296
rect 1901 3232 1917 3296
rect 1981 3232 1997 3296
rect 2061 3232 2069 3296
rect 1749 2208 2069 3232
rect 1749 2144 1757 2208
rect 1821 2144 1837 2208
rect 1901 2144 1917 2208
rect 1981 2144 1997 2208
rect 2061 2144 2069 2208
rect 1749 1120 2069 2144
rect 1749 1056 1757 1120
rect 1821 1056 1837 1120
rect 1901 1056 1917 1120
rect 1981 1056 1997 1120
rect 2061 1056 2069 1120
rect 1749 496 2069 1056
rect 3106 11456 3426 11472
rect 3106 11392 3114 11456
rect 3178 11392 3194 11456
rect 3258 11392 3274 11456
rect 3338 11392 3354 11456
rect 3418 11392 3426 11456
rect 3106 10368 3426 11392
rect 3106 10304 3114 10368
rect 3178 10304 3194 10368
rect 3258 10304 3274 10368
rect 3338 10304 3354 10368
rect 3418 10304 3426 10368
rect 3106 9280 3426 10304
rect 3106 9216 3114 9280
rect 3178 9216 3194 9280
rect 3258 9216 3274 9280
rect 3338 9216 3354 9280
rect 3418 9216 3426 9280
rect 3106 8192 3426 9216
rect 3106 8128 3114 8192
rect 3178 8128 3194 8192
rect 3258 8128 3274 8192
rect 3338 8128 3354 8192
rect 3418 8128 3426 8192
rect 3106 7104 3426 8128
rect 3106 7040 3114 7104
rect 3178 7040 3194 7104
rect 3258 7040 3274 7104
rect 3338 7040 3354 7104
rect 3418 7040 3426 7104
rect 3106 6016 3426 7040
rect 3106 5952 3114 6016
rect 3178 5952 3194 6016
rect 3258 5952 3274 6016
rect 3338 5952 3354 6016
rect 3418 5952 3426 6016
rect 3106 4928 3426 5952
rect 3106 4864 3114 4928
rect 3178 4864 3194 4928
rect 3258 4864 3274 4928
rect 3338 4864 3354 4928
rect 3418 4864 3426 4928
rect 3106 3840 3426 4864
rect 3106 3776 3114 3840
rect 3178 3776 3194 3840
rect 3258 3776 3274 3840
rect 3338 3776 3354 3840
rect 3418 3776 3426 3840
rect 3106 2752 3426 3776
rect 3106 2688 3114 2752
rect 3178 2688 3194 2752
rect 3258 2688 3274 2752
rect 3338 2688 3354 2752
rect 3418 2688 3426 2752
rect 3106 1664 3426 2688
rect 3106 1600 3114 1664
rect 3178 1600 3194 1664
rect 3258 1600 3274 1664
rect 3338 1600 3354 1664
rect 3418 1600 3426 1664
rect 3106 576 3426 1600
rect 3106 512 3114 576
rect 3178 512 3194 576
rect 3258 512 3274 576
rect 3338 512 3354 576
rect 3418 512 3426 576
rect 3106 496 3426 512
rect 4463 10912 4783 11472
rect 4463 10848 4471 10912
rect 4535 10848 4551 10912
rect 4615 10848 4631 10912
rect 4695 10848 4711 10912
rect 4775 10848 4783 10912
rect 4463 9824 4783 10848
rect 4463 9760 4471 9824
rect 4535 9760 4551 9824
rect 4615 9760 4631 9824
rect 4695 9760 4711 9824
rect 4775 9760 4783 9824
rect 4463 8736 4783 9760
rect 4463 8672 4471 8736
rect 4535 8672 4551 8736
rect 4615 8672 4631 8736
rect 4695 8672 4711 8736
rect 4775 8672 4783 8736
rect 4463 7648 4783 8672
rect 4463 7584 4471 7648
rect 4535 7584 4551 7648
rect 4615 7584 4631 7648
rect 4695 7584 4711 7648
rect 4775 7584 4783 7648
rect 4463 6560 4783 7584
rect 4463 6496 4471 6560
rect 4535 6496 4551 6560
rect 4615 6496 4631 6560
rect 4695 6496 4711 6560
rect 4775 6496 4783 6560
rect 4463 5472 4783 6496
rect 4463 5408 4471 5472
rect 4535 5408 4551 5472
rect 4615 5408 4631 5472
rect 4695 5408 4711 5472
rect 4775 5408 4783 5472
rect 4463 4384 4783 5408
rect 4463 4320 4471 4384
rect 4535 4320 4551 4384
rect 4615 4320 4631 4384
rect 4695 4320 4711 4384
rect 4775 4320 4783 4384
rect 4463 3296 4783 4320
rect 4463 3232 4471 3296
rect 4535 3232 4551 3296
rect 4615 3232 4631 3296
rect 4695 3232 4711 3296
rect 4775 3232 4783 3296
rect 4463 2208 4783 3232
rect 4463 2144 4471 2208
rect 4535 2144 4551 2208
rect 4615 2144 4631 2208
rect 4695 2144 4711 2208
rect 4775 2144 4783 2208
rect 4463 1120 4783 2144
rect 4463 1056 4471 1120
rect 4535 1056 4551 1120
rect 4615 1056 4631 1120
rect 4695 1056 4711 1120
rect 4775 1056 4783 1120
rect 4463 496 4783 1056
rect 5820 11456 6140 11472
rect 5820 11392 5828 11456
rect 5892 11392 5908 11456
rect 5972 11392 5988 11456
rect 6052 11392 6068 11456
rect 6132 11392 6140 11456
rect 5820 10368 6140 11392
rect 5820 10304 5828 10368
rect 5892 10304 5908 10368
rect 5972 10304 5988 10368
rect 6052 10304 6068 10368
rect 6132 10304 6140 10368
rect 5820 9280 6140 10304
rect 5820 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5988 9280
rect 6052 9216 6068 9280
rect 6132 9216 6140 9280
rect 5820 8192 6140 9216
rect 5820 8128 5828 8192
rect 5892 8128 5908 8192
rect 5972 8128 5988 8192
rect 6052 8128 6068 8192
rect 6132 8128 6140 8192
rect 5820 7104 6140 8128
rect 5820 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5988 7104
rect 6052 7040 6068 7104
rect 6132 7040 6140 7104
rect 5820 6016 6140 7040
rect 5820 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5988 6016
rect 6052 5952 6068 6016
rect 6132 5952 6140 6016
rect 5820 4928 6140 5952
rect 5820 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5988 4928
rect 6052 4864 6068 4928
rect 6132 4864 6140 4928
rect 5820 3840 6140 4864
rect 5820 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5988 3840
rect 6052 3776 6068 3840
rect 6132 3776 6140 3840
rect 5820 2752 6140 3776
rect 5820 2688 5828 2752
rect 5892 2688 5908 2752
rect 5972 2688 5988 2752
rect 6052 2688 6068 2752
rect 6132 2688 6140 2752
rect 5820 1664 6140 2688
rect 5820 1600 5828 1664
rect 5892 1600 5908 1664
rect 5972 1600 5988 1664
rect 6052 1600 6068 1664
rect 6132 1600 6140 1664
rect 5820 576 6140 1600
rect 5820 512 5828 576
rect 5892 512 5908 576
rect 5972 512 5988 576
rect 6052 512 6068 576
rect 6132 512 6140 576
rect 5820 496 6140 512
rect 7177 10912 7497 11472
rect 7177 10848 7185 10912
rect 7249 10848 7265 10912
rect 7329 10848 7345 10912
rect 7409 10848 7425 10912
rect 7489 10848 7497 10912
rect 7177 9824 7497 10848
rect 7177 9760 7185 9824
rect 7249 9760 7265 9824
rect 7329 9760 7345 9824
rect 7409 9760 7425 9824
rect 7489 9760 7497 9824
rect 7177 8736 7497 9760
rect 7177 8672 7185 8736
rect 7249 8672 7265 8736
rect 7329 8672 7345 8736
rect 7409 8672 7425 8736
rect 7489 8672 7497 8736
rect 7177 7648 7497 8672
rect 7177 7584 7185 7648
rect 7249 7584 7265 7648
rect 7329 7584 7345 7648
rect 7409 7584 7425 7648
rect 7489 7584 7497 7648
rect 7177 6560 7497 7584
rect 7177 6496 7185 6560
rect 7249 6496 7265 6560
rect 7329 6496 7345 6560
rect 7409 6496 7425 6560
rect 7489 6496 7497 6560
rect 7177 5472 7497 6496
rect 7177 5408 7185 5472
rect 7249 5408 7265 5472
rect 7329 5408 7345 5472
rect 7409 5408 7425 5472
rect 7489 5408 7497 5472
rect 7177 4384 7497 5408
rect 7177 4320 7185 4384
rect 7249 4320 7265 4384
rect 7329 4320 7345 4384
rect 7409 4320 7425 4384
rect 7489 4320 7497 4384
rect 7177 3296 7497 4320
rect 7177 3232 7185 3296
rect 7249 3232 7265 3296
rect 7329 3232 7345 3296
rect 7409 3232 7425 3296
rect 7489 3232 7497 3296
rect 7177 2208 7497 3232
rect 7177 2144 7185 2208
rect 7249 2144 7265 2208
rect 7329 2144 7345 2208
rect 7409 2144 7425 2208
rect 7489 2144 7497 2208
rect 7177 1120 7497 2144
rect 7177 1056 7185 1120
rect 7249 1056 7265 1120
rect 7329 1056 7345 1120
rect 7409 1056 7425 1120
rect 7489 1056 7497 1120
rect 7177 496 7497 1056
rect 8534 11456 8854 11472
rect 8534 11392 8542 11456
rect 8606 11392 8622 11456
rect 8686 11392 8702 11456
rect 8766 11392 8782 11456
rect 8846 11392 8854 11456
rect 8534 10368 8854 11392
rect 8534 10304 8542 10368
rect 8606 10304 8622 10368
rect 8686 10304 8702 10368
rect 8766 10304 8782 10368
rect 8846 10304 8854 10368
rect 8534 9280 8854 10304
rect 8534 9216 8542 9280
rect 8606 9216 8622 9280
rect 8686 9216 8702 9280
rect 8766 9216 8782 9280
rect 8846 9216 8854 9280
rect 8534 8192 8854 9216
rect 8534 8128 8542 8192
rect 8606 8128 8622 8192
rect 8686 8128 8702 8192
rect 8766 8128 8782 8192
rect 8846 8128 8854 8192
rect 8534 7104 8854 8128
rect 8534 7040 8542 7104
rect 8606 7040 8622 7104
rect 8686 7040 8702 7104
rect 8766 7040 8782 7104
rect 8846 7040 8854 7104
rect 8534 6016 8854 7040
rect 8534 5952 8542 6016
rect 8606 5952 8622 6016
rect 8686 5952 8702 6016
rect 8766 5952 8782 6016
rect 8846 5952 8854 6016
rect 8534 4928 8854 5952
rect 8534 4864 8542 4928
rect 8606 4864 8622 4928
rect 8686 4864 8702 4928
rect 8766 4864 8782 4928
rect 8846 4864 8854 4928
rect 8534 3840 8854 4864
rect 8534 3776 8542 3840
rect 8606 3776 8622 3840
rect 8686 3776 8702 3840
rect 8766 3776 8782 3840
rect 8846 3776 8854 3840
rect 8534 2752 8854 3776
rect 8534 2688 8542 2752
rect 8606 2688 8622 2752
rect 8686 2688 8702 2752
rect 8766 2688 8782 2752
rect 8846 2688 8854 2752
rect 8534 1664 8854 2688
rect 8534 1600 8542 1664
rect 8606 1600 8622 1664
rect 8686 1600 8702 1664
rect 8766 1600 8782 1664
rect 8846 1600 8854 1664
rect 8534 576 8854 1600
rect 8534 512 8542 576
rect 8606 512 8622 576
rect 8686 512 8702 576
rect 8766 512 8782 576
rect 8846 512 8854 576
rect 8534 496 8854 512
rect 9891 10912 10211 11472
rect 9891 10848 9899 10912
rect 9963 10848 9979 10912
rect 10043 10848 10059 10912
rect 10123 10848 10139 10912
rect 10203 10848 10211 10912
rect 9891 9824 10211 10848
rect 9891 9760 9899 9824
rect 9963 9760 9979 9824
rect 10043 9760 10059 9824
rect 10123 9760 10139 9824
rect 10203 9760 10211 9824
rect 9891 8736 10211 9760
rect 9891 8672 9899 8736
rect 9963 8672 9979 8736
rect 10043 8672 10059 8736
rect 10123 8672 10139 8736
rect 10203 8672 10211 8736
rect 9891 7648 10211 8672
rect 9891 7584 9899 7648
rect 9963 7584 9979 7648
rect 10043 7584 10059 7648
rect 10123 7584 10139 7648
rect 10203 7584 10211 7648
rect 9891 6560 10211 7584
rect 9891 6496 9899 6560
rect 9963 6496 9979 6560
rect 10043 6496 10059 6560
rect 10123 6496 10139 6560
rect 10203 6496 10211 6560
rect 9891 5472 10211 6496
rect 9891 5408 9899 5472
rect 9963 5408 9979 5472
rect 10043 5408 10059 5472
rect 10123 5408 10139 5472
rect 10203 5408 10211 5472
rect 9891 4384 10211 5408
rect 9891 4320 9899 4384
rect 9963 4320 9979 4384
rect 10043 4320 10059 4384
rect 10123 4320 10139 4384
rect 10203 4320 10211 4384
rect 9891 3296 10211 4320
rect 9891 3232 9899 3296
rect 9963 3232 9979 3296
rect 10043 3232 10059 3296
rect 10123 3232 10139 3296
rect 10203 3232 10211 3296
rect 9891 2208 10211 3232
rect 9891 2144 9899 2208
rect 9963 2144 9979 2208
rect 10043 2144 10059 2208
rect 10123 2144 10139 2208
rect 10203 2144 10211 2208
rect 9891 1120 10211 2144
rect 9891 1056 9899 1120
rect 9963 1056 9979 1120
rect 10043 1056 10059 1120
rect 10123 1056 10139 1120
rect 10203 1056 10211 1120
rect 9891 496 10211 1056
rect 11248 11456 11568 11472
rect 11248 11392 11256 11456
rect 11320 11392 11336 11456
rect 11400 11392 11416 11456
rect 11480 11392 11496 11456
rect 11560 11392 11568 11456
rect 11248 10368 11568 11392
rect 11248 10304 11256 10368
rect 11320 10304 11336 10368
rect 11400 10304 11416 10368
rect 11480 10304 11496 10368
rect 11560 10304 11568 10368
rect 11248 9280 11568 10304
rect 11248 9216 11256 9280
rect 11320 9216 11336 9280
rect 11400 9216 11416 9280
rect 11480 9216 11496 9280
rect 11560 9216 11568 9280
rect 11248 8192 11568 9216
rect 11248 8128 11256 8192
rect 11320 8128 11336 8192
rect 11400 8128 11416 8192
rect 11480 8128 11496 8192
rect 11560 8128 11568 8192
rect 11248 7104 11568 8128
rect 11248 7040 11256 7104
rect 11320 7040 11336 7104
rect 11400 7040 11416 7104
rect 11480 7040 11496 7104
rect 11560 7040 11568 7104
rect 11248 6016 11568 7040
rect 11248 5952 11256 6016
rect 11320 5952 11336 6016
rect 11400 5952 11416 6016
rect 11480 5952 11496 6016
rect 11560 5952 11568 6016
rect 11248 4928 11568 5952
rect 11248 4864 11256 4928
rect 11320 4864 11336 4928
rect 11400 4864 11416 4928
rect 11480 4864 11496 4928
rect 11560 4864 11568 4928
rect 11248 3840 11568 4864
rect 11248 3776 11256 3840
rect 11320 3776 11336 3840
rect 11400 3776 11416 3840
rect 11480 3776 11496 3840
rect 11560 3776 11568 3840
rect 11248 2752 11568 3776
rect 11248 2688 11256 2752
rect 11320 2688 11336 2752
rect 11400 2688 11416 2752
rect 11480 2688 11496 2752
rect 11560 2688 11568 2752
rect 11248 1664 11568 2688
rect 11248 1600 11256 1664
rect 11320 1600 11336 1664
rect 11400 1600 11416 1664
rect 11480 1600 11496 1664
rect 11560 1600 11568 1664
rect 11248 576 11568 1600
rect 11248 512 11256 576
rect 11320 512 11336 576
rect 11400 512 11416 576
rect 11480 512 11496 576
rect 11560 512 11568 576
rect 11248 496 11568 512
use sky130_fd_sc_hd__inv_2  _12_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9108 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _13_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7268 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _14_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _16_
timestamp 1688980957
transform -1 0 4416 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _17_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4324 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _18_
timestamp 1688980957
transform 1 0 4416 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _19_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6624 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _20_
timestamp 1688980957
transform 1 0 6072 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _22_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _23__2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8188 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _23_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8924 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_4  _24_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8004 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _25_
timestamp 1688980957
transform 1 0 4692 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _26_
timestamp 1688980957
transform 1 0 4048 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _27_
timestamp 1688980957
transform -1 0 8464 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1688980957
transform -1 0 5060 0 1 544
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1688980957
transform 1 0 8372 0 1 544
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5060 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 5612 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_76
timestamp 1688980957
transform 1 0 7544 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_105
timestamp 1688980957
transform 1 0 10212 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 10764 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10948 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4140 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4876 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_61
timestamp 1688980957
transform 1 0 6164 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp 1688980957
transform 1 0 10948 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3220 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_37
timestamp 1688980957
transform 1 0 3956 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_64
timestamp 1688980957
transform 1 0 6440 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_72
timestamp 1688980957
transform 1 0 7176 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_76
timestamp 1688980957
transform 1 0 7544 0 1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_109
timestamp 1688980957
transform 1 0 10580 0 1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3036 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_33
timestamp 1688980957
transform 1 0 3588 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_57
timestamp 1688980957
transform 1 0 5796 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_91
timestamp 1688980957
transform 1 0 8924 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_103
timestamp 1688980957
transform 1 0 10028 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_113
timestamp 1688980957
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3220 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_37
timestamp 1688980957
transform 1 0 3956 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8372 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_89
timestamp 1688980957
transform 1 0 8740 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_93
timestamp 1688980957
transform 1 0 9108 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_105
timestamp 1688980957
transform 1 0 10212 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_113
timestamp 1688980957
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_57
timestamp 1688980957
transform 1 0 5796 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_86
timestamp 1688980957
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_98
timestamp 1688980957
transform 1 0 9568 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_106
timestamp 1688980957
transform 1 0 10304 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_113
timestamp 1688980957
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_109
timestamp 1688980957
transform 1 0 10580 0 1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1688980957
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_109
timestamp 1688980957
transform 1 0 10580 0 1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_113
timestamp 1688980957
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_109
timestamp 1688980957
transform 1 0 10580 0 1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10212 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_113
timestamp 1688980957
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 9476 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_109
timestamp 1688980957
transform 1 0 10580 0 1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10212 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1688980957
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8372 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_109
timestamp 1688980957
transform 1 0 10580 0 1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10212 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1688980957
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 7636 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 9476 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_109
timestamp 1688980957
transform 1 0 10580 0 1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8004 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10212 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_113
timestamp 1688980957
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1688980957
transform 1 0 6532 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 9476 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_109
timestamp 1688980957
transform 1 0 10580 0 1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3036 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_29
timestamp 1688980957
transform 1 0 3220 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_41
timestamp 1688980957
transform 1 0 4324 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_53
timestamp 1688980957
transform 1 0 5428 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 5796 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_81
timestamp 1688980957
transform 1 0 8004 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_85
timestamp 1688980957
transform 1 0 8372 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_97
timestamp 1688980957
transform 1 0 9476 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1688980957
transform 1 0 10580 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_113
timestamp 1688980957
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7544 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6532 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 5704 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 6624 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 10580 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 11408 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 11408 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 11408 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 11408 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 11408 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 11408 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 11408 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 11408 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 11408 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 11408 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 11408 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 11408 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 11408 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 11408 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 11408 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 11408 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 11408 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 11408 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 11408 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 11408 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 3128 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 8280 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
<< labels >>
flabel metal4 s 3106 496 3426 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5820 496 6140 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 8534 496 8854 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11248 496 11568 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1749 496 2069 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4463 496 4783 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7177 496 7497 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9891 496 10211 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 8168 400 8288 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 7746 0 7802 400 0 FreeSans 224 90 0 0 drive_bit[0]
port 3 nsew signal tristate
flabel metal2 s 18 0 74 400 0 FreeSans 224 90 0 0 drive_bit[1]
port 4 nsew signal tristate
flabel metal2 s 3882 11600 3938 12000 0 FreeSans 224 90 0 0 drive_bit[2]
port 5 nsew signal tristate
flabel metal2 s 11610 11600 11666 12000 0 FreeSans 224 90 0 0 drive_bit[3]
port 6 nsew signal tristate
flabel metal3 s 11600 3408 12000 3528 0 FreeSans 480 0 0 0 n_rst
port 7 nsew signal input
rlabel via1 6060 11424 6060 11424 0 VGND
rlabel metal1 5980 10880 5980 10880 0 VPWR
rlabel metal1 8694 2822 8694 2822 0 _00_
rlabel metal1 7038 850 7038 850 0 _01_
rlabel metal1 5106 1530 5106 1530 0 _02_
rlabel via1 4554 1955 4554 1955 0 _03_
rlabel metal1 8004 3162 8004 3162 0 _04_
rlabel metal1 5658 1394 5658 1394 0 _05_
rlabel metal1 4646 1938 4646 1938 0 _06_
rlabel metal1 4370 1870 4370 1870 0 _07_
rlabel metal1 5106 2278 5106 2278 0 _08_
rlabel metal1 5888 3366 5888 3366 0 _09_
rlabel metal1 6946 2958 6946 2958 0 _10_
rlabel metal1 5704 2958 5704 2958 0 clk
rlabel metal1 6716 714 6716 714 0 clknet_0_clk
rlabel metal1 3910 2958 3910 2958 0 clknet_1_0__leaf_clk
rlabel metal1 8694 3502 8694 3502 0 clknet_1_1__leaf_clk
rlabel metal1 6486 3468 6486 3468 0 drive_bit[0]
rlabel metal2 46 1078 46 1078 0 drive_bit[1]
rlabel metal1 5612 2822 5612 2822 0 drive_bit[2]
rlabel metal2 6854 3910 6854 3910 0 drive_bit[3]
rlabel metal1 10810 3536 10810 3536 0 n_rst
rlabel metal1 9844 2958 9844 2958 0 net1
rlabel metal1 8234 2822 8234 2822 0 net2
rlabel metal1 4830 1462 4830 1462 0 net3
rlabel metal1 7452 986 7452 986 0 net4
rlabel metal1 4554 1802 4554 1802 0 net5
rlabel metal2 5566 1802 5566 1802 0 net6
rlabel metal1 7130 2584 7130 2584 0 rst
<< properties >>
string FIXED_BBOX 0 0 12000 12000
<< end >>
