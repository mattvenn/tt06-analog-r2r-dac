Simulation of an R2R DAC with Verilator and d_cosim

* https://sourceforge.net/p/ngspice/ngspice/ci/master/tree/examples/xspice/verilator/

* The digital portion of the circuit is specified in compiled Verilog.
* list the inputs and outputs
adut [ clk n_rst ext_data d7 d6 d5 d4 d3 d2 d1 d0 load_divider ] [b7 b6 b5 b4 b3 b2 b1 b0] null dut
.model dut d_cosim simulation="./r2r_dac_control.so"

* connect the driver to the R2R dac
* had to edit spice exported by xschem to add the subckt and ends

.include "../xschem/r2r.spice" 

xr2r b1 b0 b2 b3 b5 out b4 b6 b7 r2r

**** End of the ADC and its subcircuits.  Begin test circuit ****

.param vcc=3.3
vcc vcc 0 {vcc}

* Digital clock signal

aclock 0 clk clock
.model clock d_osc cntl_array=[-1 1] freq_array=[1Meg 1Meg]

* reset signal

Vreset n_rst 0 PULSE 3 0 1n 20p 20p 1u 500u

.control
tran 100n 400u
plot out
.endc
.end
