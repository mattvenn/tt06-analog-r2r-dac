VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_mattvenn_r2r_dac
  CLASS BLOCK ;
  FOREIGN tt_um_mattvenn_r2r_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 411.130493 ;
    ANTENNADIFFAREA 131.494949 ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 0.000 2.500 225.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 0.000 50.500 225.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 67.825 213.525 67.995 213.715 ;
        RECT 69.205 213.525 69.375 213.715 ;
        RECT 74.725 213.525 74.895 213.715 ;
        RECT 80.240 213.575 80.360 213.685 ;
        RECT 81.165 213.525 81.335 213.715 ;
        RECT 86.685 213.525 86.855 213.715 ;
        RECT 92.205 213.525 92.375 213.715 ;
        RECT 94.045 213.525 94.215 213.715 ;
        RECT 99.565 213.525 99.735 213.715 ;
        RECT 105.085 213.525 105.255 213.715 ;
        RECT 106.925 213.525 107.095 213.715 ;
        RECT 112.445 213.525 112.615 213.715 ;
        RECT 117.965 213.525 118.135 213.715 ;
        RECT 119.815 213.570 119.975 213.680 ;
        RECT 121.645 213.525 121.815 213.715 ;
        RECT 67.685 212.715 69.055 213.525 ;
        RECT 69.065 212.715 74.575 213.525 ;
        RECT 74.585 212.715 80.095 213.525 ;
        RECT 80.575 212.655 81.005 213.440 ;
        RECT 81.025 212.715 86.535 213.525 ;
        RECT 86.545 212.715 92.055 213.525 ;
        RECT 92.065 212.715 93.435 213.525 ;
        RECT 93.455 212.655 93.885 213.440 ;
        RECT 93.905 212.715 99.415 213.525 ;
        RECT 99.425 212.715 104.935 213.525 ;
        RECT 104.945 212.715 106.315 213.525 ;
        RECT 106.335 212.655 106.765 213.440 ;
        RECT 106.785 212.715 112.295 213.525 ;
        RECT 112.305 212.715 117.815 213.525 ;
        RECT 117.825 212.715 119.195 213.525 ;
        RECT 119.215 212.655 119.645 213.440 ;
        RECT 120.585 212.715 121.955 213.525 ;
      LAYER nwell ;
        RECT 67.490 209.495 122.150 212.325 ;
      LAYER pwell ;
        RECT 67.685 208.295 69.055 209.105 ;
        RECT 69.065 208.295 74.575 209.105 ;
        RECT 74.585 208.295 80.095 209.105 ;
        RECT 80.575 208.380 81.005 209.165 ;
        RECT 81.025 208.295 86.535 209.105 ;
        RECT 86.545 208.295 92.055 209.105 ;
        RECT 92.065 208.295 97.575 209.105 ;
        RECT 97.585 208.295 103.095 209.105 ;
        RECT 103.105 208.295 105.855 209.105 ;
        RECT 106.335 208.380 106.765 209.165 ;
        RECT 106.785 208.295 112.295 209.105 ;
        RECT 112.305 208.295 117.815 209.105 ;
        RECT 117.825 208.295 120.575 209.105 ;
        RECT 120.585 208.295 121.955 209.105 ;
        RECT 67.825 208.085 67.995 208.295 ;
        RECT 69.205 208.085 69.375 208.295 ;
        RECT 74.725 208.085 74.895 208.295 ;
        RECT 80.245 208.245 80.415 208.275 ;
        RECT 80.240 208.135 80.415 208.245 ;
        RECT 80.245 208.085 80.415 208.135 ;
        RECT 81.165 208.105 81.335 208.295 ;
        RECT 85.765 208.085 85.935 208.275 ;
        RECT 86.685 208.105 86.855 208.295 ;
        RECT 91.285 208.085 91.455 208.275 ;
        RECT 92.205 208.105 92.375 208.295 ;
        RECT 93.120 208.135 93.240 208.245 ;
        RECT 94.045 208.085 94.215 208.275 ;
        RECT 97.725 208.105 97.895 208.295 ;
        RECT 99.565 208.085 99.735 208.275 ;
        RECT 103.245 208.105 103.415 208.295 ;
        RECT 105.085 208.085 105.255 208.275 ;
        RECT 106.000 208.135 106.120 208.245 ;
        RECT 106.925 208.105 107.095 208.295 ;
        RECT 110.605 208.085 110.775 208.275 ;
        RECT 112.445 208.105 112.615 208.295 ;
        RECT 116.125 208.085 116.295 208.275 ;
        RECT 117.965 208.105 118.135 208.295 ;
        RECT 118.880 208.135 119.000 208.245 ;
        RECT 119.815 208.130 119.975 208.240 ;
        RECT 121.645 208.085 121.815 208.295 ;
        RECT 67.685 207.275 69.055 208.085 ;
        RECT 69.065 207.275 74.575 208.085 ;
        RECT 74.585 207.275 80.095 208.085 ;
        RECT 80.105 207.275 85.615 208.085 ;
        RECT 85.625 207.275 91.135 208.085 ;
        RECT 91.145 207.275 92.975 208.085 ;
        RECT 93.455 207.215 93.885 208.000 ;
        RECT 93.905 207.275 99.415 208.085 ;
        RECT 99.425 207.275 104.935 208.085 ;
        RECT 104.945 207.275 110.455 208.085 ;
        RECT 110.465 207.275 115.975 208.085 ;
        RECT 115.985 207.275 118.735 208.085 ;
        RECT 119.215 207.215 119.645 208.000 ;
        RECT 120.585 207.275 121.955 208.085 ;
      LAYER nwell ;
        RECT 67.490 204.055 122.150 206.885 ;
      LAYER pwell ;
        RECT 67.685 202.855 69.055 203.665 ;
        RECT 69.065 202.855 74.575 203.665 ;
        RECT 74.585 202.855 80.095 203.665 ;
        RECT 80.575 202.940 81.005 203.725 ;
        RECT 81.025 202.855 86.535 203.665 ;
        RECT 86.545 202.855 92.055 203.665 ;
        RECT 92.065 202.855 97.575 203.665 ;
        RECT 97.585 202.855 103.095 203.665 ;
        RECT 103.105 202.855 105.855 203.665 ;
        RECT 106.335 202.940 106.765 203.725 ;
        RECT 106.785 202.855 112.295 203.665 ;
        RECT 112.305 202.855 117.815 203.665 ;
        RECT 117.825 202.855 120.575 203.665 ;
        RECT 120.585 202.855 121.955 203.665 ;
        RECT 67.825 202.645 67.995 202.855 ;
        RECT 69.205 202.645 69.375 202.855 ;
        RECT 74.725 202.645 74.895 202.855 ;
        RECT 80.245 202.805 80.415 202.835 ;
        RECT 80.240 202.695 80.415 202.805 ;
        RECT 80.245 202.645 80.415 202.695 ;
        RECT 81.165 202.665 81.335 202.855 ;
        RECT 85.765 202.645 85.935 202.835 ;
        RECT 86.685 202.665 86.855 202.855 ;
        RECT 91.285 202.645 91.455 202.835 ;
        RECT 92.205 202.665 92.375 202.855 ;
        RECT 93.120 202.695 93.240 202.805 ;
        RECT 94.045 202.645 94.215 202.835 ;
        RECT 97.725 202.665 97.895 202.855 ;
        RECT 99.565 202.645 99.735 202.835 ;
        RECT 103.245 202.665 103.415 202.855 ;
        RECT 105.085 202.645 105.255 202.835 ;
        RECT 106.000 202.695 106.120 202.805 ;
        RECT 106.925 202.665 107.095 202.855 ;
        RECT 110.605 202.645 110.775 202.835 ;
        RECT 112.445 202.665 112.615 202.855 ;
        RECT 116.125 202.645 116.295 202.835 ;
        RECT 117.965 202.665 118.135 202.855 ;
        RECT 118.880 202.695 119.000 202.805 ;
        RECT 119.815 202.690 119.975 202.800 ;
        RECT 121.645 202.645 121.815 202.855 ;
        RECT 67.685 201.835 69.055 202.645 ;
        RECT 69.065 201.835 74.575 202.645 ;
        RECT 74.585 201.835 80.095 202.645 ;
        RECT 80.105 201.835 85.615 202.645 ;
        RECT 85.625 201.835 91.135 202.645 ;
        RECT 91.145 201.835 92.975 202.645 ;
        RECT 93.455 201.775 93.885 202.560 ;
        RECT 93.905 201.835 99.415 202.645 ;
        RECT 99.425 201.835 104.935 202.645 ;
        RECT 104.945 201.835 110.455 202.645 ;
        RECT 110.465 201.835 115.975 202.645 ;
        RECT 115.985 201.835 118.735 202.645 ;
        RECT 119.215 201.775 119.645 202.560 ;
        RECT 120.585 201.835 121.955 202.645 ;
      LAYER nwell ;
        RECT 67.490 198.615 122.150 201.445 ;
      LAYER pwell ;
        RECT 67.685 197.415 69.055 198.225 ;
        RECT 69.065 197.415 74.575 198.225 ;
        RECT 74.585 197.415 80.095 198.225 ;
        RECT 80.575 197.500 81.005 198.285 ;
        RECT 81.025 197.415 86.535 198.225 ;
        RECT 86.545 197.415 92.055 198.225 ;
        RECT 92.065 197.415 97.575 198.225 ;
        RECT 97.585 197.415 103.095 198.225 ;
        RECT 103.105 197.415 105.855 198.225 ;
        RECT 106.335 197.500 106.765 198.285 ;
        RECT 106.785 197.415 112.295 198.225 ;
        RECT 112.305 197.415 117.815 198.225 ;
        RECT 117.825 197.415 120.575 198.225 ;
        RECT 120.585 197.415 121.955 198.225 ;
        RECT 67.825 197.205 67.995 197.415 ;
        RECT 69.205 197.205 69.375 197.415 ;
        RECT 74.725 197.205 74.895 197.415 ;
        RECT 80.245 197.365 80.415 197.395 ;
        RECT 80.240 197.255 80.415 197.365 ;
        RECT 80.245 197.205 80.415 197.255 ;
        RECT 81.165 197.225 81.335 197.415 ;
        RECT 85.765 197.205 85.935 197.395 ;
        RECT 86.685 197.225 86.855 197.415 ;
        RECT 91.285 197.205 91.455 197.395 ;
        RECT 92.205 197.225 92.375 197.415 ;
        RECT 93.120 197.255 93.240 197.365 ;
        RECT 94.045 197.205 94.215 197.395 ;
        RECT 97.725 197.225 97.895 197.415 ;
        RECT 99.565 197.205 99.735 197.395 ;
        RECT 103.245 197.225 103.415 197.415 ;
        RECT 105.085 197.205 105.255 197.395 ;
        RECT 106.000 197.255 106.120 197.365 ;
        RECT 106.925 197.225 107.095 197.415 ;
        RECT 110.605 197.205 110.775 197.395 ;
        RECT 112.445 197.225 112.615 197.415 ;
        RECT 116.125 197.205 116.295 197.395 ;
        RECT 117.965 197.225 118.135 197.415 ;
        RECT 118.880 197.255 119.000 197.365 ;
        RECT 119.815 197.250 119.975 197.360 ;
        RECT 121.645 197.205 121.815 197.415 ;
        RECT 67.685 196.395 69.055 197.205 ;
        RECT 69.065 196.395 74.575 197.205 ;
        RECT 74.585 196.395 80.095 197.205 ;
        RECT 80.105 196.395 85.615 197.205 ;
        RECT 85.625 196.395 91.135 197.205 ;
        RECT 91.145 196.395 92.975 197.205 ;
        RECT 93.455 196.335 93.885 197.120 ;
        RECT 93.905 196.395 99.415 197.205 ;
        RECT 99.425 196.395 104.935 197.205 ;
        RECT 104.945 196.395 110.455 197.205 ;
        RECT 110.465 196.395 115.975 197.205 ;
        RECT 115.985 196.395 118.735 197.205 ;
        RECT 119.215 196.335 119.645 197.120 ;
        RECT 120.585 196.395 121.955 197.205 ;
      LAYER nwell ;
        RECT 67.490 193.175 122.150 196.005 ;
      LAYER pwell ;
        RECT 67.685 191.975 69.055 192.785 ;
        RECT 69.065 191.975 74.575 192.785 ;
        RECT 74.585 191.975 80.095 192.785 ;
        RECT 80.575 192.060 81.005 192.845 ;
        RECT 81.025 191.975 86.535 192.785 ;
        RECT 86.545 191.975 92.055 192.785 ;
        RECT 92.065 191.975 97.575 192.785 ;
        RECT 97.585 191.975 103.095 192.785 ;
        RECT 103.105 191.975 105.855 192.785 ;
        RECT 106.335 192.060 106.765 192.845 ;
        RECT 106.785 191.975 112.295 192.785 ;
        RECT 112.305 191.975 117.815 192.785 ;
        RECT 117.825 191.975 120.575 192.785 ;
        RECT 120.585 191.975 121.955 192.785 ;
        RECT 67.825 191.765 67.995 191.975 ;
        RECT 69.205 191.765 69.375 191.975 ;
        RECT 74.725 191.765 74.895 191.975 ;
        RECT 80.245 191.925 80.415 191.955 ;
        RECT 80.240 191.815 80.415 191.925 ;
        RECT 80.245 191.765 80.415 191.815 ;
        RECT 81.165 191.785 81.335 191.975 ;
        RECT 85.765 191.765 85.935 191.955 ;
        RECT 86.685 191.785 86.855 191.975 ;
        RECT 91.285 191.765 91.455 191.955 ;
        RECT 92.205 191.785 92.375 191.975 ;
        RECT 93.120 191.815 93.240 191.925 ;
        RECT 94.045 191.765 94.215 191.955 ;
        RECT 97.725 191.785 97.895 191.975 ;
        RECT 99.565 191.765 99.735 191.955 ;
        RECT 103.245 191.785 103.415 191.975 ;
        RECT 105.085 191.765 105.255 191.955 ;
        RECT 106.000 191.815 106.120 191.925 ;
        RECT 106.925 191.785 107.095 191.975 ;
        RECT 110.605 191.765 110.775 191.955 ;
        RECT 112.445 191.785 112.615 191.975 ;
        RECT 116.125 191.765 116.295 191.955 ;
        RECT 117.965 191.785 118.135 191.975 ;
        RECT 118.880 191.815 119.000 191.925 ;
        RECT 119.815 191.810 119.975 191.920 ;
        RECT 121.645 191.765 121.815 191.975 ;
        RECT 67.685 190.955 69.055 191.765 ;
        RECT 69.065 190.955 74.575 191.765 ;
        RECT 74.585 190.955 80.095 191.765 ;
        RECT 80.105 190.955 85.615 191.765 ;
        RECT 85.625 190.955 91.135 191.765 ;
        RECT 91.145 190.955 92.975 191.765 ;
        RECT 93.455 190.895 93.885 191.680 ;
        RECT 93.905 190.955 99.415 191.765 ;
        RECT 99.425 190.955 104.935 191.765 ;
        RECT 104.945 190.955 110.455 191.765 ;
        RECT 110.465 190.955 115.975 191.765 ;
        RECT 115.985 190.955 118.735 191.765 ;
        RECT 119.215 190.895 119.645 191.680 ;
        RECT 120.585 190.955 121.955 191.765 ;
      LAYER nwell ;
        RECT 67.490 187.735 122.150 190.565 ;
      LAYER pwell ;
        RECT 67.685 186.535 69.055 187.345 ;
        RECT 69.065 186.535 74.575 187.345 ;
        RECT 74.585 186.535 80.095 187.345 ;
        RECT 80.575 186.620 81.005 187.405 ;
        RECT 81.025 186.535 86.535 187.345 ;
        RECT 86.545 186.535 92.055 187.345 ;
        RECT 92.065 186.535 97.575 187.345 ;
        RECT 97.585 186.535 103.095 187.345 ;
        RECT 103.105 186.535 105.855 187.345 ;
        RECT 106.335 186.620 106.765 187.405 ;
        RECT 106.785 186.535 112.295 187.345 ;
        RECT 112.305 186.535 117.815 187.345 ;
        RECT 117.825 186.535 120.575 187.345 ;
        RECT 120.585 186.535 121.955 187.345 ;
        RECT 67.825 186.325 67.995 186.535 ;
        RECT 69.205 186.325 69.375 186.535 ;
        RECT 74.725 186.325 74.895 186.535 ;
        RECT 80.245 186.485 80.415 186.515 ;
        RECT 80.240 186.375 80.415 186.485 ;
        RECT 80.245 186.325 80.415 186.375 ;
        RECT 81.165 186.345 81.335 186.535 ;
        RECT 85.765 186.325 85.935 186.515 ;
        RECT 86.685 186.345 86.855 186.535 ;
        RECT 91.285 186.325 91.455 186.515 ;
        RECT 92.205 186.345 92.375 186.535 ;
        RECT 93.120 186.375 93.240 186.485 ;
        RECT 94.045 186.325 94.215 186.515 ;
        RECT 97.725 186.345 97.895 186.535 ;
        RECT 99.565 186.325 99.735 186.515 ;
        RECT 103.245 186.345 103.415 186.535 ;
        RECT 105.085 186.325 105.255 186.515 ;
        RECT 106.000 186.375 106.120 186.485 ;
        RECT 106.925 186.345 107.095 186.535 ;
        RECT 110.605 186.325 110.775 186.515 ;
        RECT 112.445 186.345 112.615 186.535 ;
        RECT 116.125 186.325 116.295 186.515 ;
        RECT 117.965 186.345 118.135 186.535 ;
        RECT 118.880 186.375 119.000 186.485 ;
        RECT 119.815 186.370 119.975 186.480 ;
        RECT 121.645 186.325 121.815 186.535 ;
        RECT 67.685 185.515 69.055 186.325 ;
        RECT 69.065 185.515 74.575 186.325 ;
        RECT 74.585 185.515 80.095 186.325 ;
        RECT 80.105 185.515 85.615 186.325 ;
        RECT 85.625 185.515 91.135 186.325 ;
        RECT 91.145 185.515 92.975 186.325 ;
        RECT 93.455 185.455 93.885 186.240 ;
        RECT 93.905 185.515 99.415 186.325 ;
        RECT 99.425 185.515 104.935 186.325 ;
        RECT 104.945 185.515 110.455 186.325 ;
        RECT 110.465 185.515 115.975 186.325 ;
        RECT 115.985 185.515 118.735 186.325 ;
        RECT 119.215 185.455 119.645 186.240 ;
        RECT 120.585 185.515 121.955 186.325 ;
      LAYER nwell ;
        RECT 67.490 182.295 122.150 185.125 ;
      LAYER pwell ;
        RECT 67.685 181.095 69.055 181.905 ;
        RECT 69.065 181.095 74.575 181.905 ;
        RECT 74.585 181.095 80.095 181.905 ;
        RECT 80.575 181.180 81.005 181.965 ;
        RECT 81.025 181.095 86.535 181.905 ;
        RECT 86.545 181.095 92.055 181.905 ;
        RECT 92.065 181.095 97.575 181.905 ;
        RECT 97.585 181.095 103.095 181.905 ;
        RECT 103.105 181.095 105.855 181.905 ;
        RECT 106.335 181.180 106.765 181.965 ;
        RECT 106.785 181.095 112.295 181.905 ;
        RECT 112.305 181.095 117.815 181.905 ;
        RECT 117.825 181.095 120.575 181.905 ;
        RECT 120.585 181.095 121.955 181.905 ;
        RECT 67.825 180.885 67.995 181.095 ;
        RECT 69.205 180.885 69.375 181.095 ;
        RECT 74.725 180.885 74.895 181.095 ;
        RECT 80.245 181.045 80.415 181.075 ;
        RECT 80.240 180.935 80.415 181.045 ;
        RECT 80.245 180.885 80.415 180.935 ;
        RECT 81.165 180.905 81.335 181.095 ;
        RECT 85.765 180.885 85.935 181.075 ;
        RECT 86.685 180.905 86.855 181.095 ;
        RECT 91.285 180.885 91.455 181.075 ;
        RECT 92.205 180.905 92.375 181.095 ;
        RECT 93.120 180.935 93.240 181.045 ;
        RECT 94.045 180.885 94.215 181.075 ;
        RECT 97.725 180.905 97.895 181.095 ;
        RECT 99.565 180.885 99.735 181.075 ;
        RECT 103.245 180.905 103.415 181.095 ;
        RECT 105.085 180.885 105.255 181.075 ;
        RECT 106.000 180.935 106.120 181.045 ;
        RECT 106.925 180.905 107.095 181.095 ;
        RECT 110.605 180.885 110.775 181.075 ;
        RECT 112.445 180.905 112.615 181.095 ;
        RECT 116.125 180.885 116.295 181.075 ;
        RECT 117.965 180.905 118.135 181.095 ;
        RECT 118.880 180.935 119.000 181.045 ;
        RECT 119.815 180.930 119.975 181.040 ;
        RECT 121.645 180.885 121.815 181.095 ;
        RECT 67.685 180.075 69.055 180.885 ;
        RECT 69.065 180.075 74.575 180.885 ;
        RECT 74.585 180.075 80.095 180.885 ;
        RECT 80.105 180.075 85.615 180.885 ;
        RECT 85.625 180.075 91.135 180.885 ;
        RECT 91.145 180.075 92.975 180.885 ;
        RECT 93.455 180.015 93.885 180.800 ;
        RECT 93.905 180.075 99.415 180.885 ;
        RECT 99.425 180.075 104.935 180.885 ;
        RECT 104.945 180.075 110.455 180.885 ;
        RECT 110.465 180.075 115.975 180.885 ;
        RECT 115.985 180.075 118.735 180.885 ;
        RECT 119.215 180.015 119.645 180.800 ;
        RECT 120.585 180.075 121.955 180.885 ;
      LAYER nwell ;
        RECT 67.490 176.855 122.150 179.685 ;
      LAYER pwell ;
        RECT 67.685 175.655 69.055 176.465 ;
        RECT 69.065 175.655 74.575 176.465 ;
        RECT 74.585 175.655 80.095 176.465 ;
        RECT 80.575 175.740 81.005 176.525 ;
        RECT 81.025 175.655 86.535 176.465 ;
        RECT 86.545 175.655 92.055 176.465 ;
        RECT 92.065 175.655 97.575 176.465 ;
        RECT 97.585 175.655 103.095 176.465 ;
        RECT 103.105 175.655 105.855 176.465 ;
        RECT 106.335 175.740 106.765 176.525 ;
        RECT 106.785 175.655 112.295 176.465 ;
        RECT 112.305 175.655 117.815 176.465 ;
        RECT 117.825 175.655 120.575 176.465 ;
        RECT 120.585 175.655 121.955 176.465 ;
        RECT 67.825 175.445 67.995 175.655 ;
        RECT 69.205 175.445 69.375 175.655 ;
        RECT 74.725 175.445 74.895 175.655 ;
        RECT 80.245 175.605 80.415 175.635 ;
        RECT 80.240 175.495 80.415 175.605 ;
        RECT 80.245 175.445 80.415 175.495 ;
        RECT 81.165 175.465 81.335 175.655 ;
        RECT 85.765 175.445 85.935 175.635 ;
        RECT 86.685 175.465 86.855 175.655 ;
        RECT 91.285 175.445 91.455 175.635 ;
        RECT 92.205 175.465 92.375 175.655 ;
        RECT 93.120 175.495 93.240 175.605 ;
        RECT 94.045 175.445 94.215 175.635 ;
        RECT 95.430 175.445 95.600 175.635 ;
        RECT 97.725 175.465 97.895 175.655 ;
        RECT 103.245 175.465 103.415 175.655 ;
        RECT 106.000 175.495 106.120 175.605 ;
        RECT 106.925 175.445 107.095 175.655 ;
        RECT 107.385 175.445 107.555 175.635 ;
        RECT 112.445 175.465 112.615 175.655 ;
        RECT 112.905 175.445 113.075 175.635 ;
        RECT 116.585 175.445 116.755 175.635 ;
        RECT 117.965 175.465 118.135 175.655 ;
        RECT 118.885 175.445 119.055 175.635 ;
        RECT 119.815 175.490 119.975 175.600 ;
        RECT 121.645 175.445 121.815 175.655 ;
        RECT 67.685 174.635 69.055 175.445 ;
        RECT 69.065 174.635 74.575 175.445 ;
        RECT 74.585 174.635 80.095 175.445 ;
        RECT 80.105 174.635 85.615 175.445 ;
        RECT 85.625 174.635 91.135 175.445 ;
        RECT 91.145 174.635 92.975 175.445 ;
        RECT 93.455 174.575 93.885 175.360 ;
        RECT 93.905 174.635 95.275 175.445 ;
        RECT 95.285 174.535 98.205 175.445 ;
        RECT 98.535 174.765 107.235 175.445 ;
        RECT 98.535 174.535 101.240 174.765 ;
        RECT 102.780 174.545 103.690 174.765 ;
        RECT 107.245 174.635 112.755 175.445 ;
        RECT 112.765 174.635 116.435 175.445 ;
        RECT 116.445 174.635 117.815 175.445 ;
        RECT 117.825 174.665 119.195 175.445 ;
        RECT 119.215 174.575 119.645 175.360 ;
        RECT 120.585 174.635 121.955 175.445 ;
      LAYER nwell ;
        RECT 67.490 171.415 122.150 174.245 ;
      LAYER pwell ;
        RECT 67.685 170.215 69.055 171.025 ;
        RECT 69.065 170.215 74.575 171.025 ;
        RECT 74.585 170.215 80.095 171.025 ;
        RECT 80.575 170.300 81.005 171.085 ;
        RECT 81.025 170.215 84.695 171.025 ;
        RECT 88.710 170.895 89.620 171.115 ;
        RECT 91.160 170.895 93.865 171.125 ;
        RECT 85.165 170.215 93.865 170.895 ;
        RECT 93.905 170.215 103.010 170.895 ;
        RECT 103.105 170.215 104.475 170.995 ;
        RECT 106.335 170.300 106.765 171.085 ;
        RECT 106.785 170.215 108.615 171.025 ;
        RECT 109.095 170.215 110.445 171.125 ;
        RECT 110.465 170.215 115.975 171.025 ;
        RECT 115.985 170.215 119.655 171.025 ;
        RECT 120.585 170.215 121.955 171.025 ;
        RECT 67.825 170.005 67.995 170.215 ;
        RECT 69.205 170.005 69.375 170.215 ;
        RECT 74.725 170.005 74.895 170.215 ;
        RECT 80.245 170.165 80.415 170.195 ;
        RECT 80.240 170.055 80.415 170.165 ;
        RECT 80.245 170.005 80.415 170.055 ;
        RECT 81.165 170.025 81.335 170.215 ;
        RECT 83.000 170.055 83.120 170.165 ;
        RECT 84.840 170.055 84.960 170.165 ;
        RECT 85.305 170.025 85.475 170.215 ;
        RECT 86.220 170.005 86.390 170.195 ;
        RECT 67.685 169.195 69.055 170.005 ;
        RECT 69.065 169.195 74.575 170.005 ;
        RECT 74.585 169.195 80.095 170.005 ;
        RECT 80.105 169.195 82.855 170.005 ;
        RECT 83.615 169.095 86.535 170.005 ;
        RECT 86.690 169.975 86.860 170.195 ;
        RECT 93.125 170.005 93.295 170.195 ;
        RECT 94.045 170.165 94.215 170.215 ;
        RECT 94.040 170.055 94.215 170.165 ;
        RECT 94.045 170.025 94.215 170.055 ;
        RECT 97.725 170.005 97.895 170.195 ;
        RECT 98.190 170.005 98.360 170.195 ;
        RECT 103.245 170.025 103.415 170.215 ;
        RECT 105.545 170.025 105.715 170.195 ;
        RECT 106.000 170.055 106.120 170.165 ;
        RECT 106.925 170.025 107.095 170.215 ;
        RECT 108.760 170.055 108.880 170.165 ;
        RECT 109.225 170.005 109.395 170.195 ;
        RECT 109.685 170.005 109.855 170.195 ;
        RECT 110.145 170.025 110.315 170.215 ;
        RECT 110.605 170.025 110.775 170.215 ;
        RECT 115.205 170.005 115.375 170.195 ;
        RECT 116.125 170.025 116.295 170.215 ;
        RECT 118.880 170.055 119.000 170.165 ;
        RECT 119.815 170.050 119.975 170.170 ;
        RECT 121.645 170.005 121.815 170.215 ;
        RECT 88.820 169.975 89.755 170.005 ;
        RECT 86.690 169.775 89.755 169.975 ;
        RECT 86.545 169.295 89.755 169.775 ;
        RECT 86.545 169.095 87.475 169.295 ;
        RECT 88.805 169.095 89.755 169.295 ;
        RECT 89.860 169.325 93.325 170.005 ;
        RECT 89.860 169.095 90.780 169.325 ;
        RECT 93.455 169.135 93.885 169.920 ;
        RECT 94.460 169.325 97.925 170.005 ;
        RECT 94.460 169.095 95.380 169.325 ;
        RECT 98.045 169.095 100.335 170.005 ;
        RECT 100.345 169.325 109.535 170.005 ;
        RECT 100.345 169.095 101.265 169.325 ;
        RECT 104.095 169.105 105.025 169.325 ;
        RECT 109.545 169.195 115.055 170.005 ;
        RECT 115.065 169.195 118.735 170.005 ;
        RECT 119.215 169.135 119.645 169.920 ;
        RECT 120.585 169.195 121.955 170.005 ;
      LAYER nwell ;
        RECT 67.490 165.975 122.150 168.805 ;
      LAYER pwell ;
        RECT 67.685 164.775 69.055 165.585 ;
        RECT 69.065 164.775 74.575 165.585 ;
        RECT 74.585 164.775 80.095 165.585 ;
        RECT 80.575 164.860 81.005 165.645 ;
        RECT 81.025 164.775 84.695 165.585 ;
        RECT 85.165 164.775 86.980 165.685 ;
        RECT 87.005 164.775 88.355 165.685 ;
        RECT 91.930 165.455 92.840 165.675 ;
        RECT 94.380 165.455 97.085 165.685 ;
        RECT 88.385 164.775 97.085 165.455 ;
        RECT 97.125 164.775 100.795 165.585 ;
        RECT 101.265 164.775 102.635 165.555 ;
        RECT 102.645 164.775 106.315 165.585 ;
        RECT 106.335 164.860 106.765 165.645 ;
        RECT 106.785 164.775 112.295 165.585 ;
        RECT 112.305 164.775 117.815 165.585 ;
        RECT 117.825 164.775 120.575 165.585 ;
        RECT 120.585 164.775 121.955 165.585 ;
        RECT 67.825 164.565 67.995 164.775 ;
        RECT 69.205 164.565 69.375 164.775 ;
        RECT 74.725 164.565 74.895 164.775 ;
        RECT 80.245 164.725 80.415 164.755 ;
        RECT 80.240 164.615 80.415 164.725 ;
        RECT 80.245 164.565 80.415 164.615 ;
        RECT 81.165 164.585 81.335 164.775 ;
        RECT 84.840 164.615 84.960 164.725 ;
        RECT 85.765 164.565 85.935 164.755 ;
        RECT 86.685 164.585 86.855 164.775 ;
        RECT 87.150 164.585 87.320 164.775 ;
        RECT 88.525 164.585 88.695 164.775 ;
        RECT 89.445 164.565 89.615 164.755 ;
        RECT 90.825 164.565 90.995 164.755 ;
        RECT 94.045 164.565 94.215 164.755 ;
        RECT 95.880 164.615 96.000 164.725 ;
        RECT 97.265 164.585 97.435 164.775 ;
        RECT 100.940 164.615 101.060 164.725 ;
        RECT 102.315 164.585 102.485 164.775 ;
        RECT 102.785 164.585 102.955 164.775 ;
        RECT 104.625 164.565 104.795 164.755 ;
        RECT 105.085 164.565 105.255 164.755 ;
        RECT 106.925 164.585 107.095 164.775 ;
        RECT 110.605 164.565 110.775 164.755 ;
        RECT 112.445 164.585 112.615 164.775 ;
        RECT 116.125 164.565 116.295 164.755 ;
        RECT 117.965 164.585 118.135 164.775 ;
        RECT 118.880 164.615 119.000 164.725 ;
        RECT 119.815 164.610 119.975 164.720 ;
        RECT 121.645 164.565 121.815 164.775 ;
        RECT 67.685 163.755 69.055 164.565 ;
        RECT 69.065 163.755 74.575 164.565 ;
        RECT 74.585 163.755 80.095 164.565 ;
        RECT 80.105 163.755 85.615 164.565 ;
        RECT 85.625 163.755 89.295 164.565 ;
        RECT 89.305 163.755 90.675 164.565 ;
        RECT 90.685 163.655 93.435 164.565 ;
        RECT 93.455 163.695 93.885 164.480 ;
        RECT 93.920 163.655 95.735 164.565 ;
        RECT 96.235 163.885 104.935 164.565 ;
        RECT 96.235 163.655 98.940 163.885 ;
        RECT 100.480 163.665 101.390 163.885 ;
        RECT 104.945 163.755 110.455 164.565 ;
        RECT 110.465 163.755 115.975 164.565 ;
        RECT 115.985 163.755 118.735 164.565 ;
        RECT 119.215 163.695 119.645 164.480 ;
        RECT 120.585 163.755 121.955 164.565 ;
      LAYER nwell ;
        RECT 67.490 160.535 122.150 163.365 ;
      LAYER pwell ;
        RECT 67.685 159.335 69.055 160.145 ;
        RECT 69.065 159.335 74.575 160.145 ;
        RECT 74.585 159.335 80.095 160.145 ;
        RECT 80.575 159.420 81.005 160.205 ;
        RECT 81.110 159.335 90.215 160.015 ;
        RECT 90.225 159.335 92.975 160.145 ;
        RECT 93.455 159.420 93.885 160.205 ;
        RECT 93.905 159.335 97.575 160.145 ;
        RECT 100.240 160.015 101.160 160.245 ;
        RECT 97.695 159.335 101.160 160.015 ;
        RECT 101.265 159.335 102.615 160.245 ;
        RECT 102.645 159.335 106.315 160.145 ;
        RECT 106.335 159.420 106.765 160.205 ;
        RECT 106.785 159.335 115.890 160.015 ;
        RECT 115.985 159.335 118.735 160.145 ;
        RECT 119.215 159.420 119.645 160.205 ;
        RECT 120.585 159.335 121.955 160.145 ;
        RECT 67.825 159.145 67.995 159.335 ;
        RECT 69.205 159.145 69.375 159.335 ;
        RECT 74.725 159.145 74.895 159.335 ;
        RECT 80.240 159.175 80.360 159.285 ;
        RECT 89.905 159.145 90.075 159.335 ;
        RECT 90.365 159.145 90.535 159.335 ;
        RECT 93.120 159.175 93.240 159.285 ;
        RECT 94.045 159.145 94.215 159.335 ;
        RECT 97.725 159.145 97.895 159.335 ;
        RECT 101.410 159.145 101.580 159.335 ;
        RECT 102.785 159.145 102.955 159.335 ;
        RECT 106.925 159.145 107.095 159.335 ;
        RECT 116.125 159.145 116.295 159.335 ;
        RECT 118.880 159.175 119.000 159.285 ;
        RECT 119.815 159.180 119.975 159.290 ;
        RECT 121.645 159.145 121.815 159.335 ;
      LAYER li1 ;
        RECT 67.680 213.545 121.960 213.715 ;
        RECT 67.765 212.795 68.975 213.545 ;
        RECT 69.145 213.000 74.490 213.545 ;
        RECT 74.665 213.000 80.010 213.545 ;
        RECT 67.765 212.255 68.285 212.795 ;
        RECT 68.455 212.085 68.975 212.625 ;
        RECT 70.730 212.170 71.070 213.000 ;
        RECT 67.765 210.995 68.975 212.085 ;
        RECT 72.550 211.430 72.900 212.680 ;
        RECT 76.250 212.170 76.590 213.000 ;
        RECT 80.645 212.820 80.935 213.545 ;
        RECT 81.105 213.000 86.450 213.545 ;
        RECT 86.625 213.000 91.970 213.545 ;
        RECT 78.070 211.430 78.420 212.680 ;
        RECT 82.690 212.170 83.030 213.000 ;
        RECT 69.145 210.995 74.490 211.430 ;
        RECT 74.665 210.995 80.010 211.430 ;
        RECT 80.645 210.995 80.935 212.160 ;
        RECT 84.510 211.430 84.860 212.680 ;
        RECT 88.210 212.170 88.550 213.000 ;
        RECT 92.145 212.795 93.355 213.545 ;
        RECT 93.525 212.820 93.815 213.545 ;
        RECT 93.985 213.000 99.330 213.545 ;
        RECT 99.505 213.000 104.850 213.545 ;
        RECT 90.030 211.430 90.380 212.680 ;
        RECT 92.145 212.255 92.665 212.795 ;
        RECT 92.835 212.085 93.355 212.625 ;
        RECT 95.570 212.170 95.910 213.000 ;
        RECT 81.105 210.995 86.450 211.430 ;
        RECT 86.625 210.995 91.970 211.430 ;
        RECT 92.145 210.995 93.355 212.085 ;
        RECT 93.525 210.995 93.815 212.160 ;
        RECT 97.390 211.430 97.740 212.680 ;
        RECT 101.090 212.170 101.430 213.000 ;
        RECT 105.025 212.795 106.235 213.545 ;
        RECT 106.405 212.820 106.695 213.545 ;
        RECT 106.865 213.000 112.210 213.545 ;
        RECT 112.385 213.000 117.730 213.545 ;
        RECT 102.910 211.430 103.260 212.680 ;
        RECT 105.025 212.255 105.545 212.795 ;
        RECT 105.715 212.085 106.235 212.625 ;
        RECT 108.450 212.170 108.790 213.000 ;
        RECT 93.985 210.995 99.330 211.430 ;
        RECT 99.505 210.995 104.850 211.430 ;
        RECT 105.025 210.995 106.235 212.085 ;
        RECT 106.405 210.995 106.695 212.160 ;
        RECT 110.270 211.430 110.620 212.680 ;
        RECT 113.970 212.170 114.310 213.000 ;
        RECT 117.905 212.795 119.115 213.545 ;
        RECT 119.285 212.820 119.575 213.545 ;
        RECT 120.665 212.795 121.875 213.545 ;
        RECT 115.790 211.430 116.140 212.680 ;
        RECT 117.905 212.255 118.425 212.795 ;
        RECT 118.595 212.085 119.115 212.625 ;
        RECT 106.865 210.995 112.210 211.430 ;
        RECT 112.385 210.995 117.730 211.430 ;
        RECT 117.905 210.995 119.115 212.085 ;
        RECT 119.285 210.995 119.575 212.160 ;
        RECT 120.665 212.085 121.185 212.625 ;
        RECT 121.355 212.255 121.875 212.795 ;
        RECT 120.665 210.995 121.875 212.085 ;
        RECT 67.680 210.825 121.960 210.995 ;
        RECT 67.765 209.735 68.975 210.825 ;
        RECT 69.145 210.390 74.490 210.825 ;
        RECT 74.665 210.390 80.010 210.825 ;
        RECT 67.765 209.025 68.285 209.565 ;
        RECT 68.455 209.195 68.975 209.735 ;
        RECT 67.765 208.275 68.975 209.025 ;
        RECT 70.730 208.820 71.070 209.650 ;
        RECT 72.550 209.140 72.900 210.390 ;
        RECT 76.250 208.820 76.590 209.650 ;
        RECT 78.070 209.140 78.420 210.390 ;
        RECT 80.645 209.660 80.935 210.825 ;
        RECT 81.105 210.390 86.450 210.825 ;
        RECT 86.625 210.390 91.970 210.825 ;
        RECT 92.145 210.390 97.490 210.825 ;
        RECT 97.665 210.390 103.010 210.825 ;
        RECT 69.145 208.275 74.490 208.820 ;
        RECT 74.665 208.275 80.010 208.820 ;
        RECT 80.645 208.275 80.935 209.000 ;
        RECT 82.690 208.820 83.030 209.650 ;
        RECT 84.510 209.140 84.860 210.390 ;
        RECT 88.210 208.820 88.550 209.650 ;
        RECT 90.030 209.140 90.380 210.390 ;
        RECT 93.730 208.820 94.070 209.650 ;
        RECT 95.550 209.140 95.900 210.390 ;
        RECT 99.250 208.820 99.590 209.650 ;
        RECT 101.070 209.140 101.420 210.390 ;
        RECT 103.185 209.735 105.775 210.825 ;
        RECT 103.185 209.045 104.395 209.565 ;
        RECT 104.565 209.215 105.775 209.735 ;
        RECT 106.405 209.660 106.695 210.825 ;
        RECT 106.865 210.390 112.210 210.825 ;
        RECT 112.385 210.390 117.730 210.825 ;
        RECT 81.105 208.275 86.450 208.820 ;
        RECT 86.625 208.275 91.970 208.820 ;
        RECT 92.145 208.275 97.490 208.820 ;
        RECT 97.665 208.275 103.010 208.820 ;
        RECT 103.185 208.275 105.775 209.045 ;
        RECT 106.405 208.275 106.695 209.000 ;
        RECT 108.450 208.820 108.790 209.650 ;
        RECT 110.270 209.140 110.620 210.390 ;
        RECT 113.970 208.820 114.310 209.650 ;
        RECT 115.790 209.140 116.140 210.390 ;
        RECT 117.905 209.735 120.495 210.825 ;
        RECT 117.905 209.045 119.115 209.565 ;
        RECT 119.285 209.215 120.495 209.735 ;
        RECT 120.665 209.735 121.875 210.825 ;
        RECT 120.665 209.195 121.185 209.735 ;
        RECT 106.865 208.275 112.210 208.820 ;
        RECT 112.385 208.275 117.730 208.820 ;
        RECT 117.905 208.275 120.495 209.045 ;
        RECT 121.355 209.025 121.875 209.565 ;
        RECT 120.665 208.275 121.875 209.025 ;
        RECT 67.680 208.105 121.960 208.275 ;
        RECT 67.765 207.355 68.975 208.105 ;
        RECT 69.145 207.560 74.490 208.105 ;
        RECT 74.665 207.560 80.010 208.105 ;
        RECT 80.185 207.560 85.530 208.105 ;
        RECT 85.705 207.560 91.050 208.105 ;
        RECT 67.765 206.815 68.285 207.355 ;
        RECT 68.455 206.645 68.975 207.185 ;
        RECT 70.730 206.730 71.070 207.560 ;
        RECT 67.765 205.555 68.975 206.645 ;
        RECT 72.550 205.990 72.900 207.240 ;
        RECT 76.250 206.730 76.590 207.560 ;
        RECT 78.070 205.990 78.420 207.240 ;
        RECT 81.770 206.730 82.110 207.560 ;
        RECT 83.590 205.990 83.940 207.240 ;
        RECT 87.290 206.730 87.630 207.560 ;
        RECT 91.225 207.335 92.895 208.105 ;
        RECT 93.525 207.380 93.815 208.105 ;
        RECT 93.985 207.560 99.330 208.105 ;
        RECT 99.505 207.560 104.850 208.105 ;
        RECT 105.025 207.560 110.370 208.105 ;
        RECT 110.545 207.560 115.890 208.105 ;
        RECT 89.110 205.990 89.460 207.240 ;
        RECT 91.225 206.815 91.975 207.335 ;
        RECT 92.145 206.645 92.895 207.165 ;
        RECT 95.570 206.730 95.910 207.560 ;
        RECT 69.145 205.555 74.490 205.990 ;
        RECT 74.665 205.555 80.010 205.990 ;
        RECT 80.185 205.555 85.530 205.990 ;
        RECT 85.705 205.555 91.050 205.990 ;
        RECT 91.225 205.555 92.895 206.645 ;
        RECT 93.525 205.555 93.815 206.720 ;
        RECT 97.390 205.990 97.740 207.240 ;
        RECT 101.090 206.730 101.430 207.560 ;
        RECT 102.910 205.990 103.260 207.240 ;
        RECT 106.610 206.730 106.950 207.560 ;
        RECT 108.430 205.990 108.780 207.240 ;
        RECT 112.130 206.730 112.470 207.560 ;
        RECT 116.065 207.335 118.655 208.105 ;
        RECT 119.285 207.380 119.575 208.105 ;
        RECT 120.665 207.355 121.875 208.105 ;
        RECT 113.950 205.990 114.300 207.240 ;
        RECT 116.065 206.815 117.275 207.335 ;
        RECT 117.445 206.645 118.655 207.165 ;
        RECT 93.985 205.555 99.330 205.990 ;
        RECT 99.505 205.555 104.850 205.990 ;
        RECT 105.025 205.555 110.370 205.990 ;
        RECT 110.545 205.555 115.890 205.990 ;
        RECT 116.065 205.555 118.655 206.645 ;
        RECT 119.285 205.555 119.575 206.720 ;
        RECT 120.665 206.645 121.185 207.185 ;
        RECT 121.355 206.815 121.875 207.355 ;
        RECT 120.665 205.555 121.875 206.645 ;
        RECT 67.680 205.385 121.960 205.555 ;
        RECT 67.765 204.295 68.975 205.385 ;
        RECT 69.145 204.950 74.490 205.385 ;
        RECT 74.665 204.950 80.010 205.385 ;
        RECT 67.765 203.585 68.285 204.125 ;
        RECT 68.455 203.755 68.975 204.295 ;
        RECT 67.765 202.835 68.975 203.585 ;
        RECT 70.730 203.380 71.070 204.210 ;
        RECT 72.550 203.700 72.900 204.950 ;
        RECT 76.250 203.380 76.590 204.210 ;
        RECT 78.070 203.700 78.420 204.950 ;
        RECT 80.645 204.220 80.935 205.385 ;
        RECT 81.105 204.950 86.450 205.385 ;
        RECT 86.625 204.950 91.970 205.385 ;
        RECT 92.145 204.950 97.490 205.385 ;
        RECT 97.665 204.950 103.010 205.385 ;
        RECT 69.145 202.835 74.490 203.380 ;
        RECT 74.665 202.835 80.010 203.380 ;
        RECT 80.645 202.835 80.935 203.560 ;
        RECT 82.690 203.380 83.030 204.210 ;
        RECT 84.510 203.700 84.860 204.950 ;
        RECT 88.210 203.380 88.550 204.210 ;
        RECT 90.030 203.700 90.380 204.950 ;
        RECT 93.730 203.380 94.070 204.210 ;
        RECT 95.550 203.700 95.900 204.950 ;
        RECT 99.250 203.380 99.590 204.210 ;
        RECT 101.070 203.700 101.420 204.950 ;
        RECT 103.185 204.295 105.775 205.385 ;
        RECT 103.185 203.605 104.395 204.125 ;
        RECT 104.565 203.775 105.775 204.295 ;
        RECT 106.405 204.220 106.695 205.385 ;
        RECT 106.865 204.950 112.210 205.385 ;
        RECT 112.385 204.950 117.730 205.385 ;
        RECT 81.105 202.835 86.450 203.380 ;
        RECT 86.625 202.835 91.970 203.380 ;
        RECT 92.145 202.835 97.490 203.380 ;
        RECT 97.665 202.835 103.010 203.380 ;
        RECT 103.185 202.835 105.775 203.605 ;
        RECT 106.405 202.835 106.695 203.560 ;
        RECT 108.450 203.380 108.790 204.210 ;
        RECT 110.270 203.700 110.620 204.950 ;
        RECT 113.970 203.380 114.310 204.210 ;
        RECT 115.790 203.700 116.140 204.950 ;
        RECT 117.905 204.295 120.495 205.385 ;
        RECT 117.905 203.605 119.115 204.125 ;
        RECT 119.285 203.775 120.495 204.295 ;
        RECT 120.665 204.295 121.875 205.385 ;
        RECT 120.665 203.755 121.185 204.295 ;
        RECT 106.865 202.835 112.210 203.380 ;
        RECT 112.385 202.835 117.730 203.380 ;
        RECT 117.905 202.835 120.495 203.605 ;
        RECT 121.355 203.585 121.875 204.125 ;
        RECT 120.665 202.835 121.875 203.585 ;
        RECT 67.680 202.665 121.960 202.835 ;
        RECT 67.765 201.915 68.975 202.665 ;
        RECT 69.145 202.120 74.490 202.665 ;
        RECT 74.665 202.120 80.010 202.665 ;
        RECT 80.185 202.120 85.530 202.665 ;
        RECT 85.705 202.120 91.050 202.665 ;
        RECT 67.765 201.375 68.285 201.915 ;
        RECT 68.455 201.205 68.975 201.745 ;
        RECT 70.730 201.290 71.070 202.120 ;
        RECT 67.765 200.115 68.975 201.205 ;
        RECT 72.550 200.550 72.900 201.800 ;
        RECT 76.250 201.290 76.590 202.120 ;
        RECT 78.070 200.550 78.420 201.800 ;
        RECT 81.770 201.290 82.110 202.120 ;
        RECT 83.590 200.550 83.940 201.800 ;
        RECT 87.290 201.290 87.630 202.120 ;
        RECT 91.225 201.895 92.895 202.665 ;
        RECT 93.525 201.940 93.815 202.665 ;
        RECT 93.985 202.120 99.330 202.665 ;
        RECT 99.505 202.120 104.850 202.665 ;
        RECT 105.025 202.120 110.370 202.665 ;
        RECT 110.545 202.120 115.890 202.665 ;
        RECT 89.110 200.550 89.460 201.800 ;
        RECT 91.225 201.375 91.975 201.895 ;
        RECT 92.145 201.205 92.895 201.725 ;
        RECT 95.570 201.290 95.910 202.120 ;
        RECT 69.145 200.115 74.490 200.550 ;
        RECT 74.665 200.115 80.010 200.550 ;
        RECT 80.185 200.115 85.530 200.550 ;
        RECT 85.705 200.115 91.050 200.550 ;
        RECT 91.225 200.115 92.895 201.205 ;
        RECT 93.525 200.115 93.815 201.280 ;
        RECT 97.390 200.550 97.740 201.800 ;
        RECT 101.090 201.290 101.430 202.120 ;
        RECT 102.910 200.550 103.260 201.800 ;
        RECT 106.610 201.290 106.950 202.120 ;
        RECT 108.430 200.550 108.780 201.800 ;
        RECT 112.130 201.290 112.470 202.120 ;
        RECT 116.065 201.895 118.655 202.665 ;
        RECT 119.285 201.940 119.575 202.665 ;
        RECT 120.665 201.915 121.875 202.665 ;
        RECT 113.950 200.550 114.300 201.800 ;
        RECT 116.065 201.375 117.275 201.895 ;
        RECT 117.445 201.205 118.655 201.725 ;
        RECT 93.985 200.115 99.330 200.550 ;
        RECT 99.505 200.115 104.850 200.550 ;
        RECT 105.025 200.115 110.370 200.550 ;
        RECT 110.545 200.115 115.890 200.550 ;
        RECT 116.065 200.115 118.655 201.205 ;
        RECT 119.285 200.115 119.575 201.280 ;
        RECT 120.665 201.205 121.185 201.745 ;
        RECT 121.355 201.375 121.875 201.915 ;
        RECT 120.665 200.115 121.875 201.205 ;
        RECT 67.680 199.945 121.960 200.115 ;
        RECT 67.765 198.855 68.975 199.945 ;
        RECT 69.145 199.510 74.490 199.945 ;
        RECT 74.665 199.510 80.010 199.945 ;
        RECT 67.765 198.145 68.285 198.685 ;
        RECT 68.455 198.315 68.975 198.855 ;
        RECT 67.765 197.395 68.975 198.145 ;
        RECT 70.730 197.940 71.070 198.770 ;
        RECT 72.550 198.260 72.900 199.510 ;
        RECT 76.250 197.940 76.590 198.770 ;
        RECT 78.070 198.260 78.420 199.510 ;
        RECT 80.645 198.780 80.935 199.945 ;
        RECT 81.105 199.510 86.450 199.945 ;
        RECT 86.625 199.510 91.970 199.945 ;
        RECT 92.145 199.510 97.490 199.945 ;
        RECT 97.665 199.510 103.010 199.945 ;
        RECT 69.145 197.395 74.490 197.940 ;
        RECT 74.665 197.395 80.010 197.940 ;
        RECT 80.645 197.395 80.935 198.120 ;
        RECT 82.690 197.940 83.030 198.770 ;
        RECT 84.510 198.260 84.860 199.510 ;
        RECT 88.210 197.940 88.550 198.770 ;
        RECT 90.030 198.260 90.380 199.510 ;
        RECT 93.730 197.940 94.070 198.770 ;
        RECT 95.550 198.260 95.900 199.510 ;
        RECT 99.250 197.940 99.590 198.770 ;
        RECT 101.070 198.260 101.420 199.510 ;
        RECT 103.185 198.855 105.775 199.945 ;
        RECT 103.185 198.165 104.395 198.685 ;
        RECT 104.565 198.335 105.775 198.855 ;
        RECT 106.405 198.780 106.695 199.945 ;
        RECT 106.865 199.510 112.210 199.945 ;
        RECT 112.385 199.510 117.730 199.945 ;
        RECT 81.105 197.395 86.450 197.940 ;
        RECT 86.625 197.395 91.970 197.940 ;
        RECT 92.145 197.395 97.490 197.940 ;
        RECT 97.665 197.395 103.010 197.940 ;
        RECT 103.185 197.395 105.775 198.165 ;
        RECT 106.405 197.395 106.695 198.120 ;
        RECT 108.450 197.940 108.790 198.770 ;
        RECT 110.270 198.260 110.620 199.510 ;
        RECT 113.970 197.940 114.310 198.770 ;
        RECT 115.790 198.260 116.140 199.510 ;
        RECT 117.905 198.855 120.495 199.945 ;
        RECT 117.905 198.165 119.115 198.685 ;
        RECT 119.285 198.335 120.495 198.855 ;
        RECT 120.665 198.855 121.875 199.945 ;
        RECT 120.665 198.315 121.185 198.855 ;
        RECT 106.865 197.395 112.210 197.940 ;
        RECT 112.385 197.395 117.730 197.940 ;
        RECT 117.905 197.395 120.495 198.165 ;
        RECT 121.355 198.145 121.875 198.685 ;
        RECT 120.665 197.395 121.875 198.145 ;
        RECT 67.680 197.225 121.960 197.395 ;
        RECT 67.765 196.475 68.975 197.225 ;
        RECT 69.145 196.680 74.490 197.225 ;
        RECT 74.665 196.680 80.010 197.225 ;
        RECT 80.185 196.680 85.530 197.225 ;
        RECT 85.705 196.680 91.050 197.225 ;
        RECT 67.765 195.935 68.285 196.475 ;
        RECT 68.455 195.765 68.975 196.305 ;
        RECT 70.730 195.850 71.070 196.680 ;
        RECT 67.765 194.675 68.975 195.765 ;
        RECT 72.550 195.110 72.900 196.360 ;
        RECT 76.250 195.850 76.590 196.680 ;
        RECT 78.070 195.110 78.420 196.360 ;
        RECT 81.770 195.850 82.110 196.680 ;
        RECT 83.590 195.110 83.940 196.360 ;
        RECT 87.290 195.850 87.630 196.680 ;
        RECT 91.225 196.455 92.895 197.225 ;
        RECT 93.525 196.500 93.815 197.225 ;
        RECT 93.985 196.680 99.330 197.225 ;
        RECT 99.505 196.680 104.850 197.225 ;
        RECT 105.025 196.680 110.370 197.225 ;
        RECT 110.545 196.680 115.890 197.225 ;
        RECT 89.110 195.110 89.460 196.360 ;
        RECT 91.225 195.935 91.975 196.455 ;
        RECT 92.145 195.765 92.895 196.285 ;
        RECT 95.570 195.850 95.910 196.680 ;
        RECT 69.145 194.675 74.490 195.110 ;
        RECT 74.665 194.675 80.010 195.110 ;
        RECT 80.185 194.675 85.530 195.110 ;
        RECT 85.705 194.675 91.050 195.110 ;
        RECT 91.225 194.675 92.895 195.765 ;
        RECT 93.525 194.675 93.815 195.840 ;
        RECT 97.390 195.110 97.740 196.360 ;
        RECT 101.090 195.850 101.430 196.680 ;
        RECT 102.910 195.110 103.260 196.360 ;
        RECT 106.610 195.850 106.950 196.680 ;
        RECT 108.430 195.110 108.780 196.360 ;
        RECT 112.130 195.850 112.470 196.680 ;
        RECT 116.065 196.455 118.655 197.225 ;
        RECT 119.285 196.500 119.575 197.225 ;
        RECT 120.665 196.475 121.875 197.225 ;
        RECT 113.950 195.110 114.300 196.360 ;
        RECT 116.065 195.935 117.275 196.455 ;
        RECT 117.445 195.765 118.655 196.285 ;
        RECT 93.985 194.675 99.330 195.110 ;
        RECT 99.505 194.675 104.850 195.110 ;
        RECT 105.025 194.675 110.370 195.110 ;
        RECT 110.545 194.675 115.890 195.110 ;
        RECT 116.065 194.675 118.655 195.765 ;
        RECT 119.285 194.675 119.575 195.840 ;
        RECT 120.665 195.765 121.185 196.305 ;
        RECT 121.355 195.935 121.875 196.475 ;
        RECT 120.665 194.675 121.875 195.765 ;
        RECT 67.680 194.505 121.960 194.675 ;
        RECT 67.765 193.415 68.975 194.505 ;
        RECT 69.145 194.070 74.490 194.505 ;
        RECT 74.665 194.070 80.010 194.505 ;
        RECT 67.765 192.705 68.285 193.245 ;
        RECT 68.455 192.875 68.975 193.415 ;
        RECT 67.765 191.955 68.975 192.705 ;
        RECT 70.730 192.500 71.070 193.330 ;
        RECT 72.550 192.820 72.900 194.070 ;
        RECT 76.250 192.500 76.590 193.330 ;
        RECT 78.070 192.820 78.420 194.070 ;
        RECT 80.645 193.340 80.935 194.505 ;
        RECT 81.105 194.070 86.450 194.505 ;
        RECT 86.625 194.070 91.970 194.505 ;
        RECT 92.145 194.070 97.490 194.505 ;
        RECT 97.665 194.070 103.010 194.505 ;
        RECT 69.145 191.955 74.490 192.500 ;
        RECT 74.665 191.955 80.010 192.500 ;
        RECT 80.645 191.955 80.935 192.680 ;
        RECT 82.690 192.500 83.030 193.330 ;
        RECT 84.510 192.820 84.860 194.070 ;
        RECT 88.210 192.500 88.550 193.330 ;
        RECT 90.030 192.820 90.380 194.070 ;
        RECT 93.730 192.500 94.070 193.330 ;
        RECT 95.550 192.820 95.900 194.070 ;
        RECT 99.250 192.500 99.590 193.330 ;
        RECT 101.070 192.820 101.420 194.070 ;
        RECT 103.185 193.415 105.775 194.505 ;
        RECT 103.185 192.725 104.395 193.245 ;
        RECT 104.565 192.895 105.775 193.415 ;
        RECT 106.405 193.340 106.695 194.505 ;
        RECT 106.865 194.070 112.210 194.505 ;
        RECT 112.385 194.070 117.730 194.505 ;
        RECT 81.105 191.955 86.450 192.500 ;
        RECT 86.625 191.955 91.970 192.500 ;
        RECT 92.145 191.955 97.490 192.500 ;
        RECT 97.665 191.955 103.010 192.500 ;
        RECT 103.185 191.955 105.775 192.725 ;
        RECT 106.405 191.955 106.695 192.680 ;
        RECT 108.450 192.500 108.790 193.330 ;
        RECT 110.270 192.820 110.620 194.070 ;
        RECT 113.970 192.500 114.310 193.330 ;
        RECT 115.790 192.820 116.140 194.070 ;
        RECT 117.905 193.415 120.495 194.505 ;
        RECT 117.905 192.725 119.115 193.245 ;
        RECT 119.285 192.895 120.495 193.415 ;
        RECT 120.665 193.415 121.875 194.505 ;
        RECT 120.665 192.875 121.185 193.415 ;
        RECT 106.865 191.955 112.210 192.500 ;
        RECT 112.385 191.955 117.730 192.500 ;
        RECT 117.905 191.955 120.495 192.725 ;
        RECT 121.355 192.705 121.875 193.245 ;
        RECT 120.665 191.955 121.875 192.705 ;
        RECT 67.680 191.785 121.960 191.955 ;
        RECT 67.765 191.035 68.975 191.785 ;
        RECT 69.145 191.240 74.490 191.785 ;
        RECT 74.665 191.240 80.010 191.785 ;
        RECT 80.185 191.240 85.530 191.785 ;
        RECT 85.705 191.240 91.050 191.785 ;
        RECT 67.765 190.495 68.285 191.035 ;
        RECT 68.455 190.325 68.975 190.865 ;
        RECT 70.730 190.410 71.070 191.240 ;
        RECT 67.765 189.235 68.975 190.325 ;
        RECT 72.550 189.670 72.900 190.920 ;
        RECT 76.250 190.410 76.590 191.240 ;
        RECT 78.070 189.670 78.420 190.920 ;
        RECT 81.770 190.410 82.110 191.240 ;
        RECT 83.590 189.670 83.940 190.920 ;
        RECT 87.290 190.410 87.630 191.240 ;
        RECT 91.225 191.015 92.895 191.785 ;
        RECT 93.525 191.060 93.815 191.785 ;
        RECT 93.985 191.240 99.330 191.785 ;
        RECT 99.505 191.240 104.850 191.785 ;
        RECT 105.025 191.240 110.370 191.785 ;
        RECT 110.545 191.240 115.890 191.785 ;
        RECT 89.110 189.670 89.460 190.920 ;
        RECT 91.225 190.495 91.975 191.015 ;
        RECT 92.145 190.325 92.895 190.845 ;
        RECT 95.570 190.410 95.910 191.240 ;
        RECT 69.145 189.235 74.490 189.670 ;
        RECT 74.665 189.235 80.010 189.670 ;
        RECT 80.185 189.235 85.530 189.670 ;
        RECT 85.705 189.235 91.050 189.670 ;
        RECT 91.225 189.235 92.895 190.325 ;
        RECT 93.525 189.235 93.815 190.400 ;
        RECT 97.390 189.670 97.740 190.920 ;
        RECT 101.090 190.410 101.430 191.240 ;
        RECT 102.910 189.670 103.260 190.920 ;
        RECT 106.610 190.410 106.950 191.240 ;
        RECT 108.430 189.670 108.780 190.920 ;
        RECT 112.130 190.410 112.470 191.240 ;
        RECT 116.065 191.015 118.655 191.785 ;
        RECT 119.285 191.060 119.575 191.785 ;
        RECT 120.665 191.035 121.875 191.785 ;
        RECT 113.950 189.670 114.300 190.920 ;
        RECT 116.065 190.495 117.275 191.015 ;
        RECT 117.445 190.325 118.655 190.845 ;
        RECT 93.985 189.235 99.330 189.670 ;
        RECT 99.505 189.235 104.850 189.670 ;
        RECT 105.025 189.235 110.370 189.670 ;
        RECT 110.545 189.235 115.890 189.670 ;
        RECT 116.065 189.235 118.655 190.325 ;
        RECT 119.285 189.235 119.575 190.400 ;
        RECT 120.665 190.325 121.185 190.865 ;
        RECT 121.355 190.495 121.875 191.035 ;
        RECT 120.665 189.235 121.875 190.325 ;
        RECT 67.680 189.065 121.960 189.235 ;
        RECT 67.765 187.975 68.975 189.065 ;
        RECT 69.145 188.630 74.490 189.065 ;
        RECT 74.665 188.630 80.010 189.065 ;
        RECT 67.765 187.265 68.285 187.805 ;
        RECT 68.455 187.435 68.975 187.975 ;
        RECT 67.765 186.515 68.975 187.265 ;
        RECT 70.730 187.060 71.070 187.890 ;
        RECT 72.550 187.380 72.900 188.630 ;
        RECT 76.250 187.060 76.590 187.890 ;
        RECT 78.070 187.380 78.420 188.630 ;
        RECT 80.645 187.900 80.935 189.065 ;
        RECT 81.105 188.630 86.450 189.065 ;
        RECT 86.625 188.630 91.970 189.065 ;
        RECT 92.145 188.630 97.490 189.065 ;
        RECT 97.665 188.630 103.010 189.065 ;
        RECT 69.145 186.515 74.490 187.060 ;
        RECT 74.665 186.515 80.010 187.060 ;
        RECT 80.645 186.515 80.935 187.240 ;
        RECT 82.690 187.060 83.030 187.890 ;
        RECT 84.510 187.380 84.860 188.630 ;
        RECT 88.210 187.060 88.550 187.890 ;
        RECT 90.030 187.380 90.380 188.630 ;
        RECT 93.730 187.060 94.070 187.890 ;
        RECT 95.550 187.380 95.900 188.630 ;
        RECT 99.250 187.060 99.590 187.890 ;
        RECT 101.070 187.380 101.420 188.630 ;
        RECT 103.185 187.975 105.775 189.065 ;
        RECT 103.185 187.285 104.395 187.805 ;
        RECT 104.565 187.455 105.775 187.975 ;
        RECT 106.405 187.900 106.695 189.065 ;
        RECT 106.865 188.630 112.210 189.065 ;
        RECT 112.385 188.630 117.730 189.065 ;
        RECT 81.105 186.515 86.450 187.060 ;
        RECT 86.625 186.515 91.970 187.060 ;
        RECT 92.145 186.515 97.490 187.060 ;
        RECT 97.665 186.515 103.010 187.060 ;
        RECT 103.185 186.515 105.775 187.285 ;
        RECT 106.405 186.515 106.695 187.240 ;
        RECT 108.450 187.060 108.790 187.890 ;
        RECT 110.270 187.380 110.620 188.630 ;
        RECT 113.970 187.060 114.310 187.890 ;
        RECT 115.790 187.380 116.140 188.630 ;
        RECT 117.905 187.975 120.495 189.065 ;
        RECT 117.905 187.285 119.115 187.805 ;
        RECT 119.285 187.455 120.495 187.975 ;
        RECT 120.665 187.975 121.875 189.065 ;
        RECT 120.665 187.435 121.185 187.975 ;
        RECT 106.865 186.515 112.210 187.060 ;
        RECT 112.385 186.515 117.730 187.060 ;
        RECT 117.905 186.515 120.495 187.285 ;
        RECT 121.355 187.265 121.875 187.805 ;
        RECT 120.665 186.515 121.875 187.265 ;
        RECT 67.680 186.345 121.960 186.515 ;
        RECT 67.765 185.595 68.975 186.345 ;
        RECT 69.145 185.800 74.490 186.345 ;
        RECT 74.665 185.800 80.010 186.345 ;
        RECT 80.185 185.800 85.530 186.345 ;
        RECT 85.705 185.800 91.050 186.345 ;
        RECT 67.765 185.055 68.285 185.595 ;
        RECT 68.455 184.885 68.975 185.425 ;
        RECT 70.730 184.970 71.070 185.800 ;
        RECT 67.765 183.795 68.975 184.885 ;
        RECT 72.550 184.230 72.900 185.480 ;
        RECT 76.250 184.970 76.590 185.800 ;
        RECT 78.070 184.230 78.420 185.480 ;
        RECT 81.770 184.970 82.110 185.800 ;
        RECT 83.590 184.230 83.940 185.480 ;
        RECT 87.290 184.970 87.630 185.800 ;
        RECT 91.225 185.575 92.895 186.345 ;
        RECT 93.525 185.620 93.815 186.345 ;
        RECT 93.985 185.800 99.330 186.345 ;
        RECT 99.505 185.800 104.850 186.345 ;
        RECT 105.025 185.800 110.370 186.345 ;
        RECT 110.545 185.800 115.890 186.345 ;
        RECT 89.110 184.230 89.460 185.480 ;
        RECT 91.225 185.055 91.975 185.575 ;
        RECT 92.145 184.885 92.895 185.405 ;
        RECT 95.570 184.970 95.910 185.800 ;
        RECT 69.145 183.795 74.490 184.230 ;
        RECT 74.665 183.795 80.010 184.230 ;
        RECT 80.185 183.795 85.530 184.230 ;
        RECT 85.705 183.795 91.050 184.230 ;
        RECT 91.225 183.795 92.895 184.885 ;
        RECT 93.525 183.795 93.815 184.960 ;
        RECT 97.390 184.230 97.740 185.480 ;
        RECT 101.090 184.970 101.430 185.800 ;
        RECT 102.910 184.230 103.260 185.480 ;
        RECT 106.610 184.970 106.950 185.800 ;
        RECT 108.430 184.230 108.780 185.480 ;
        RECT 112.130 184.970 112.470 185.800 ;
        RECT 116.065 185.575 118.655 186.345 ;
        RECT 119.285 185.620 119.575 186.345 ;
        RECT 120.665 185.595 121.875 186.345 ;
        RECT 113.950 184.230 114.300 185.480 ;
        RECT 116.065 185.055 117.275 185.575 ;
        RECT 117.445 184.885 118.655 185.405 ;
        RECT 93.985 183.795 99.330 184.230 ;
        RECT 99.505 183.795 104.850 184.230 ;
        RECT 105.025 183.795 110.370 184.230 ;
        RECT 110.545 183.795 115.890 184.230 ;
        RECT 116.065 183.795 118.655 184.885 ;
        RECT 119.285 183.795 119.575 184.960 ;
        RECT 120.665 184.885 121.185 185.425 ;
        RECT 121.355 185.055 121.875 185.595 ;
        RECT 120.665 183.795 121.875 184.885 ;
        RECT 67.680 183.625 121.960 183.795 ;
        RECT 67.765 182.535 68.975 183.625 ;
        RECT 69.145 183.190 74.490 183.625 ;
        RECT 74.665 183.190 80.010 183.625 ;
        RECT 67.765 181.825 68.285 182.365 ;
        RECT 68.455 181.995 68.975 182.535 ;
        RECT 67.765 181.075 68.975 181.825 ;
        RECT 70.730 181.620 71.070 182.450 ;
        RECT 72.550 181.940 72.900 183.190 ;
        RECT 76.250 181.620 76.590 182.450 ;
        RECT 78.070 181.940 78.420 183.190 ;
        RECT 80.645 182.460 80.935 183.625 ;
        RECT 81.105 183.190 86.450 183.625 ;
        RECT 86.625 183.190 91.970 183.625 ;
        RECT 92.145 183.190 97.490 183.625 ;
        RECT 97.665 183.190 103.010 183.625 ;
        RECT 69.145 181.075 74.490 181.620 ;
        RECT 74.665 181.075 80.010 181.620 ;
        RECT 80.645 181.075 80.935 181.800 ;
        RECT 82.690 181.620 83.030 182.450 ;
        RECT 84.510 181.940 84.860 183.190 ;
        RECT 88.210 181.620 88.550 182.450 ;
        RECT 90.030 181.940 90.380 183.190 ;
        RECT 93.730 181.620 94.070 182.450 ;
        RECT 95.550 181.940 95.900 183.190 ;
        RECT 99.250 181.620 99.590 182.450 ;
        RECT 101.070 181.940 101.420 183.190 ;
        RECT 103.185 182.535 105.775 183.625 ;
        RECT 103.185 181.845 104.395 182.365 ;
        RECT 104.565 182.015 105.775 182.535 ;
        RECT 106.405 182.460 106.695 183.625 ;
        RECT 106.865 183.190 112.210 183.625 ;
        RECT 112.385 183.190 117.730 183.625 ;
        RECT 81.105 181.075 86.450 181.620 ;
        RECT 86.625 181.075 91.970 181.620 ;
        RECT 92.145 181.075 97.490 181.620 ;
        RECT 97.665 181.075 103.010 181.620 ;
        RECT 103.185 181.075 105.775 181.845 ;
        RECT 106.405 181.075 106.695 181.800 ;
        RECT 108.450 181.620 108.790 182.450 ;
        RECT 110.270 181.940 110.620 183.190 ;
        RECT 113.970 181.620 114.310 182.450 ;
        RECT 115.790 181.940 116.140 183.190 ;
        RECT 117.905 182.535 120.495 183.625 ;
        RECT 117.905 181.845 119.115 182.365 ;
        RECT 119.285 182.015 120.495 182.535 ;
        RECT 120.665 182.535 121.875 183.625 ;
        RECT 120.665 181.995 121.185 182.535 ;
        RECT 106.865 181.075 112.210 181.620 ;
        RECT 112.385 181.075 117.730 181.620 ;
        RECT 117.905 181.075 120.495 181.845 ;
        RECT 121.355 181.825 121.875 182.365 ;
        RECT 120.665 181.075 121.875 181.825 ;
        RECT 67.680 180.905 121.960 181.075 ;
        RECT 67.765 180.155 68.975 180.905 ;
        RECT 69.145 180.360 74.490 180.905 ;
        RECT 74.665 180.360 80.010 180.905 ;
        RECT 80.185 180.360 85.530 180.905 ;
        RECT 85.705 180.360 91.050 180.905 ;
        RECT 67.765 179.615 68.285 180.155 ;
        RECT 68.455 179.445 68.975 179.985 ;
        RECT 70.730 179.530 71.070 180.360 ;
        RECT 67.765 178.355 68.975 179.445 ;
        RECT 72.550 178.790 72.900 180.040 ;
        RECT 76.250 179.530 76.590 180.360 ;
        RECT 78.070 178.790 78.420 180.040 ;
        RECT 81.770 179.530 82.110 180.360 ;
        RECT 83.590 178.790 83.940 180.040 ;
        RECT 87.290 179.530 87.630 180.360 ;
        RECT 91.225 180.135 92.895 180.905 ;
        RECT 93.525 180.180 93.815 180.905 ;
        RECT 93.985 180.360 99.330 180.905 ;
        RECT 99.505 180.360 104.850 180.905 ;
        RECT 105.025 180.360 110.370 180.905 ;
        RECT 110.545 180.360 115.890 180.905 ;
        RECT 89.110 178.790 89.460 180.040 ;
        RECT 91.225 179.615 91.975 180.135 ;
        RECT 92.145 179.445 92.895 179.965 ;
        RECT 95.570 179.530 95.910 180.360 ;
        RECT 69.145 178.355 74.490 178.790 ;
        RECT 74.665 178.355 80.010 178.790 ;
        RECT 80.185 178.355 85.530 178.790 ;
        RECT 85.705 178.355 91.050 178.790 ;
        RECT 91.225 178.355 92.895 179.445 ;
        RECT 93.525 178.355 93.815 179.520 ;
        RECT 97.390 178.790 97.740 180.040 ;
        RECT 101.090 179.530 101.430 180.360 ;
        RECT 102.910 178.790 103.260 180.040 ;
        RECT 106.610 179.530 106.950 180.360 ;
        RECT 108.430 178.790 108.780 180.040 ;
        RECT 112.130 179.530 112.470 180.360 ;
        RECT 116.065 180.135 118.655 180.905 ;
        RECT 119.285 180.180 119.575 180.905 ;
        RECT 120.665 180.155 121.875 180.905 ;
        RECT 113.950 178.790 114.300 180.040 ;
        RECT 116.065 179.615 117.275 180.135 ;
        RECT 117.445 179.445 118.655 179.965 ;
        RECT 93.985 178.355 99.330 178.790 ;
        RECT 99.505 178.355 104.850 178.790 ;
        RECT 105.025 178.355 110.370 178.790 ;
        RECT 110.545 178.355 115.890 178.790 ;
        RECT 116.065 178.355 118.655 179.445 ;
        RECT 119.285 178.355 119.575 179.520 ;
        RECT 120.665 179.445 121.185 179.985 ;
        RECT 121.355 179.615 121.875 180.155 ;
        RECT 120.665 178.355 121.875 179.445 ;
        RECT 67.680 178.185 121.960 178.355 ;
        RECT 67.765 177.095 68.975 178.185 ;
        RECT 69.145 177.750 74.490 178.185 ;
        RECT 74.665 177.750 80.010 178.185 ;
        RECT 67.765 176.385 68.285 176.925 ;
        RECT 68.455 176.555 68.975 177.095 ;
        RECT 67.765 175.635 68.975 176.385 ;
        RECT 70.730 176.180 71.070 177.010 ;
        RECT 72.550 176.500 72.900 177.750 ;
        RECT 76.250 176.180 76.590 177.010 ;
        RECT 78.070 176.500 78.420 177.750 ;
        RECT 80.645 177.020 80.935 178.185 ;
        RECT 81.105 177.750 86.450 178.185 ;
        RECT 86.625 177.750 91.970 178.185 ;
        RECT 92.145 177.750 97.490 178.185 ;
        RECT 97.665 177.750 103.010 178.185 ;
        RECT 69.145 175.635 74.490 176.180 ;
        RECT 74.665 175.635 80.010 176.180 ;
        RECT 80.645 175.635 80.935 176.360 ;
        RECT 82.690 176.180 83.030 177.010 ;
        RECT 84.510 176.500 84.860 177.750 ;
        RECT 88.210 176.180 88.550 177.010 ;
        RECT 90.030 176.500 90.380 177.750 ;
        RECT 93.730 176.180 94.070 177.010 ;
        RECT 95.550 176.500 95.900 177.750 ;
        RECT 99.250 176.180 99.590 177.010 ;
        RECT 101.070 176.500 101.420 177.750 ;
        RECT 103.185 177.095 105.775 178.185 ;
        RECT 103.185 176.405 104.395 176.925 ;
        RECT 104.565 176.575 105.775 177.095 ;
        RECT 106.405 177.020 106.695 178.185 ;
        RECT 106.865 177.750 112.210 178.185 ;
        RECT 112.385 177.750 117.730 178.185 ;
        RECT 81.105 175.635 86.450 176.180 ;
        RECT 86.625 175.635 91.970 176.180 ;
        RECT 92.145 175.635 97.490 176.180 ;
        RECT 97.665 175.635 103.010 176.180 ;
        RECT 103.185 175.635 105.775 176.405 ;
        RECT 106.405 175.635 106.695 176.360 ;
        RECT 108.450 176.180 108.790 177.010 ;
        RECT 110.270 176.500 110.620 177.750 ;
        RECT 113.970 176.180 114.310 177.010 ;
        RECT 115.790 176.500 116.140 177.750 ;
        RECT 117.905 177.095 120.495 178.185 ;
        RECT 117.905 176.405 119.115 176.925 ;
        RECT 119.285 176.575 120.495 177.095 ;
        RECT 120.665 177.095 121.875 178.185 ;
        RECT 120.665 176.555 121.185 177.095 ;
        RECT 106.865 175.635 112.210 176.180 ;
        RECT 112.385 175.635 117.730 176.180 ;
        RECT 117.905 175.635 120.495 176.405 ;
        RECT 121.355 176.385 121.875 176.925 ;
        RECT 120.665 175.635 121.875 176.385 ;
        RECT 67.680 175.465 121.960 175.635 ;
        RECT 67.765 174.715 68.975 175.465 ;
        RECT 69.145 174.920 74.490 175.465 ;
        RECT 74.665 174.920 80.010 175.465 ;
        RECT 80.185 174.920 85.530 175.465 ;
        RECT 85.705 174.920 91.050 175.465 ;
        RECT 67.765 174.175 68.285 174.715 ;
        RECT 68.455 174.005 68.975 174.545 ;
        RECT 70.730 174.090 71.070 174.920 ;
        RECT 67.765 172.915 68.975 174.005 ;
        RECT 72.550 173.350 72.900 174.600 ;
        RECT 76.250 174.090 76.590 174.920 ;
        RECT 78.070 173.350 78.420 174.600 ;
        RECT 81.770 174.090 82.110 174.920 ;
        RECT 83.590 173.350 83.940 174.600 ;
        RECT 87.290 174.090 87.630 174.920 ;
        RECT 91.225 174.695 92.895 175.465 ;
        RECT 93.525 174.740 93.815 175.465 ;
        RECT 93.985 174.715 95.195 175.465 ;
        RECT 95.375 174.740 95.705 175.250 ;
        RECT 95.875 175.065 96.205 175.465 ;
        RECT 97.255 174.895 97.585 175.235 ;
        RECT 97.755 175.065 98.085 175.465 ;
        RECT 98.725 174.990 98.895 175.465 ;
        RECT 89.110 173.350 89.460 174.600 ;
        RECT 91.225 174.175 91.975 174.695 ;
        RECT 92.145 174.005 92.895 174.525 ;
        RECT 93.985 174.175 94.505 174.715 ;
        RECT 69.145 172.915 74.490 173.350 ;
        RECT 74.665 172.915 80.010 173.350 ;
        RECT 80.185 172.915 85.530 173.350 ;
        RECT 85.705 172.915 91.050 173.350 ;
        RECT 91.225 172.915 92.895 174.005 ;
        RECT 93.525 172.915 93.815 174.080 ;
        RECT 94.675 174.005 95.195 174.545 ;
        RECT 93.985 172.915 95.195 174.005 ;
        RECT 95.375 173.975 95.565 174.740 ;
        RECT 95.875 174.725 98.240 174.895 ;
        RECT 99.065 174.820 99.400 175.245 ;
        RECT 99.575 174.990 99.745 175.465 ;
        RECT 99.920 174.820 100.255 175.245 ;
        RECT 100.445 174.985 100.615 175.465 ;
        RECT 95.875 174.555 96.045 174.725 ;
        RECT 95.735 174.225 96.045 174.555 ;
        RECT 96.215 174.225 96.520 174.555 ;
        RECT 95.375 173.125 95.705 173.975 ;
        RECT 95.875 172.915 96.125 174.055 ;
        RECT 96.305 173.895 96.520 174.225 ;
        RECT 96.695 173.895 96.980 174.555 ;
        RECT 97.175 173.895 97.440 174.555 ;
        RECT 97.655 173.895 97.900 174.555 ;
        RECT 98.070 173.725 98.240 174.725 ;
        RECT 98.585 174.650 100.255 174.820 ;
        RECT 100.790 174.815 101.150 175.255 ;
        RECT 101.445 174.935 101.615 175.465 ;
        RECT 101.930 175.015 102.600 175.185 ;
        RECT 102.830 175.015 103.290 175.185 ;
        RECT 98.585 174.085 98.830 174.650 ;
        RECT 100.650 174.645 101.150 174.815 ;
        RECT 100.650 174.475 100.820 174.645 ;
        RECT 101.930 174.475 102.100 175.015 ;
        RECT 99.000 174.305 100.820 174.475 ;
        RECT 101.010 174.305 102.100 174.475 ;
        RECT 98.585 173.915 100.255 174.085 ;
        RECT 96.315 173.555 97.605 173.725 ;
        RECT 96.315 173.135 96.565 173.555 ;
        RECT 96.795 172.915 97.125 173.385 ;
        RECT 97.355 173.135 97.605 173.555 ;
        RECT 97.785 173.555 98.240 173.725 ;
        RECT 97.785 173.125 98.115 173.555 ;
        RECT 98.730 172.915 98.900 173.745 ;
        RECT 99.070 173.155 99.400 173.915 ;
        RECT 99.570 172.915 99.740 173.745 ;
        RECT 99.920 173.155 100.255 173.915 ;
        RECT 100.650 174.050 100.820 174.305 ;
        RECT 100.650 173.880 101.760 174.050 ;
        RECT 100.900 173.720 101.760 173.880 ;
        RECT 100.435 172.915 100.615 173.695 ;
        RECT 100.900 173.095 101.070 173.720 ;
        RECT 101.535 172.915 101.750 173.415 ;
        RECT 101.930 173.385 102.100 174.305 ;
        RECT 102.400 174.515 102.950 174.845 ;
        RECT 103.120 174.785 103.290 175.015 ;
        RECT 103.470 174.965 103.840 175.465 ;
        RECT 104.090 175.015 104.840 175.185 ;
        RECT 105.020 175.015 105.350 175.185 ;
        RECT 102.400 173.975 102.590 174.515 ;
        RECT 103.120 174.485 103.920 174.785 ;
        RECT 102.270 173.645 102.590 173.975 ;
        RECT 102.760 173.585 102.950 174.305 ;
        RECT 103.120 173.415 103.290 174.485 ;
        RECT 103.750 174.455 103.920 174.485 ;
        RECT 103.460 174.235 103.630 174.305 ;
        RECT 104.090 174.235 104.260 175.015 ;
        RECT 104.430 174.515 105.010 174.845 ;
        RECT 103.460 174.065 104.260 174.235 ;
        RECT 103.460 173.975 103.970 174.065 ;
        RECT 101.930 173.215 102.815 173.385 ;
        RECT 103.040 173.085 103.290 173.415 ;
        RECT 103.460 172.915 103.630 173.715 ;
        RECT 103.800 173.360 103.970 173.975 ;
        RECT 104.140 173.540 104.580 173.895 ;
        RECT 104.770 173.645 105.010 174.515 ;
        RECT 105.180 173.485 105.350 175.015 ;
        RECT 105.535 175.005 105.785 175.465 ;
        RECT 105.520 173.885 105.800 174.485 ;
        RECT 103.800 173.190 104.870 173.360 ;
        RECT 105.115 173.110 105.350 173.485 ;
        RECT 105.535 172.915 105.800 173.375 ;
        RECT 106.000 173.085 106.225 175.205 ;
        RECT 106.395 175.085 106.725 175.465 ;
        RECT 106.895 174.915 107.065 175.205 ;
        RECT 107.325 174.920 112.670 175.465 ;
        RECT 106.400 174.745 107.065 174.915 ;
        RECT 106.400 173.755 106.630 174.745 ;
        RECT 106.800 173.925 107.150 174.575 ;
        RECT 108.910 174.090 109.250 174.920 ;
        RECT 112.845 174.695 116.355 175.465 ;
        RECT 116.525 174.715 117.735 175.465 ;
        RECT 117.905 174.790 118.165 175.295 ;
        RECT 118.345 175.085 118.675 175.465 ;
        RECT 118.855 174.915 119.025 175.295 ;
        RECT 106.400 173.585 107.065 173.755 ;
        RECT 106.395 172.915 106.725 173.415 ;
        RECT 106.895 173.085 107.065 173.585 ;
        RECT 110.730 173.350 111.080 174.600 ;
        RECT 112.845 174.175 114.495 174.695 ;
        RECT 114.665 174.005 116.355 174.525 ;
        RECT 116.525 174.175 117.045 174.715 ;
        RECT 117.215 174.005 117.735 174.545 ;
        RECT 107.325 172.915 112.670 173.350 ;
        RECT 112.845 172.915 116.355 174.005 ;
        RECT 116.525 172.915 117.735 174.005 ;
        RECT 117.905 173.990 118.075 174.790 ;
        RECT 118.360 174.745 119.025 174.915 ;
        RECT 118.360 174.490 118.530 174.745 ;
        RECT 119.285 174.740 119.575 175.465 ;
        RECT 120.665 174.715 121.875 175.465 ;
        RECT 118.245 174.160 118.530 174.490 ;
        RECT 118.765 174.195 119.095 174.565 ;
        RECT 118.360 174.015 118.530 174.160 ;
        RECT 117.905 173.085 118.175 173.990 ;
        RECT 118.360 173.845 119.025 174.015 ;
        RECT 118.345 172.915 118.675 173.675 ;
        RECT 118.855 173.085 119.025 173.845 ;
        RECT 119.285 172.915 119.575 174.080 ;
        RECT 120.665 174.005 121.185 174.545 ;
        RECT 121.355 174.175 121.875 174.715 ;
        RECT 120.665 172.915 121.875 174.005 ;
        RECT 67.680 172.745 121.960 172.915 ;
        RECT 67.765 171.655 68.975 172.745 ;
        RECT 69.145 172.310 74.490 172.745 ;
        RECT 74.665 172.310 80.010 172.745 ;
        RECT 67.765 170.945 68.285 171.485 ;
        RECT 68.455 171.115 68.975 171.655 ;
        RECT 67.765 170.195 68.975 170.945 ;
        RECT 70.730 170.740 71.070 171.570 ;
        RECT 72.550 171.060 72.900 172.310 ;
        RECT 76.250 170.740 76.590 171.570 ;
        RECT 78.070 171.060 78.420 172.310 ;
        RECT 80.645 171.580 80.935 172.745 ;
        RECT 81.105 171.655 84.615 172.745 ;
        RECT 85.335 172.075 85.505 172.575 ;
        RECT 85.675 172.245 86.005 172.745 ;
        RECT 85.335 171.905 86.000 172.075 ;
        RECT 81.105 170.965 82.755 171.485 ;
        RECT 82.925 171.135 84.615 171.655 ;
        RECT 85.250 171.085 85.600 171.735 ;
        RECT 69.145 170.195 74.490 170.740 ;
        RECT 74.665 170.195 80.010 170.740 ;
        RECT 80.645 170.195 80.935 170.920 ;
        RECT 81.105 170.195 84.615 170.965 ;
        RECT 85.770 170.915 86.000 171.905 ;
        RECT 85.335 170.745 86.000 170.915 ;
        RECT 85.335 170.455 85.505 170.745 ;
        RECT 85.675 170.195 86.005 170.575 ;
        RECT 86.175 170.455 86.400 172.575 ;
        RECT 86.600 172.285 86.865 172.745 ;
        RECT 87.050 172.175 87.285 172.550 ;
        RECT 87.530 172.300 88.600 172.470 ;
        RECT 86.600 171.175 86.880 171.775 ;
        RECT 86.615 170.195 86.865 170.655 ;
        RECT 87.050 170.645 87.220 172.175 ;
        RECT 87.390 171.145 87.630 172.015 ;
        RECT 87.820 171.765 88.260 172.120 ;
        RECT 88.430 171.685 88.600 172.300 ;
        RECT 88.770 171.945 88.940 172.745 ;
        RECT 89.110 172.245 89.360 172.575 ;
        RECT 89.585 172.275 90.470 172.445 ;
        RECT 88.430 171.595 88.940 171.685 ;
        RECT 88.140 171.425 88.940 171.595 ;
        RECT 87.390 170.815 87.970 171.145 ;
        RECT 88.140 170.645 88.310 171.425 ;
        RECT 88.770 171.355 88.940 171.425 ;
        RECT 88.480 171.175 88.650 171.205 ;
        RECT 89.110 171.175 89.280 172.245 ;
        RECT 89.450 171.355 89.640 172.075 ;
        RECT 89.810 171.685 90.130 172.015 ;
        RECT 88.480 170.875 89.280 171.175 ;
        RECT 89.810 171.145 90.000 171.685 ;
        RECT 87.050 170.475 87.380 170.645 ;
        RECT 87.560 170.475 88.310 170.645 ;
        RECT 88.560 170.195 88.930 170.695 ;
        RECT 89.110 170.645 89.280 170.875 ;
        RECT 89.450 170.815 90.000 171.145 ;
        RECT 90.300 171.355 90.470 172.275 ;
        RECT 90.650 172.245 90.865 172.745 ;
        RECT 91.330 171.940 91.500 172.565 ;
        RECT 91.785 171.965 91.965 172.745 ;
        RECT 90.640 171.780 91.500 171.940 ;
        RECT 90.640 171.610 91.750 171.780 ;
        RECT 91.580 171.355 91.750 171.610 ;
        RECT 92.145 171.745 92.480 172.505 ;
        RECT 92.660 171.915 92.830 172.745 ;
        RECT 93.000 171.745 93.330 172.505 ;
        RECT 93.500 171.915 93.670 172.745 ;
        RECT 93.995 171.935 94.290 172.745 ;
        RECT 92.145 171.575 93.815 171.745 ;
        RECT 90.300 171.185 91.390 171.355 ;
        RECT 91.580 171.185 93.400 171.355 ;
        RECT 90.300 170.645 90.470 171.185 ;
        RECT 91.580 171.015 91.750 171.185 ;
        RECT 91.250 170.845 91.750 171.015 ;
        RECT 93.570 171.010 93.815 171.575 ;
        RECT 94.470 171.435 94.715 172.575 ;
        RECT 94.890 171.935 95.150 172.745 ;
        RECT 95.750 172.740 102.025 172.745 ;
        RECT 95.330 171.435 95.580 172.570 ;
        RECT 95.750 171.945 96.010 172.740 ;
        RECT 96.180 171.845 96.440 172.570 ;
        RECT 96.610 172.015 96.870 172.740 ;
        RECT 97.040 171.845 97.300 172.570 ;
        RECT 97.470 172.015 97.730 172.740 ;
        RECT 97.900 171.845 98.160 172.570 ;
        RECT 98.330 172.015 98.590 172.740 ;
        RECT 98.760 171.845 99.020 172.570 ;
        RECT 99.190 172.015 99.435 172.740 ;
        RECT 99.605 171.845 99.865 172.570 ;
        RECT 100.050 172.015 100.295 172.740 ;
        RECT 100.465 171.845 100.725 172.570 ;
        RECT 100.910 172.015 101.155 172.740 ;
        RECT 101.325 171.845 101.585 172.570 ;
        RECT 101.770 172.015 102.025 172.740 ;
        RECT 96.180 171.830 101.585 171.845 ;
        RECT 102.195 171.830 102.485 172.570 ;
        RECT 102.655 172.000 102.925 172.745 ;
        RECT 96.180 171.605 102.925 171.830 ;
        RECT 103.275 171.815 103.445 172.575 ;
        RECT 103.625 171.985 103.955 172.745 ;
        RECT 103.275 171.645 103.940 171.815 ;
        RECT 104.125 171.670 104.395 172.575 ;
        RECT 89.110 170.475 89.570 170.645 ;
        RECT 89.800 170.475 90.470 170.645 ;
        RECT 90.785 170.195 90.955 170.725 ;
        RECT 91.250 170.405 91.610 170.845 ;
        RECT 92.145 170.840 93.815 171.010 ;
        RECT 93.985 170.875 94.300 171.435 ;
        RECT 94.470 171.185 101.590 171.435 ;
        RECT 91.785 170.195 91.955 170.675 ;
        RECT 92.145 170.415 92.480 170.840 ;
        RECT 92.655 170.195 92.825 170.670 ;
        RECT 93.000 170.415 93.335 170.840 ;
        RECT 93.505 170.195 93.675 170.670 ;
        RECT 93.985 170.195 94.290 170.705 ;
        RECT 94.470 170.375 94.720 171.185 ;
        RECT 94.890 170.195 95.150 170.720 ;
        RECT 95.330 170.375 95.580 171.185 ;
        RECT 101.760 171.015 102.925 171.605 ;
        RECT 103.770 171.500 103.940 171.645 ;
        RECT 103.205 171.095 103.535 171.465 ;
        RECT 103.770 171.170 104.055 171.500 ;
        RECT 96.180 170.845 102.925 171.015 ;
        RECT 103.770 170.915 103.940 171.170 ;
        RECT 95.750 170.195 96.010 170.755 ;
        RECT 96.180 170.390 96.440 170.845 ;
        RECT 96.610 170.195 96.870 170.675 ;
        RECT 97.040 170.390 97.300 170.845 ;
        RECT 97.470 170.195 97.730 170.675 ;
        RECT 97.900 170.390 98.160 170.845 ;
        RECT 98.330 170.195 98.575 170.675 ;
        RECT 98.745 170.390 99.020 170.845 ;
        RECT 99.190 170.195 99.435 170.675 ;
        RECT 99.605 170.390 99.865 170.845 ;
        RECT 100.045 170.195 100.295 170.675 ;
        RECT 100.465 170.390 100.725 170.845 ;
        RECT 100.905 170.195 101.155 170.675 ;
        RECT 101.325 170.390 101.585 170.845 ;
        RECT 101.765 170.195 102.025 170.675 ;
        RECT 102.195 170.390 102.455 170.845 ;
        RECT 103.275 170.745 103.940 170.915 ;
        RECT 104.225 170.870 104.395 171.670 ;
        RECT 104.565 171.025 105.085 172.575 ;
        RECT 105.255 172.020 105.585 172.745 ;
        RECT 102.625 170.195 102.925 170.675 ;
        RECT 103.275 170.365 103.445 170.745 ;
        RECT 103.625 170.195 103.955 170.575 ;
        RECT 104.135 170.365 104.395 170.870 ;
        RECT 104.745 170.195 105.085 170.855 ;
        RECT 105.255 170.365 105.775 171.850 ;
        RECT 106.405 171.580 106.695 172.745 ;
        RECT 106.865 171.655 108.535 172.745 ;
        RECT 106.865 170.965 107.615 171.485 ;
        RECT 107.785 171.135 108.535 171.655 ;
        RECT 109.225 171.605 109.435 172.745 ;
        RECT 109.605 171.595 109.935 172.575 ;
        RECT 110.105 171.605 110.335 172.745 ;
        RECT 110.545 172.310 115.890 172.745 ;
        RECT 106.405 170.195 106.695 170.920 ;
        RECT 106.865 170.195 108.535 170.965 ;
        RECT 109.225 170.195 109.435 171.015 ;
        RECT 109.605 170.995 109.855 171.595 ;
        RECT 110.025 171.185 110.355 171.435 ;
        RECT 109.605 170.365 109.935 170.995 ;
        RECT 110.105 170.195 110.335 171.015 ;
        RECT 112.130 170.740 112.470 171.570 ;
        RECT 113.950 171.060 114.300 172.310 ;
        RECT 116.065 171.655 119.575 172.745 ;
        RECT 116.065 170.965 117.715 171.485 ;
        RECT 117.885 171.135 119.575 171.655 ;
        RECT 120.665 171.655 121.875 172.745 ;
        RECT 120.665 171.115 121.185 171.655 ;
        RECT 110.545 170.195 115.890 170.740 ;
        RECT 116.065 170.195 119.575 170.965 ;
        RECT 121.355 170.945 121.875 171.485 ;
        RECT 120.665 170.195 121.875 170.945 ;
        RECT 67.680 170.025 121.960 170.195 ;
        RECT 67.765 169.275 68.975 170.025 ;
        RECT 69.145 169.480 74.490 170.025 ;
        RECT 74.665 169.480 80.010 170.025 ;
        RECT 67.765 168.735 68.285 169.275 ;
        RECT 68.455 168.565 68.975 169.105 ;
        RECT 70.730 168.650 71.070 169.480 ;
        RECT 67.765 167.475 68.975 168.565 ;
        RECT 72.550 167.910 72.900 169.160 ;
        RECT 76.250 168.650 76.590 169.480 ;
        RECT 80.185 169.255 82.775 170.025 ;
        RECT 83.735 169.625 84.065 170.025 ;
        RECT 84.235 169.455 84.565 169.795 ;
        RECT 85.615 169.625 85.945 170.025 ;
        RECT 83.580 169.285 85.945 169.455 ;
        RECT 86.115 169.300 86.445 169.810 ;
        RECT 78.070 167.910 78.420 169.160 ;
        RECT 80.185 168.735 81.395 169.255 ;
        RECT 81.565 168.565 82.775 169.085 ;
        RECT 69.145 167.475 74.490 167.910 ;
        RECT 74.665 167.475 80.010 167.910 ;
        RECT 80.185 167.475 82.775 168.565 ;
        RECT 83.580 168.285 83.750 169.285 ;
        RECT 85.775 169.115 85.945 169.285 ;
        RECT 83.920 168.455 84.165 169.115 ;
        RECT 84.380 168.455 84.645 169.115 ;
        RECT 84.840 168.455 85.125 169.115 ;
        RECT 85.300 168.785 85.605 169.115 ;
        RECT 85.775 168.785 86.085 169.115 ;
        RECT 85.300 168.455 85.515 168.785 ;
        RECT 83.580 168.115 84.035 168.285 ;
        RECT 83.705 167.685 84.035 168.115 ;
        RECT 84.215 168.115 85.505 168.285 ;
        RECT 84.215 167.695 84.465 168.115 ;
        RECT 84.695 167.475 85.025 167.945 ;
        RECT 85.255 167.695 85.505 168.115 ;
        RECT 85.695 167.475 85.945 168.615 ;
        RECT 86.255 168.535 86.445 169.300 ;
        RECT 86.625 169.205 86.885 170.025 ;
        RECT 87.055 169.205 87.385 169.625 ;
        RECT 87.565 169.540 88.355 169.805 ;
        RECT 87.135 169.115 87.385 169.205 ;
        RECT 86.115 167.685 86.445 168.535 ;
        RECT 86.625 168.155 86.965 169.035 ;
        RECT 87.135 168.865 87.930 169.115 ;
        RECT 86.625 167.475 86.885 167.985 ;
        RECT 87.135 167.645 87.305 168.865 ;
        RECT 88.100 168.685 88.355 169.540 ;
        RECT 88.525 169.385 88.725 169.805 ;
        RECT 88.915 169.565 89.245 170.025 ;
        RECT 88.525 168.865 88.935 169.385 ;
        RECT 89.415 169.375 89.675 169.855 ;
        RECT 89.105 168.685 89.335 169.115 ;
        RECT 87.545 168.515 89.335 168.685 ;
        RECT 87.545 168.150 87.795 168.515 ;
        RECT 87.965 168.155 88.295 168.345 ;
        RECT 88.515 168.220 89.230 168.515 ;
        RECT 89.505 168.345 89.675 169.375 ;
        RECT 87.965 167.980 88.160 168.155 ;
        RECT 87.545 167.475 88.160 167.980 ;
        RECT 88.330 167.645 88.805 167.985 ;
        RECT 88.975 167.475 89.190 168.020 ;
        RECT 89.400 167.645 89.675 168.345 ;
        RECT 89.845 169.285 90.230 169.855 ;
        RECT 90.400 169.565 90.725 170.025 ;
        RECT 91.245 169.395 91.525 169.855 ;
        RECT 89.845 168.615 90.125 169.285 ;
        RECT 90.400 169.225 91.525 169.395 ;
        RECT 90.400 169.115 90.850 169.225 ;
        RECT 90.295 168.785 90.850 169.115 ;
        RECT 91.715 169.055 92.115 169.855 ;
        RECT 92.515 169.565 92.785 170.025 ;
        RECT 92.955 169.395 93.240 169.855 ;
        RECT 89.845 167.645 90.230 168.615 ;
        RECT 90.400 168.325 90.850 168.785 ;
        RECT 91.020 168.495 92.115 169.055 ;
        RECT 90.400 168.105 91.525 168.325 ;
        RECT 90.400 167.475 90.725 167.935 ;
        RECT 91.245 167.645 91.525 168.105 ;
        RECT 91.715 167.645 92.115 168.495 ;
        RECT 92.285 169.225 93.240 169.395 ;
        RECT 93.525 169.300 93.815 170.025 ;
        RECT 94.445 169.285 94.830 169.855 ;
        RECT 95.000 169.565 95.325 170.025 ;
        RECT 95.845 169.395 96.125 169.855 ;
        RECT 92.285 168.325 92.495 169.225 ;
        RECT 92.665 168.495 93.355 169.055 ;
        RECT 92.285 168.105 93.240 168.325 ;
        RECT 92.515 167.475 92.785 167.935 ;
        RECT 92.955 167.645 93.240 168.105 ;
        RECT 93.525 167.475 93.815 168.640 ;
        RECT 94.445 168.615 94.725 169.285 ;
        RECT 95.000 169.225 96.125 169.395 ;
        RECT 95.000 169.115 95.450 169.225 ;
        RECT 94.895 168.785 95.450 169.115 ;
        RECT 96.315 169.055 96.715 169.855 ;
        RECT 97.115 169.565 97.385 170.025 ;
        RECT 97.555 169.395 97.840 169.855 ;
        RECT 94.445 167.645 94.830 168.615 ;
        RECT 95.000 168.325 95.450 168.785 ;
        RECT 95.620 168.495 96.715 169.055 ;
        RECT 95.000 168.105 96.125 168.325 ;
        RECT 95.000 167.475 95.325 167.935 ;
        RECT 95.845 167.645 96.125 168.105 ;
        RECT 96.315 167.645 96.715 168.495 ;
        RECT 96.885 169.225 97.840 169.395 ;
        RECT 98.130 169.285 98.465 170.025 ;
        RECT 96.885 168.325 97.095 169.225 ;
        RECT 98.635 169.115 98.850 169.810 ;
        RECT 99.040 169.285 99.390 169.810 ;
        RECT 99.560 169.285 100.255 169.855 ;
        RECT 100.430 169.315 100.685 169.845 ;
        RECT 100.855 169.565 101.160 170.025 ;
        RECT 101.405 169.645 102.475 169.815 ;
        RECT 99.185 169.115 99.390 169.285 ;
        RECT 97.265 168.495 97.955 169.055 ;
        RECT 98.150 168.785 98.435 169.115 ;
        RECT 98.635 168.785 99.015 169.115 ;
        RECT 99.185 168.785 99.495 169.115 ;
        RECT 99.665 168.615 99.835 169.285 ;
        RECT 96.885 168.105 97.840 168.325 ;
        RECT 97.115 167.475 97.385 167.935 ;
        RECT 97.555 167.645 97.840 168.105 ;
        RECT 98.125 167.475 98.385 168.615 ;
        RECT 98.555 168.445 99.835 168.615 ;
        RECT 100.015 168.445 100.255 169.115 ;
        RECT 100.430 168.665 100.640 169.315 ;
        RECT 101.405 169.290 101.725 169.645 ;
        RECT 101.400 169.115 101.725 169.290 ;
        RECT 100.810 168.815 101.725 169.115 ;
        RECT 101.895 169.075 102.135 169.475 ;
        RECT 102.305 169.415 102.475 169.645 ;
        RECT 102.645 169.585 102.835 170.025 ;
        RECT 103.005 169.575 103.955 169.855 ;
        RECT 104.175 169.665 104.525 169.835 ;
        RECT 102.305 169.245 102.835 169.415 ;
        RECT 100.810 168.785 101.550 168.815 ;
        RECT 98.555 167.645 98.885 168.445 ;
        RECT 99.055 167.475 99.225 168.275 ;
        RECT 99.425 167.645 99.755 168.445 ;
        RECT 99.955 167.475 100.235 168.275 ;
        RECT 100.430 167.785 100.685 168.665 ;
        RECT 100.855 167.475 101.160 168.615 ;
        RECT 101.380 168.195 101.550 168.785 ;
        RECT 101.895 168.705 102.435 169.075 ;
        RECT 102.615 168.965 102.835 169.245 ;
        RECT 103.005 168.795 103.175 169.575 ;
        RECT 102.770 168.625 103.175 168.795 ;
        RECT 103.345 168.785 103.695 169.405 ;
        RECT 102.770 168.535 102.940 168.625 ;
        RECT 103.865 168.615 104.075 169.405 ;
        RECT 101.720 168.365 102.940 168.535 ;
        RECT 103.400 168.455 104.075 168.615 ;
        RECT 101.380 168.025 102.180 168.195 ;
        RECT 101.500 167.475 101.830 167.855 ;
        RECT 102.010 167.735 102.180 168.025 ;
        RECT 102.770 167.985 102.940 168.365 ;
        RECT 103.110 168.445 104.075 168.455 ;
        RECT 104.265 169.275 104.525 169.665 ;
        RECT 104.735 169.565 105.065 170.025 ;
        RECT 105.940 169.635 106.795 169.805 ;
        RECT 107.000 169.635 107.495 169.805 ;
        RECT 107.665 169.665 107.995 170.025 ;
        RECT 104.265 168.585 104.435 169.275 ;
        RECT 104.605 168.925 104.775 169.105 ;
        RECT 104.945 169.095 105.735 169.345 ;
        RECT 105.940 168.925 106.110 169.635 ;
        RECT 106.280 169.125 106.635 169.345 ;
        RECT 104.605 168.755 106.295 168.925 ;
        RECT 103.110 168.155 103.570 168.445 ;
        RECT 104.265 168.415 105.765 168.585 ;
        RECT 104.265 168.275 104.435 168.415 ;
        RECT 103.875 168.105 104.435 168.275 ;
        RECT 102.350 167.475 102.600 167.935 ;
        RECT 102.770 167.645 103.640 167.985 ;
        RECT 103.875 167.645 104.045 168.105 ;
        RECT 104.880 168.075 105.955 168.245 ;
        RECT 104.215 167.475 104.585 167.935 ;
        RECT 104.880 167.735 105.050 168.075 ;
        RECT 105.220 167.475 105.550 167.905 ;
        RECT 105.785 167.735 105.955 168.075 ;
        RECT 106.125 167.975 106.295 168.755 ;
        RECT 106.465 168.535 106.635 169.125 ;
        RECT 106.805 168.725 107.155 169.345 ;
        RECT 106.465 168.145 106.930 168.535 ;
        RECT 107.325 168.275 107.495 169.635 ;
        RECT 107.665 168.445 108.125 169.495 ;
        RECT 107.100 168.105 107.495 168.275 ;
        RECT 107.100 167.975 107.270 168.105 ;
        RECT 106.125 167.645 106.805 167.975 ;
        RECT 107.020 167.645 107.270 167.975 ;
        RECT 107.440 167.475 107.690 167.935 ;
        RECT 107.860 167.660 108.185 168.445 ;
        RECT 108.355 167.645 108.525 169.765 ;
        RECT 108.695 169.645 109.025 170.025 ;
        RECT 109.195 169.475 109.450 169.765 ;
        RECT 109.625 169.480 114.970 170.025 ;
        RECT 108.700 169.305 109.450 169.475 ;
        RECT 108.700 168.315 108.930 169.305 ;
        RECT 109.100 168.485 109.450 169.135 ;
        RECT 111.210 168.650 111.550 169.480 ;
        RECT 115.145 169.255 118.655 170.025 ;
        RECT 119.285 169.300 119.575 170.025 ;
        RECT 120.665 169.275 121.875 170.025 ;
        RECT 108.700 168.145 109.450 168.315 ;
        RECT 108.695 167.475 109.025 167.975 ;
        RECT 109.195 167.645 109.450 168.145 ;
        RECT 113.030 167.910 113.380 169.160 ;
        RECT 115.145 168.735 116.795 169.255 ;
        RECT 116.965 168.565 118.655 169.085 ;
        RECT 109.625 167.475 114.970 167.910 ;
        RECT 115.145 167.475 118.655 168.565 ;
        RECT 119.285 167.475 119.575 168.640 ;
        RECT 120.665 168.565 121.185 169.105 ;
        RECT 121.355 168.735 121.875 169.275 ;
        RECT 120.665 167.475 121.875 168.565 ;
        RECT 67.680 167.305 121.960 167.475 ;
        RECT 67.765 166.215 68.975 167.305 ;
        RECT 69.145 166.870 74.490 167.305 ;
        RECT 74.665 166.870 80.010 167.305 ;
        RECT 67.765 165.505 68.285 166.045 ;
        RECT 68.455 165.675 68.975 166.215 ;
        RECT 67.765 164.755 68.975 165.505 ;
        RECT 70.730 165.300 71.070 166.130 ;
        RECT 72.550 165.620 72.900 166.870 ;
        RECT 76.250 165.300 76.590 166.130 ;
        RECT 78.070 165.620 78.420 166.870 ;
        RECT 80.645 166.140 80.935 167.305 ;
        RECT 81.105 166.215 84.615 167.305 ;
        RECT 81.105 165.525 82.755 166.045 ;
        RECT 82.925 165.695 84.615 166.215 ;
        RECT 85.255 166.695 85.585 167.125 ;
        RECT 85.765 166.865 85.960 167.305 ;
        RECT 86.130 166.695 86.460 167.125 ;
        RECT 85.255 166.525 86.460 166.695 ;
        RECT 85.255 166.195 86.150 166.525 ;
        RECT 86.630 166.355 86.905 167.125 ;
        RECT 86.320 166.165 86.905 166.355 ;
        RECT 87.095 166.335 87.425 167.120 ;
        RECT 87.095 166.165 87.775 166.335 ;
        RECT 87.955 166.165 88.285 167.305 ;
        RECT 88.555 166.635 88.725 167.135 ;
        RECT 88.895 166.805 89.225 167.305 ;
        RECT 88.555 166.465 89.220 166.635 ;
        RECT 85.260 165.665 85.555 165.995 ;
        RECT 85.735 165.665 86.150 165.995 ;
        RECT 69.145 164.755 74.490 165.300 ;
        RECT 74.665 164.755 80.010 165.300 ;
        RECT 80.645 164.755 80.935 165.480 ;
        RECT 81.105 164.755 84.615 165.525 ;
        RECT 85.255 164.755 85.555 165.485 ;
        RECT 85.735 165.045 85.965 165.665 ;
        RECT 86.320 165.495 86.495 166.165 ;
        RECT 86.165 165.315 86.495 165.495 ;
        RECT 86.665 165.345 86.905 165.995 ;
        RECT 87.085 165.745 87.435 165.995 ;
        RECT 87.605 165.565 87.775 166.165 ;
        RECT 87.945 165.745 88.295 165.995 ;
        RECT 88.470 165.645 88.820 166.295 ;
        RECT 86.165 164.935 86.390 165.315 ;
        RECT 86.560 164.755 86.890 165.145 ;
        RECT 87.105 164.755 87.345 165.565 ;
        RECT 87.515 164.925 87.845 165.565 ;
        RECT 88.015 164.755 88.285 165.565 ;
        RECT 88.990 165.475 89.220 166.465 ;
        RECT 88.555 165.305 89.220 165.475 ;
        RECT 88.555 165.015 88.725 165.305 ;
        RECT 88.895 164.755 89.225 165.135 ;
        RECT 89.395 165.015 89.620 167.135 ;
        RECT 89.820 166.845 90.085 167.305 ;
        RECT 90.270 166.735 90.505 167.110 ;
        RECT 90.750 166.860 91.820 167.030 ;
        RECT 89.820 165.735 90.100 166.335 ;
        RECT 89.835 164.755 90.085 165.215 ;
        RECT 90.270 165.205 90.440 166.735 ;
        RECT 90.610 165.705 90.850 166.575 ;
        RECT 91.040 166.325 91.480 166.680 ;
        RECT 91.650 166.245 91.820 166.860 ;
        RECT 91.990 166.505 92.160 167.305 ;
        RECT 92.330 166.805 92.580 167.135 ;
        RECT 92.805 166.835 93.690 167.005 ;
        RECT 91.650 166.155 92.160 166.245 ;
        RECT 91.360 165.985 92.160 166.155 ;
        RECT 90.610 165.375 91.190 165.705 ;
        RECT 91.360 165.205 91.530 165.985 ;
        RECT 91.990 165.915 92.160 165.985 ;
        RECT 91.700 165.735 91.870 165.765 ;
        RECT 92.330 165.735 92.500 166.805 ;
        RECT 92.670 165.915 92.860 166.635 ;
        RECT 93.030 166.245 93.350 166.575 ;
        RECT 91.700 165.435 92.500 165.735 ;
        RECT 93.030 165.705 93.220 166.245 ;
        RECT 90.270 165.035 90.600 165.205 ;
        RECT 90.780 165.035 91.530 165.205 ;
        RECT 91.780 164.755 92.150 165.255 ;
        RECT 92.330 165.205 92.500 165.435 ;
        RECT 92.670 165.375 93.220 165.705 ;
        RECT 93.520 165.915 93.690 166.835 ;
        RECT 93.870 166.805 94.085 167.305 ;
        RECT 94.550 166.500 94.720 167.125 ;
        RECT 95.005 166.525 95.185 167.305 ;
        RECT 93.860 166.340 94.720 166.500 ;
        RECT 93.860 166.170 94.970 166.340 ;
        RECT 94.800 165.915 94.970 166.170 ;
        RECT 95.365 166.305 95.700 167.065 ;
        RECT 95.880 166.475 96.050 167.305 ;
        RECT 96.220 166.305 96.550 167.065 ;
        RECT 96.720 166.475 96.890 167.305 ;
        RECT 95.365 166.135 97.035 166.305 ;
        RECT 97.205 166.215 100.715 167.305 ;
        RECT 93.520 165.745 94.610 165.915 ;
        RECT 94.800 165.745 96.620 165.915 ;
        RECT 93.520 165.205 93.690 165.745 ;
        RECT 94.800 165.575 94.970 165.745 ;
        RECT 94.470 165.405 94.970 165.575 ;
        RECT 96.790 165.570 97.035 166.135 ;
        RECT 92.330 165.035 92.790 165.205 ;
        RECT 93.020 165.035 93.690 165.205 ;
        RECT 94.005 164.755 94.175 165.285 ;
        RECT 94.470 164.965 94.830 165.405 ;
        RECT 95.365 165.400 97.035 165.570 ;
        RECT 97.205 165.525 98.855 166.045 ;
        RECT 99.025 165.695 100.715 166.215 ;
        RECT 101.345 166.230 101.615 167.135 ;
        RECT 101.785 166.545 102.115 167.305 ;
        RECT 102.295 166.375 102.475 167.135 ;
        RECT 95.005 164.755 95.175 165.235 ;
        RECT 95.365 164.975 95.700 165.400 ;
        RECT 95.875 164.755 96.045 165.230 ;
        RECT 96.220 164.975 96.555 165.400 ;
        RECT 96.725 164.755 96.895 165.230 ;
        RECT 97.205 164.755 100.715 165.525 ;
        RECT 101.345 165.430 101.525 166.230 ;
        RECT 101.800 166.205 102.475 166.375 ;
        RECT 102.725 166.215 106.235 167.305 ;
        RECT 101.800 166.060 101.970 166.205 ;
        RECT 101.695 165.730 101.970 166.060 ;
        RECT 101.800 165.475 101.970 165.730 ;
        RECT 102.195 165.655 102.535 166.025 ;
        RECT 102.725 165.525 104.375 166.045 ;
        RECT 104.545 165.695 106.235 166.215 ;
        RECT 106.405 166.140 106.695 167.305 ;
        RECT 106.865 166.870 112.210 167.305 ;
        RECT 112.385 166.870 117.730 167.305 ;
        RECT 101.345 164.925 101.605 165.430 ;
        RECT 101.800 165.305 102.465 165.475 ;
        RECT 101.785 164.755 102.115 165.135 ;
        RECT 102.295 164.925 102.465 165.305 ;
        RECT 102.725 164.755 106.235 165.525 ;
        RECT 106.405 164.755 106.695 165.480 ;
        RECT 108.450 165.300 108.790 166.130 ;
        RECT 110.270 165.620 110.620 166.870 ;
        RECT 113.970 165.300 114.310 166.130 ;
        RECT 115.790 165.620 116.140 166.870 ;
        RECT 117.905 166.215 120.495 167.305 ;
        RECT 117.905 165.525 119.115 166.045 ;
        RECT 119.285 165.695 120.495 166.215 ;
        RECT 120.665 166.215 121.875 167.305 ;
        RECT 120.665 165.675 121.185 166.215 ;
        RECT 106.865 164.755 112.210 165.300 ;
        RECT 112.385 164.755 117.730 165.300 ;
        RECT 117.905 164.755 120.495 165.525 ;
        RECT 121.355 165.505 121.875 166.045 ;
        RECT 120.665 164.755 121.875 165.505 ;
        RECT 67.680 164.585 121.960 164.755 ;
        RECT 67.765 163.835 68.975 164.585 ;
        RECT 69.145 164.040 74.490 164.585 ;
        RECT 74.665 164.040 80.010 164.585 ;
        RECT 80.185 164.040 85.530 164.585 ;
        RECT 67.765 163.295 68.285 163.835 ;
        RECT 68.455 163.125 68.975 163.665 ;
        RECT 70.730 163.210 71.070 164.040 ;
        RECT 67.765 162.035 68.975 163.125 ;
        RECT 72.550 162.470 72.900 163.720 ;
        RECT 76.250 163.210 76.590 164.040 ;
        RECT 78.070 162.470 78.420 163.720 ;
        RECT 81.770 163.210 82.110 164.040 ;
        RECT 85.705 163.815 89.215 164.585 ;
        RECT 89.385 163.835 90.595 164.585 ;
        RECT 83.590 162.470 83.940 163.720 ;
        RECT 85.705 163.295 87.355 163.815 ;
        RECT 87.525 163.125 89.215 163.645 ;
        RECT 89.385 163.295 89.905 163.835 ;
        RECT 90.075 163.125 90.595 163.665 ;
        RECT 69.145 162.035 74.490 162.470 ;
        RECT 74.665 162.035 80.010 162.470 ;
        RECT 80.185 162.035 85.530 162.470 ;
        RECT 85.705 162.035 89.215 163.125 ;
        RECT 89.385 162.035 90.595 163.125 ;
        RECT 90.765 163.640 91.105 164.415 ;
        RECT 91.275 164.125 91.445 164.585 ;
        RECT 91.685 164.150 92.045 164.415 ;
        RECT 91.685 164.145 92.040 164.150 ;
        RECT 91.685 164.135 92.035 164.145 ;
        RECT 91.685 164.130 92.030 164.135 ;
        RECT 91.685 164.120 92.025 164.130 ;
        RECT 92.675 164.125 92.845 164.585 ;
        RECT 91.685 164.115 92.020 164.120 ;
        RECT 91.685 164.105 92.010 164.115 ;
        RECT 91.685 164.095 92.000 164.105 ;
        RECT 91.685 163.955 91.985 164.095 ;
        RECT 91.275 163.765 91.985 163.955 ;
        RECT 92.175 163.955 92.505 164.035 ;
        RECT 93.015 163.955 93.355 164.415 ;
        RECT 92.175 163.765 93.355 163.955 ;
        RECT 93.525 163.860 93.815 164.585 ;
        RECT 94.010 164.195 94.340 164.585 ;
        RECT 94.510 164.025 94.735 164.405 ;
        RECT 90.765 162.205 91.045 163.640 ;
        RECT 91.275 163.195 91.560 163.765 ;
        RECT 91.745 163.365 92.215 163.595 ;
        RECT 92.385 163.575 92.715 163.595 ;
        RECT 92.385 163.395 92.835 163.575 ;
        RECT 93.025 163.395 93.355 163.595 ;
        RECT 91.275 162.980 92.425 163.195 ;
        RECT 91.215 162.035 91.925 162.810 ;
        RECT 92.095 162.205 92.425 162.980 ;
        RECT 92.620 162.280 92.835 163.395 ;
        RECT 93.125 163.055 93.355 163.395 ;
        RECT 93.995 163.345 94.235 163.995 ;
        RECT 94.405 163.845 94.735 164.025 ;
        RECT 93.015 162.035 93.345 162.755 ;
        RECT 93.525 162.035 93.815 163.200 ;
        RECT 94.405 163.175 94.580 163.845 ;
        RECT 94.935 163.675 95.165 164.295 ;
        RECT 95.345 163.855 95.645 164.585 ;
        RECT 96.425 164.110 96.595 164.585 ;
        RECT 96.765 163.940 97.100 164.365 ;
        RECT 97.275 164.110 97.445 164.585 ;
        RECT 97.620 163.940 97.955 164.365 ;
        RECT 98.145 164.105 98.315 164.585 ;
        RECT 96.285 163.770 97.955 163.940 ;
        RECT 98.490 163.935 98.850 164.375 ;
        RECT 99.145 164.055 99.315 164.585 ;
        RECT 99.630 164.135 100.300 164.305 ;
        RECT 100.530 164.135 100.990 164.305 ;
        RECT 94.750 163.345 95.165 163.675 ;
        RECT 95.345 163.345 95.640 163.675 ;
        RECT 93.995 162.985 94.580 163.175 ;
        RECT 96.285 163.205 96.530 163.770 ;
        RECT 98.350 163.765 98.850 163.935 ;
        RECT 98.350 163.595 98.520 163.765 ;
        RECT 99.630 163.595 99.800 164.135 ;
        RECT 96.700 163.425 98.520 163.595 ;
        RECT 98.710 163.425 99.800 163.595 ;
        RECT 93.995 162.215 94.270 162.985 ;
        RECT 94.750 162.815 95.645 163.145 ;
        RECT 96.285 163.035 97.955 163.205 ;
        RECT 94.440 162.645 95.645 162.815 ;
        RECT 94.440 162.215 94.770 162.645 ;
        RECT 94.940 162.035 95.135 162.475 ;
        RECT 95.315 162.215 95.645 162.645 ;
        RECT 96.430 162.035 96.600 162.865 ;
        RECT 96.770 162.275 97.100 163.035 ;
        RECT 97.270 162.035 97.440 162.865 ;
        RECT 97.620 162.275 97.955 163.035 ;
        RECT 98.350 163.170 98.520 163.425 ;
        RECT 98.350 163.000 99.460 163.170 ;
        RECT 98.600 162.840 99.460 163.000 ;
        RECT 98.135 162.035 98.315 162.815 ;
        RECT 98.600 162.215 98.770 162.840 ;
        RECT 99.235 162.035 99.450 162.535 ;
        RECT 99.630 162.505 99.800 163.425 ;
        RECT 100.100 163.635 100.650 163.965 ;
        RECT 100.820 163.905 100.990 164.135 ;
        RECT 101.170 164.085 101.540 164.585 ;
        RECT 101.790 164.135 102.540 164.305 ;
        RECT 102.720 164.135 103.050 164.305 ;
        RECT 100.100 163.095 100.290 163.635 ;
        RECT 100.820 163.605 101.620 163.905 ;
        RECT 99.970 162.765 100.290 163.095 ;
        RECT 100.460 162.705 100.650 163.425 ;
        RECT 100.820 162.535 100.990 163.605 ;
        RECT 101.450 163.575 101.620 163.605 ;
        RECT 101.160 163.355 101.330 163.425 ;
        RECT 101.790 163.355 101.960 164.135 ;
        RECT 102.130 163.635 102.710 163.965 ;
        RECT 101.160 163.185 101.960 163.355 ;
        RECT 101.160 163.095 101.670 163.185 ;
        RECT 99.630 162.335 100.515 162.505 ;
        RECT 100.740 162.205 100.990 162.535 ;
        RECT 101.160 162.035 101.330 162.835 ;
        RECT 101.500 162.480 101.670 163.095 ;
        RECT 101.840 162.660 102.280 163.015 ;
        RECT 102.470 162.765 102.710 163.635 ;
        RECT 102.880 162.605 103.050 164.135 ;
        RECT 103.235 164.125 103.485 164.585 ;
        RECT 103.220 163.005 103.500 163.605 ;
        RECT 101.500 162.310 102.570 162.480 ;
        RECT 102.815 162.230 103.050 162.605 ;
        RECT 103.235 162.035 103.500 162.495 ;
        RECT 103.700 162.205 103.925 164.325 ;
        RECT 104.095 164.205 104.425 164.585 ;
        RECT 104.595 164.035 104.765 164.325 ;
        RECT 105.025 164.040 110.370 164.585 ;
        RECT 110.545 164.040 115.890 164.585 ;
        RECT 104.100 163.865 104.765 164.035 ;
        RECT 104.100 162.875 104.330 163.865 ;
        RECT 104.500 163.045 104.850 163.695 ;
        RECT 106.610 163.210 106.950 164.040 ;
        RECT 104.100 162.705 104.765 162.875 ;
        RECT 104.095 162.035 104.425 162.535 ;
        RECT 104.595 162.205 104.765 162.705 ;
        RECT 108.430 162.470 108.780 163.720 ;
        RECT 112.130 163.210 112.470 164.040 ;
        RECT 116.065 163.815 118.655 164.585 ;
        RECT 119.285 163.860 119.575 164.585 ;
        RECT 120.665 163.835 121.875 164.585 ;
        RECT 113.950 162.470 114.300 163.720 ;
        RECT 116.065 163.295 117.275 163.815 ;
        RECT 117.445 163.125 118.655 163.645 ;
        RECT 105.025 162.035 110.370 162.470 ;
        RECT 110.545 162.035 115.890 162.470 ;
        RECT 116.065 162.035 118.655 163.125 ;
        RECT 119.285 162.035 119.575 163.200 ;
        RECT 120.665 163.125 121.185 163.665 ;
        RECT 121.355 163.295 121.875 163.835 ;
        RECT 120.665 162.035 121.875 163.125 ;
        RECT 67.680 161.865 121.960 162.035 ;
        RECT 67.765 160.775 68.975 161.865 ;
        RECT 69.145 161.430 74.490 161.865 ;
        RECT 74.665 161.430 80.010 161.865 ;
        RECT 67.765 160.065 68.285 160.605 ;
        RECT 68.455 160.235 68.975 160.775 ;
        RECT 67.765 159.315 68.975 160.065 ;
        RECT 70.730 159.860 71.070 160.690 ;
        RECT 72.550 160.180 72.900 161.430 ;
        RECT 76.250 159.860 76.590 160.690 ;
        RECT 78.070 160.180 78.420 161.430 ;
        RECT 80.645 160.700 80.935 161.865 ;
        RECT 81.195 161.120 81.465 161.865 ;
        RECT 82.095 161.860 88.370 161.865 ;
        RECT 81.635 160.950 81.925 161.690 ;
        RECT 82.095 161.135 82.350 161.860 ;
        RECT 82.535 160.965 82.795 161.690 ;
        RECT 82.965 161.135 83.210 161.860 ;
        RECT 83.395 160.965 83.655 161.690 ;
        RECT 83.825 161.135 84.070 161.860 ;
        RECT 84.255 160.965 84.515 161.690 ;
        RECT 84.685 161.135 84.930 161.860 ;
        RECT 85.100 160.965 85.360 161.690 ;
        RECT 85.530 161.135 85.790 161.860 ;
        RECT 85.960 160.965 86.220 161.690 ;
        RECT 86.390 161.135 86.650 161.860 ;
        RECT 86.820 160.965 87.080 161.690 ;
        RECT 87.250 161.135 87.510 161.860 ;
        RECT 87.680 160.965 87.940 161.690 ;
        RECT 88.110 161.065 88.370 161.860 ;
        RECT 82.535 160.950 87.940 160.965 ;
        RECT 81.195 160.725 87.940 160.950 ;
        RECT 81.195 160.135 82.360 160.725 ;
        RECT 88.540 160.555 88.790 161.690 ;
        RECT 88.970 161.055 89.230 161.865 ;
        RECT 89.405 160.555 89.650 161.695 ;
        RECT 89.830 161.055 90.125 161.865 ;
        RECT 90.305 160.775 92.895 161.865 ;
        RECT 82.530 160.305 89.650 160.555 ;
        RECT 69.145 159.315 74.490 159.860 ;
        RECT 74.665 159.315 80.010 159.860 ;
        RECT 80.645 159.315 80.935 160.040 ;
        RECT 81.195 159.965 87.940 160.135 ;
        RECT 81.195 159.315 81.495 159.795 ;
        RECT 81.665 159.510 81.925 159.965 ;
        RECT 82.095 159.315 82.355 159.795 ;
        RECT 82.535 159.510 82.795 159.965 ;
        RECT 82.965 159.315 83.215 159.795 ;
        RECT 83.395 159.510 83.655 159.965 ;
        RECT 83.825 159.315 84.075 159.795 ;
        RECT 84.255 159.510 84.515 159.965 ;
        RECT 84.685 159.315 84.930 159.795 ;
        RECT 85.100 159.510 85.375 159.965 ;
        RECT 85.545 159.315 85.790 159.795 ;
        RECT 85.960 159.510 86.220 159.965 ;
        RECT 86.390 159.315 86.650 159.795 ;
        RECT 86.820 159.510 87.080 159.965 ;
        RECT 87.250 159.315 87.510 159.795 ;
        RECT 87.680 159.510 87.940 159.965 ;
        RECT 88.110 159.315 88.370 159.875 ;
        RECT 88.540 159.495 88.790 160.305 ;
        RECT 88.970 159.315 89.230 159.840 ;
        RECT 89.400 159.495 89.650 160.305 ;
        RECT 89.820 159.995 90.135 160.555 ;
        RECT 90.305 160.085 91.515 160.605 ;
        RECT 91.685 160.255 92.895 160.775 ;
        RECT 93.525 160.700 93.815 161.865 ;
        RECT 93.985 160.775 97.495 161.865 ;
        RECT 97.780 161.235 98.065 161.695 ;
        RECT 98.235 161.405 98.505 161.865 ;
        RECT 97.780 161.015 98.735 161.235 ;
        RECT 93.985 160.085 95.635 160.605 ;
        RECT 95.805 160.255 97.495 160.775 ;
        RECT 97.665 160.285 98.355 160.845 ;
        RECT 98.525 160.115 98.735 161.015 ;
        RECT 89.830 159.315 90.135 159.825 ;
        RECT 90.305 159.315 92.895 160.085 ;
        RECT 93.525 159.315 93.815 160.040 ;
        RECT 93.985 159.315 97.495 160.085 ;
        RECT 97.780 159.945 98.735 160.115 ;
        RECT 98.905 160.845 99.305 161.695 ;
        RECT 99.495 161.235 99.775 161.695 ;
        RECT 100.295 161.405 100.620 161.865 ;
        RECT 99.495 161.015 100.620 161.235 ;
        RECT 98.905 160.285 100.000 160.845 ;
        RECT 100.170 160.555 100.620 161.015 ;
        RECT 100.790 160.725 101.175 161.695 ;
        RECT 101.355 160.895 101.685 161.680 ;
        RECT 101.355 160.725 102.035 160.895 ;
        RECT 102.215 160.725 102.545 161.865 ;
        RECT 102.725 160.775 106.235 161.865 ;
        RECT 97.780 159.485 98.065 159.945 ;
        RECT 98.235 159.315 98.505 159.775 ;
        RECT 98.905 159.485 99.305 160.285 ;
        RECT 100.170 160.225 100.725 160.555 ;
        RECT 100.170 160.115 100.620 160.225 ;
        RECT 99.495 159.945 100.620 160.115 ;
        RECT 100.895 160.055 101.175 160.725 ;
        RECT 101.345 160.305 101.695 160.555 ;
        RECT 101.865 160.125 102.035 160.725 ;
        RECT 102.205 160.305 102.555 160.555 ;
        RECT 99.495 159.485 99.775 159.945 ;
        RECT 100.295 159.315 100.620 159.775 ;
        RECT 100.790 159.485 101.175 160.055 ;
        RECT 101.365 159.315 101.605 160.125 ;
        RECT 101.775 159.485 102.105 160.125 ;
        RECT 102.275 159.315 102.545 160.125 ;
        RECT 102.725 160.085 104.375 160.605 ;
        RECT 104.545 160.255 106.235 160.775 ;
        RECT 106.405 160.700 106.695 161.865 ;
        RECT 106.875 161.055 107.170 161.865 ;
        RECT 107.350 160.555 107.595 161.695 ;
        RECT 107.770 161.055 108.030 161.865 ;
        RECT 108.630 161.860 114.905 161.865 ;
        RECT 108.210 160.555 108.460 161.690 ;
        RECT 108.630 161.065 108.890 161.860 ;
        RECT 109.060 160.965 109.320 161.690 ;
        RECT 109.490 161.135 109.750 161.860 ;
        RECT 109.920 160.965 110.180 161.690 ;
        RECT 110.350 161.135 110.610 161.860 ;
        RECT 110.780 160.965 111.040 161.690 ;
        RECT 111.210 161.135 111.470 161.860 ;
        RECT 111.640 160.965 111.900 161.690 ;
        RECT 112.070 161.135 112.315 161.860 ;
        RECT 112.485 160.965 112.745 161.690 ;
        RECT 112.930 161.135 113.175 161.860 ;
        RECT 113.345 160.965 113.605 161.690 ;
        RECT 113.790 161.135 114.035 161.860 ;
        RECT 114.205 160.965 114.465 161.690 ;
        RECT 114.650 161.135 114.905 161.860 ;
        RECT 109.060 160.950 114.465 160.965 ;
        RECT 115.075 160.950 115.365 161.690 ;
        RECT 115.535 161.120 115.805 161.865 ;
        RECT 109.060 160.725 115.805 160.950 ;
        RECT 116.065 160.775 118.655 161.865 ;
        RECT 102.725 159.315 106.235 160.085 ;
        RECT 106.405 159.315 106.695 160.040 ;
        RECT 106.865 159.995 107.180 160.555 ;
        RECT 107.350 160.305 114.470 160.555 ;
        RECT 106.865 159.315 107.170 159.825 ;
        RECT 107.350 159.495 107.600 160.305 ;
        RECT 107.770 159.315 108.030 159.840 ;
        RECT 108.210 159.495 108.460 160.305 ;
        RECT 114.640 160.135 115.805 160.725 ;
        RECT 109.060 159.965 115.805 160.135 ;
        RECT 116.065 160.085 117.275 160.605 ;
        RECT 117.445 160.255 118.655 160.775 ;
        RECT 119.285 160.700 119.575 161.865 ;
        RECT 120.665 160.775 121.875 161.865 ;
        RECT 120.665 160.235 121.185 160.775 ;
        RECT 108.630 159.315 108.890 159.875 ;
        RECT 109.060 159.510 109.320 159.965 ;
        RECT 109.490 159.315 109.750 159.795 ;
        RECT 109.920 159.510 110.180 159.965 ;
        RECT 110.350 159.315 110.610 159.795 ;
        RECT 110.780 159.510 111.040 159.965 ;
        RECT 111.210 159.315 111.455 159.795 ;
        RECT 111.625 159.510 111.900 159.965 ;
        RECT 112.070 159.315 112.315 159.795 ;
        RECT 112.485 159.510 112.745 159.965 ;
        RECT 112.925 159.315 113.175 159.795 ;
        RECT 113.345 159.510 113.605 159.965 ;
        RECT 113.785 159.315 114.035 159.795 ;
        RECT 114.205 159.510 114.465 159.965 ;
        RECT 114.645 159.315 114.905 159.795 ;
        RECT 115.075 159.510 115.335 159.965 ;
        RECT 115.505 159.315 115.805 159.795 ;
        RECT 116.065 159.315 118.655 160.085 ;
        RECT 121.355 160.065 121.875 160.605 ;
        RECT 119.285 159.315 119.575 160.040 ;
        RECT 120.665 159.315 121.875 160.065 ;
        RECT 67.680 159.145 121.960 159.315 ;
        RECT 86.550 91.940 86.880 92.110 ;
        RECT 86.630 90.125 86.800 91.940 ;
        RECT 88.640 91.900 88.970 92.070 ;
        RECT 95.400 92.000 95.730 92.170 ;
        RECT 88.720 90.085 88.890 91.900 ;
        RECT 90.760 91.750 91.090 91.920 ;
        RECT 93.030 91.750 93.360 91.920 ;
        RECT 90.840 89.935 91.010 91.750 ;
        RECT 93.110 89.935 93.280 91.750 ;
        RECT 95.480 90.185 95.650 92.000 ;
        RECT 86.630 74.450 86.800 76.265 ;
        RECT 86.550 74.280 86.880 74.450 ;
        RECT 88.720 74.410 88.890 76.225 ;
        RECT 88.640 74.240 88.970 74.410 ;
        RECT 90.840 74.260 91.010 76.075 ;
        RECT 93.110 74.260 93.280 76.075 ;
        RECT 95.480 74.510 95.650 76.325 ;
        RECT 95.400 74.340 95.730 74.510 ;
        RECT 90.760 74.090 91.090 74.260 ;
        RECT 93.030 74.090 93.360 74.260 ;
        RECT 90.760 71.230 91.090 71.400 ;
        RECT 93.130 71.380 93.460 71.550 ;
        RECT 90.840 69.415 91.010 71.230 ;
        RECT 93.210 69.565 93.380 71.380 ;
        RECT 95.500 71.130 95.830 71.300 ;
        RECT 95.580 69.315 95.750 71.130 ;
        RECT 90.840 60.580 91.010 62.395 ;
        RECT 93.210 60.730 93.380 62.545 ;
        RECT 90.760 60.410 91.090 60.580 ;
        RECT 93.130 60.560 93.460 60.730 ;
        RECT 95.580 60.480 95.750 62.295 ;
        RECT 95.500 60.310 95.830 60.480 ;
      LAYER mcon ;
        RECT 67.825 213.545 67.995 213.715 ;
        RECT 68.285 213.545 68.455 213.715 ;
        RECT 68.745 213.545 68.915 213.715 ;
        RECT 69.205 213.545 69.375 213.715 ;
        RECT 69.665 213.545 69.835 213.715 ;
        RECT 70.125 213.545 70.295 213.715 ;
        RECT 70.585 213.545 70.755 213.715 ;
        RECT 71.045 213.545 71.215 213.715 ;
        RECT 71.505 213.545 71.675 213.715 ;
        RECT 71.965 213.545 72.135 213.715 ;
        RECT 72.425 213.545 72.595 213.715 ;
        RECT 72.885 213.545 73.055 213.715 ;
        RECT 73.345 213.545 73.515 213.715 ;
        RECT 73.805 213.545 73.975 213.715 ;
        RECT 74.265 213.545 74.435 213.715 ;
        RECT 74.725 213.545 74.895 213.715 ;
        RECT 75.185 213.545 75.355 213.715 ;
        RECT 75.645 213.545 75.815 213.715 ;
        RECT 76.105 213.545 76.275 213.715 ;
        RECT 76.565 213.545 76.735 213.715 ;
        RECT 77.025 213.545 77.195 213.715 ;
        RECT 77.485 213.545 77.655 213.715 ;
        RECT 77.945 213.545 78.115 213.715 ;
        RECT 78.405 213.545 78.575 213.715 ;
        RECT 78.865 213.545 79.035 213.715 ;
        RECT 79.325 213.545 79.495 213.715 ;
        RECT 79.785 213.545 79.955 213.715 ;
        RECT 80.245 213.545 80.415 213.715 ;
        RECT 80.705 213.545 80.875 213.715 ;
        RECT 81.165 213.545 81.335 213.715 ;
        RECT 81.625 213.545 81.795 213.715 ;
        RECT 82.085 213.545 82.255 213.715 ;
        RECT 82.545 213.545 82.715 213.715 ;
        RECT 83.005 213.545 83.175 213.715 ;
        RECT 83.465 213.545 83.635 213.715 ;
        RECT 83.925 213.545 84.095 213.715 ;
        RECT 84.385 213.545 84.555 213.715 ;
        RECT 84.845 213.545 85.015 213.715 ;
        RECT 85.305 213.545 85.475 213.715 ;
        RECT 85.765 213.545 85.935 213.715 ;
        RECT 86.225 213.545 86.395 213.715 ;
        RECT 86.685 213.545 86.855 213.715 ;
        RECT 87.145 213.545 87.315 213.715 ;
        RECT 87.605 213.545 87.775 213.715 ;
        RECT 88.065 213.545 88.235 213.715 ;
        RECT 88.525 213.545 88.695 213.715 ;
        RECT 88.985 213.545 89.155 213.715 ;
        RECT 89.445 213.545 89.615 213.715 ;
        RECT 89.905 213.545 90.075 213.715 ;
        RECT 90.365 213.545 90.535 213.715 ;
        RECT 90.825 213.545 90.995 213.715 ;
        RECT 91.285 213.545 91.455 213.715 ;
        RECT 91.745 213.545 91.915 213.715 ;
        RECT 92.205 213.545 92.375 213.715 ;
        RECT 92.665 213.545 92.835 213.715 ;
        RECT 93.125 213.545 93.295 213.715 ;
        RECT 93.585 213.545 93.755 213.715 ;
        RECT 94.045 213.545 94.215 213.715 ;
        RECT 94.505 213.545 94.675 213.715 ;
        RECT 94.965 213.545 95.135 213.715 ;
        RECT 95.425 213.545 95.595 213.715 ;
        RECT 95.885 213.545 96.055 213.715 ;
        RECT 96.345 213.545 96.515 213.715 ;
        RECT 96.805 213.545 96.975 213.715 ;
        RECT 97.265 213.545 97.435 213.715 ;
        RECT 97.725 213.545 97.895 213.715 ;
        RECT 98.185 213.545 98.355 213.715 ;
        RECT 98.645 213.545 98.815 213.715 ;
        RECT 99.105 213.545 99.275 213.715 ;
        RECT 99.565 213.545 99.735 213.715 ;
        RECT 100.025 213.545 100.195 213.715 ;
        RECT 100.485 213.545 100.655 213.715 ;
        RECT 100.945 213.545 101.115 213.715 ;
        RECT 101.405 213.545 101.575 213.715 ;
        RECT 101.865 213.545 102.035 213.715 ;
        RECT 102.325 213.545 102.495 213.715 ;
        RECT 102.785 213.545 102.955 213.715 ;
        RECT 103.245 213.545 103.415 213.715 ;
        RECT 103.705 213.545 103.875 213.715 ;
        RECT 104.165 213.545 104.335 213.715 ;
        RECT 104.625 213.545 104.795 213.715 ;
        RECT 105.085 213.545 105.255 213.715 ;
        RECT 105.545 213.545 105.715 213.715 ;
        RECT 106.005 213.545 106.175 213.715 ;
        RECT 106.465 213.545 106.635 213.715 ;
        RECT 106.925 213.545 107.095 213.715 ;
        RECT 107.385 213.545 107.555 213.715 ;
        RECT 107.845 213.545 108.015 213.715 ;
        RECT 108.305 213.545 108.475 213.715 ;
        RECT 108.765 213.545 108.935 213.715 ;
        RECT 109.225 213.545 109.395 213.715 ;
        RECT 109.685 213.545 109.855 213.715 ;
        RECT 110.145 213.545 110.315 213.715 ;
        RECT 110.605 213.545 110.775 213.715 ;
        RECT 111.065 213.545 111.235 213.715 ;
        RECT 111.525 213.545 111.695 213.715 ;
        RECT 111.985 213.545 112.155 213.715 ;
        RECT 112.445 213.545 112.615 213.715 ;
        RECT 112.905 213.545 113.075 213.715 ;
        RECT 113.365 213.545 113.535 213.715 ;
        RECT 113.825 213.545 113.995 213.715 ;
        RECT 114.285 213.545 114.455 213.715 ;
        RECT 114.745 213.545 114.915 213.715 ;
        RECT 115.205 213.545 115.375 213.715 ;
        RECT 115.665 213.545 115.835 213.715 ;
        RECT 116.125 213.545 116.295 213.715 ;
        RECT 116.585 213.545 116.755 213.715 ;
        RECT 117.045 213.545 117.215 213.715 ;
        RECT 117.505 213.545 117.675 213.715 ;
        RECT 117.965 213.545 118.135 213.715 ;
        RECT 118.425 213.545 118.595 213.715 ;
        RECT 118.885 213.545 119.055 213.715 ;
        RECT 119.345 213.545 119.515 213.715 ;
        RECT 119.805 213.545 119.975 213.715 ;
        RECT 120.265 213.545 120.435 213.715 ;
        RECT 120.725 213.545 120.895 213.715 ;
        RECT 121.185 213.545 121.355 213.715 ;
        RECT 121.645 213.545 121.815 213.715 ;
        RECT 67.825 210.825 67.995 210.995 ;
        RECT 68.285 210.825 68.455 210.995 ;
        RECT 68.745 210.825 68.915 210.995 ;
        RECT 69.205 210.825 69.375 210.995 ;
        RECT 69.665 210.825 69.835 210.995 ;
        RECT 70.125 210.825 70.295 210.995 ;
        RECT 70.585 210.825 70.755 210.995 ;
        RECT 71.045 210.825 71.215 210.995 ;
        RECT 71.505 210.825 71.675 210.995 ;
        RECT 71.965 210.825 72.135 210.995 ;
        RECT 72.425 210.825 72.595 210.995 ;
        RECT 72.885 210.825 73.055 210.995 ;
        RECT 73.345 210.825 73.515 210.995 ;
        RECT 73.805 210.825 73.975 210.995 ;
        RECT 74.265 210.825 74.435 210.995 ;
        RECT 74.725 210.825 74.895 210.995 ;
        RECT 75.185 210.825 75.355 210.995 ;
        RECT 75.645 210.825 75.815 210.995 ;
        RECT 76.105 210.825 76.275 210.995 ;
        RECT 76.565 210.825 76.735 210.995 ;
        RECT 77.025 210.825 77.195 210.995 ;
        RECT 77.485 210.825 77.655 210.995 ;
        RECT 77.945 210.825 78.115 210.995 ;
        RECT 78.405 210.825 78.575 210.995 ;
        RECT 78.865 210.825 79.035 210.995 ;
        RECT 79.325 210.825 79.495 210.995 ;
        RECT 79.785 210.825 79.955 210.995 ;
        RECT 80.245 210.825 80.415 210.995 ;
        RECT 80.705 210.825 80.875 210.995 ;
        RECT 81.165 210.825 81.335 210.995 ;
        RECT 81.625 210.825 81.795 210.995 ;
        RECT 82.085 210.825 82.255 210.995 ;
        RECT 82.545 210.825 82.715 210.995 ;
        RECT 83.005 210.825 83.175 210.995 ;
        RECT 83.465 210.825 83.635 210.995 ;
        RECT 83.925 210.825 84.095 210.995 ;
        RECT 84.385 210.825 84.555 210.995 ;
        RECT 84.845 210.825 85.015 210.995 ;
        RECT 85.305 210.825 85.475 210.995 ;
        RECT 85.765 210.825 85.935 210.995 ;
        RECT 86.225 210.825 86.395 210.995 ;
        RECT 86.685 210.825 86.855 210.995 ;
        RECT 87.145 210.825 87.315 210.995 ;
        RECT 87.605 210.825 87.775 210.995 ;
        RECT 88.065 210.825 88.235 210.995 ;
        RECT 88.525 210.825 88.695 210.995 ;
        RECT 88.985 210.825 89.155 210.995 ;
        RECT 89.445 210.825 89.615 210.995 ;
        RECT 89.905 210.825 90.075 210.995 ;
        RECT 90.365 210.825 90.535 210.995 ;
        RECT 90.825 210.825 90.995 210.995 ;
        RECT 91.285 210.825 91.455 210.995 ;
        RECT 91.745 210.825 91.915 210.995 ;
        RECT 92.205 210.825 92.375 210.995 ;
        RECT 92.665 210.825 92.835 210.995 ;
        RECT 93.125 210.825 93.295 210.995 ;
        RECT 93.585 210.825 93.755 210.995 ;
        RECT 94.045 210.825 94.215 210.995 ;
        RECT 94.505 210.825 94.675 210.995 ;
        RECT 94.965 210.825 95.135 210.995 ;
        RECT 95.425 210.825 95.595 210.995 ;
        RECT 95.885 210.825 96.055 210.995 ;
        RECT 96.345 210.825 96.515 210.995 ;
        RECT 96.805 210.825 96.975 210.995 ;
        RECT 97.265 210.825 97.435 210.995 ;
        RECT 97.725 210.825 97.895 210.995 ;
        RECT 98.185 210.825 98.355 210.995 ;
        RECT 98.645 210.825 98.815 210.995 ;
        RECT 99.105 210.825 99.275 210.995 ;
        RECT 99.565 210.825 99.735 210.995 ;
        RECT 100.025 210.825 100.195 210.995 ;
        RECT 100.485 210.825 100.655 210.995 ;
        RECT 100.945 210.825 101.115 210.995 ;
        RECT 101.405 210.825 101.575 210.995 ;
        RECT 101.865 210.825 102.035 210.995 ;
        RECT 102.325 210.825 102.495 210.995 ;
        RECT 102.785 210.825 102.955 210.995 ;
        RECT 103.245 210.825 103.415 210.995 ;
        RECT 103.705 210.825 103.875 210.995 ;
        RECT 104.165 210.825 104.335 210.995 ;
        RECT 104.625 210.825 104.795 210.995 ;
        RECT 105.085 210.825 105.255 210.995 ;
        RECT 105.545 210.825 105.715 210.995 ;
        RECT 106.005 210.825 106.175 210.995 ;
        RECT 106.465 210.825 106.635 210.995 ;
        RECT 106.925 210.825 107.095 210.995 ;
        RECT 107.385 210.825 107.555 210.995 ;
        RECT 107.845 210.825 108.015 210.995 ;
        RECT 108.305 210.825 108.475 210.995 ;
        RECT 108.765 210.825 108.935 210.995 ;
        RECT 109.225 210.825 109.395 210.995 ;
        RECT 109.685 210.825 109.855 210.995 ;
        RECT 110.145 210.825 110.315 210.995 ;
        RECT 110.605 210.825 110.775 210.995 ;
        RECT 111.065 210.825 111.235 210.995 ;
        RECT 111.525 210.825 111.695 210.995 ;
        RECT 111.985 210.825 112.155 210.995 ;
        RECT 112.445 210.825 112.615 210.995 ;
        RECT 112.905 210.825 113.075 210.995 ;
        RECT 113.365 210.825 113.535 210.995 ;
        RECT 113.825 210.825 113.995 210.995 ;
        RECT 114.285 210.825 114.455 210.995 ;
        RECT 114.745 210.825 114.915 210.995 ;
        RECT 115.205 210.825 115.375 210.995 ;
        RECT 115.665 210.825 115.835 210.995 ;
        RECT 116.125 210.825 116.295 210.995 ;
        RECT 116.585 210.825 116.755 210.995 ;
        RECT 117.045 210.825 117.215 210.995 ;
        RECT 117.505 210.825 117.675 210.995 ;
        RECT 117.965 210.825 118.135 210.995 ;
        RECT 118.425 210.825 118.595 210.995 ;
        RECT 118.885 210.825 119.055 210.995 ;
        RECT 119.345 210.825 119.515 210.995 ;
        RECT 119.805 210.825 119.975 210.995 ;
        RECT 120.265 210.825 120.435 210.995 ;
        RECT 120.725 210.825 120.895 210.995 ;
        RECT 121.185 210.825 121.355 210.995 ;
        RECT 121.645 210.825 121.815 210.995 ;
        RECT 67.825 208.105 67.995 208.275 ;
        RECT 68.285 208.105 68.455 208.275 ;
        RECT 68.745 208.105 68.915 208.275 ;
        RECT 69.205 208.105 69.375 208.275 ;
        RECT 69.665 208.105 69.835 208.275 ;
        RECT 70.125 208.105 70.295 208.275 ;
        RECT 70.585 208.105 70.755 208.275 ;
        RECT 71.045 208.105 71.215 208.275 ;
        RECT 71.505 208.105 71.675 208.275 ;
        RECT 71.965 208.105 72.135 208.275 ;
        RECT 72.425 208.105 72.595 208.275 ;
        RECT 72.885 208.105 73.055 208.275 ;
        RECT 73.345 208.105 73.515 208.275 ;
        RECT 73.805 208.105 73.975 208.275 ;
        RECT 74.265 208.105 74.435 208.275 ;
        RECT 74.725 208.105 74.895 208.275 ;
        RECT 75.185 208.105 75.355 208.275 ;
        RECT 75.645 208.105 75.815 208.275 ;
        RECT 76.105 208.105 76.275 208.275 ;
        RECT 76.565 208.105 76.735 208.275 ;
        RECT 77.025 208.105 77.195 208.275 ;
        RECT 77.485 208.105 77.655 208.275 ;
        RECT 77.945 208.105 78.115 208.275 ;
        RECT 78.405 208.105 78.575 208.275 ;
        RECT 78.865 208.105 79.035 208.275 ;
        RECT 79.325 208.105 79.495 208.275 ;
        RECT 79.785 208.105 79.955 208.275 ;
        RECT 80.245 208.105 80.415 208.275 ;
        RECT 80.705 208.105 80.875 208.275 ;
        RECT 81.165 208.105 81.335 208.275 ;
        RECT 81.625 208.105 81.795 208.275 ;
        RECT 82.085 208.105 82.255 208.275 ;
        RECT 82.545 208.105 82.715 208.275 ;
        RECT 83.005 208.105 83.175 208.275 ;
        RECT 83.465 208.105 83.635 208.275 ;
        RECT 83.925 208.105 84.095 208.275 ;
        RECT 84.385 208.105 84.555 208.275 ;
        RECT 84.845 208.105 85.015 208.275 ;
        RECT 85.305 208.105 85.475 208.275 ;
        RECT 85.765 208.105 85.935 208.275 ;
        RECT 86.225 208.105 86.395 208.275 ;
        RECT 86.685 208.105 86.855 208.275 ;
        RECT 87.145 208.105 87.315 208.275 ;
        RECT 87.605 208.105 87.775 208.275 ;
        RECT 88.065 208.105 88.235 208.275 ;
        RECT 88.525 208.105 88.695 208.275 ;
        RECT 88.985 208.105 89.155 208.275 ;
        RECT 89.445 208.105 89.615 208.275 ;
        RECT 89.905 208.105 90.075 208.275 ;
        RECT 90.365 208.105 90.535 208.275 ;
        RECT 90.825 208.105 90.995 208.275 ;
        RECT 91.285 208.105 91.455 208.275 ;
        RECT 91.745 208.105 91.915 208.275 ;
        RECT 92.205 208.105 92.375 208.275 ;
        RECT 92.665 208.105 92.835 208.275 ;
        RECT 93.125 208.105 93.295 208.275 ;
        RECT 93.585 208.105 93.755 208.275 ;
        RECT 94.045 208.105 94.215 208.275 ;
        RECT 94.505 208.105 94.675 208.275 ;
        RECT 94.965 208.105 95.135 208.275 ;
        RECT 95.425 208.105 95.595 208.275 ;
        RECT 95.885 208.105 96.055 208.275 ;
        RECT 96.345 208.105 96.515 208.275 ;
        RECT 96.805 208.105 96.975 208.275 ;
        RECT 97.265 208.105 97.435 208.275 ;
        RECT 97.725 208.105 97.895 208.275 ;
        RECT 98.185 208.105 98.355 208.275 ;
        RECT 98.645 208.105 98.815 208.275 ;
        RECT 99.105 208.105 99.275 208.275 ;
        RECT 99.565 208.105 99.735 208.275 ;
        RECT 100.025 208.105 100.195 208.275 ;
        RECT 100.485 208.105 100.655 208.275 ;
        RECT 100.945 208.105 101.115 208.275 ;
        RECT 101.405 208.105 101.575 208.275 ;
        RECT 101.865 208.105 102.035 208.275 ;
        RECT 102.325 208.105 102.495 208.275 ;
        RECT 102.785 208.105 102.955 208.275 ;
        RECT 103.245 208.105 103.415 208.275 ;
        RECT 103.705 208.105 103.875 208.275 ;
        RECT 104.165 208.105 104.335 208.275 ;
        RECT 104.625 208.105 104.795 208.275 ;
        RECT 105.085 208.105 105.255 208.275 ;
        RECT 105.545 208.105 105.715 208.275 ;
        RECT 106.005 208.105 106.175 208.275 ;
        RECT 106.465 208.105 106.635 208.275 ;
        RECT 106.925 208.105 107.095 208.275 ;
        RECT 107.385 208.105 107.555 208.275 ;
        RECT 107.845 208.105 108.015 208.275 ;
        RECT 108.305 208.105 108.475 208.275 ;
        RECT 108.765 208.105 108.935 208.275 ;
        RECT 109.225 208.105 109.395 208.275 ;
        RECT 109.685 208.105 109.855 208.275 ;
        RECT 110.145 208.105 110.315 208.275 ;
        RECT 110.605 208.105 110.775 208.275 ;
        RECT 111.065 208.105 111.235 208.275 ;
        RECT 111.525 208.105 111.695 208.275 ;
        RECT 111.985 208.105 112.155 208.275 ;
        RECT 112.445 208.105 112.615 208.275 ;
        RECT 112.905 208.105 113.075 208.275 ;
        RECT 113.365 208.105 113.535 208.275 ;
        RECT 113.825 208.105 113.995 208.275 ;
        RECT 114.285 208.105 114.455 208.275 ;
        RECT 114.745 208.105 114.915 208.275 ;
        RECT 115.205 208.105 115.375 208.275 ;
        RECT 115.665 208.105 115.835 208.275 ;
        RECT 116.125 208.105 116.295 208.275 ;
        RECT 116.585 208.105 116.755 208.275 ;
        RECT 117.045 208.105 117.215 208.275 ;
        RECT 117.505 208.105 117.675 208.275 ;
        RECT 117.965 208.105 118.135 208.275 ;
        RECT 118.425 208.105 118.595 208.275 ;
        RECT 118.885 208.105 119.055 208.275 ;
        RECT 119.345 208.105 119.515 208.275 ;
        RECT 119.805 208.105 119.975 208.275 ;
        RECT 120.265 208.105 120.435 208.275 ;
        RECT 120.725 208.105 120.895 208.275 ;
        RECT 121.185 208.105 121.355 208.275 ;
        RECT 121.645 208.105 121.815 208.275 ;
        RECT 67.825 205.385 67.995 205.555 ;
        RECT 68.285 205.385 68.455 205.555 ;
        RECT 68.745 205.385 68.915 205.555 ;
        RECT 69.205 205.385 69.375 205.555 ;
        RECT 69.665 205.385 69.835 205.555 ;
        RECT 70.125 205.385 70.295 205.555 ;
        RECT 70.585 205.385 70.755 205.555 ;
        RECT 71.045 205.385 71.215 205.555 ;
        RECT 71.505 205.385 71.675 205.555 ;
        RECT 71.965 205.385 72.135 205.555 ;
        RECT 72.425 205.385 72.595 205.555 ;
        RECT 72.885 205.385 73.055 205.555 ;
        RECT 73.345 205.385 73.515 205.555 ;
        RECT 73.805 205.385 73.975 205.555 ;
        RECT 74.265 205.385 74.435 205.555 ;
        RECT 74.725 205.385 74.895 205.555 ;
        RECT 75.185 205.385 75.355 205.555 ;
        RECT 75.645 205.385 75.815 205.555 ;
        RECT 76.105 205.385 76.275 205.555 ;
        RECT 76.565 205.385 76.735 205.555 ;
        RECT 77.025 205.385 77.195 205.555 ;
        RECT 77.485 205.385 77.655 205.555 ;
        RECT 77.945 205.385 78.115 205.555 ;
        RECT 78.405 205.385 78.575 205.555 ;
        RECT 78.865 205.385 79.035 205.555 ;
        RECT 79.325 205.385 79.495 205.555 ;
        RECT 79.785 205.385 79.955 205.555 ;
        RECT 80.245 205.385 80.415 205.555 ;
        RECT 80.705 205.385 80.875 205.555 ;
        RECT 81.165 205.385 81.335 205.555 ;
        RECT 81.625 205.385 81.795 205.555 ;
        RECT 82.085 205.385 82.255 205.555 ;
        RECT 82.545 205.385 82.715 205.555 ;
        RECT 83.005 205.385 83.175 205.555 ;
        RECT 83.465 205.385 83.635 205.555 ;
        RECT 83.925 205.385 84.095 205.555 ;
        RECT 84.385 205.385 84.555 205.555 ;
        RECT 84.845 205.385 85.015 205.555 ;
        RECT 85.305 205.385 85.475 205.555 ;
        RECT 85.765 205.385 85.935 205.555 ;
        RECT 86.225 205.385 86.395 205.555 ;
        RECT 86.685 205.385 86.855 205.555 ;
        RECT 87.145 205.385 87.315 205.555 ;
        RECT 87.605 205.385 87.775 205.555 ;
        RECT 88.065 205.385 88.235 205.555 ;
        RECT 88.525 205.385 88.695 205.555 ;
        RECT 88.985 205.385 89.155 205.555 ;
        RECT 89.445 205.385 89.615 205.555 ;
        RECT 89.905 205.385 90.075 205.555 ;
        RECT 90.365 205.385 90.535 205.555 ;
        RECT 90.825 205.385 90.995 205.555 ;
        RECT 91.285 205.385 91.455 205.555 ;
        RECT 91.745 205.385 91.915 205.555 ;
        RECT 92.205 205.385 92.375 205.555 ;
        RECT 92.665 205.385 92.835 205.555 ;
        RECT 93.125 205.385 93.295 205.555 ;
        RECT 93.585 205.385 93.755 205.555 ;
        RECT 94.045 205.385 94.215 205.555 ;
        RECT 94.505 205.385 94.675 205.555 ;
        RECT 94.965 205.385 95.135 205.555 ;
        RECT 95.425 205.385 95.595 205.555 ;
        RECT 95.885 205.385 96.055 205.555 ;
        RECT 96.345 205.385 96.515 205.555 ;
        RECT 96.805 205.385 96.975 205.555 ;
        RECT 97.265 205.385 97.435 205.555 ;
        RECT 97.725 205.385 97.895 205.555 ;
        RECT 98.185 205.385 98.355 205.555 ;
        RECT 98.645 205.385 98.815 205.555 ;
        RECT 99.105 205.385 99.275 205.555 ;
        RECT 99.565 205.385 99.735 205.555 ;
        RECT 100.025 205.385 100.195 205.555 ;
        RECT 100.485 205.385 100.655 205.555 ;
        RECT 100.945 205.385 101.115 205.555 ;
        RECT 101.405 205.385 101.575 205.555 ;
        RECT 101.865 205.385 102.035 205.555 ;
        RECT 102.325 205.385 102.495 205.555 ;
        RECT 102.785 205.385 102.955 205.555 ;
        RECT 103.245 205.385 103.415 205.555 ;
        RECT 103.705 205.385 103.875 205.555 ;
        RECT 104.165 205.385 104.335 205.555 ;
        RECT 104.625 205.385 104.795 205.555 ;
        RECT 105.085 205.385 105.255 205.555 ;
        RECT 105.545 205.385 105.715 205.555 ;
        RECT 106.005 205.385 106.175 205.555 ;
        RECT 106.465 205.385 106.635 205.555 ;
        RECT 106.925 205.385 107.095 205.555 ;
        RECT 107.385 205.385 107.555 205.555 ;
        RECT 107.845 205.385 108.015 205.555 ;
        RECT 108.305 205.385 108.475 205.555 ;
        RECT 108.765 205.385 108.935 205.555 ;
        RECT 109.225 205.385 109.395 205.555 ;
        RECT 109.685 205.385 109.855 205.555 ;
        RECT 110.145 205.385 110.315 205.555 ;
        RECT 110.605 205.385 110.775 205.555 ;
        RECT 111.065 205.385 111.235 205.555 ;
        RECT 111.525 205.385 111.695 205.555 ;
        RECT 111.985 205.385 112.155 205.555 ;
        RECT 112.445 205.385 112.615 205.555 ;
        RECT 112.905 205.385 113.075 205.555 ;
        RECT 113.365 205.385 113.535 205.555 ;
        RECT 113.825 205.385 113.995 205.555 ;
        RECT 114.285 205.385 114.455 205.555 ;
        RECT 114.745 205.385 114.915 205.555 ;
        RECT 115.205 205.385 115.375 205.555 ;
        RECT 115.665 205.385 115.835 205.555 ;
        RECT 116.125 205.385 116.295 205.555 ;
        RECT 116.585 205.385 116.755 205.555 ;
        RECT 117.045 205.385 117.215 205.555 ;
        RECT 117.505 205.385 117.675 205.555 ;
        RECT 117.965 205.385 118.135 205.555 ;
        RECT 118.425 205.385 118.595 205.555 ;
        RECT 118.885 205.385 119.055 205.555 ;
        RECT 119.345 205.385 119.515 205.555 ;
        RECT 119.805 205.385 119.975 205.555 ;
        RECT 120.265 205.385 120.435 205.555 ;
        RECT 120.725 205.385 120.895 205.555 ;
        RECT 121.185 205.385 121.355 205.555 ;
        RECT 121.645 205.385 121.815 205.555 ;
        RECT 67.825 202.665 67.995 202.835 ;
        RECT 68.285 202.665 68.455 202.835 ;
        RECT 68.745 202.665 68.915 202.835 ;
        RECT 69.205 202.665 69.375 202.835 ;
        RECT 69.665 202.665 69.835 202.835 ;
        RECT 70.125 202.665 70.295 202.835 ;
        RECT 70.585 202.665 70.755 202.835 ;
        RECT 71.045 202.665 71.215 202.835 ;
        RECT 71.505 202.665 71.675 202.835 ;
        RECT 71.965 202.665 72.135 202.835 ;
        RECT 72.425 202.665 72.595 202.835 ;
        RECT 72.885 202.665 73.055 202.835 ;
        RECT 73.345 202.665 73.515 202.835 ;
        RECT 73.805 202.665 73.975 202.835 ;
        RECT 74.265 202.665 74.435 202.835 ;
        RECT 74.725 202.665 74.895 202.835 ;
        RECT 75.185 202.665 75.355 202.835 ;
        RECT 75.645 202.665 75.815 202.835 ;
        RECT 76.105 202.665 76.275 202.835 ;
        RECT 76.565 202.665 76.735 202.835 ;
        RECT 77.025 202.665 77.195 202.835 ;
        RECT 77.485 202.665 77.655 202.835 ;
        RECT 77.945 202.665 78.115 202.835 ;
        RECT 78.405 202.665 78.575 202.835 ;
        RECT 78.865 202.665 79.035 202.835 ;
        RECT 79.325 202.665 79.495 202.835 ;
        RECT 79.785 202.665 79.955 202.835 ;
        RECT 80.245 202.665 80.415 202.835 ;
        RECT 80.705 202.665 80.875 202.835 ;
        RECT 81.165 202.665 81.335 202.835 ;
        RECT 81.625 202.665 81.795 202.835 ;
        RECT 82.085 202.665 82.255 202.835 ;
        RECT 82.545 202.665 82.715 202.835 ;
        RECT 83.005 202.665 83.175 202.835 ;
        RECT 83.465 202.665 83.635 202.835 ;
        RECT 83.925 202.665 84.095 202.835 ;
        RECT 84.385 202.665 84.555 202.835 ;
        RECT 84.845 202.665 85.015 202.835 ;
        RECT 85.305 202.665 85.475 202.835 ;
        RECT 85.765 202.665 85.935 202.835 ;
        RECT 86.225 202.665 86.395 202.835 ;
        RECT 86.685 202.665 86.855 202.835 ;
        RECT 87.145 202.665 87.315 202.835 ;
        RECT 87.605 202.665 87.775 202.835 ;
        RECT 88.065 202.665 88.235 202.835 ;
        RECT 88.525 202.665 88.695 202.835 ;
        RECT 88.985 202.665 89.155 202.835 ;
        RECT 89.445 202.665 89.615 202.835 ;
        RECT 89.905 202.665 90.075 202.835 ;
        RECT 90.365 202.665 90.535 202.835 ;
        RECT 90.825 202.665 90.995 202.835 ;
        RECT 91.285 202.665 91.455 202.835 ;
        RECT 91.745 202.665 91.915 202.835 ;
        RECT 92.205 202.665 92.375 202.835 ;
        RECT 92.665 202.665 92.835 202.835 ;
        RECT 93.125 202.665 93.295 202.835 ;
        RECT 93.585 202.665 93.755 202.835 ;
        RECT 94.045 202.665 94.215 202.835 ;
        RECT 94.505 202.665 94.675 202.835 ;
        RECT 94.965 202.665 95.135 202.835 ;
        RECT 95.425 202.665 95.595 202.835 ;
        RECT 95.885 202.665 96.055 202.835 ;
        RECT 96.345 202.665 96.515 202.835 ;
        RECT 96.805 202.665 96.975 202.835 ;
        RECT 97.265 202.665 97.435 202.835 ;
        RECT 97.725 202.665 97.895 202.835 ;
        RECT 98.185 202.665 98.355 202.835 ;
        RECT 98.645 202.665 98.815 202.835 ;
        RECT 99.105 202.665 99.275 202.835 ;
        RECT 99.565 202.665 99.735 202.835 ;
        RECT 100.025 202.665 100.195 202.835 ;
        RECT 100.485 202.665 100.655 202.835 ;
        RECT 100.945 202.665 101.115 202.835 ;
        RECT 101.405 202.665 101.575 202.835 ;
        RECT 101.865 202.665 102.035 202.835 ;
        RECT 102.325 202.665 102.495 202.835 ;
        RECT 102.785 202.665 102.955 202.835 ;
        RECT 103.245 202.665 103.415 202.835 ;
        RECT 103.705 202.665 103.875 202.835 ;
        RECT 104.165 202.665 104.335 202.835 ;
        RECT 104.625 202.665 104.795 202.835 ;
        RECT 105.085 202.665 105.255 202.835 ;
        RECT 105.545 202.665 105.715 202.835 ;
        RECT 106.005 202.665 106.175 202.835 ;
        RECT 106.465 202.665 106.635 202.835 ;
        RECT 106.925 202.665 107.095 202.835 ;
        RECT 107.385 202.665 107.555 202.835 ;
        RECT 107.845 202.665 108.015 202.835 ;
        RECT 108.305 202.665 108.475 202.835 ;
        RECT 108.765 202.665 108.935 202.835 ;
        RECT 109.225 202.665 109.395 202.835 ;
        RECT 109.685 202.665 109.855 202.835 ;
        RECT 110.145 202.665 110.315 202.835 ;
        RECT 110.605 202.665 110.775 202.835 ;
        RECT 111.065 202.665 111.235 202.835 ;
        RECT 111.525 202.665 111.695 202.835 ;
        RECT 111.985 202.665 112.155 202.835 ;
        RECT 112.445 202.665 112.615 202.835 ;
        RECT 112.905 202.665 113.075 202.835 ;
        RECT 113.365 202.665 113.535 202.835 ;
        RECT 113.825 202.665 113.995 202.835 ;
        RECT 114.285 202.665 114.455 202.835 ;
        RECT 114.745 202.665 114.915 202.835 ;
        RECT 115.205 202.665 115.375 202.835 ;
        RECT 115.665 202.665 115.835 202.835 ;
        RECT 116.125 202.665 116.295 202.835 ;
        RECT 116.585 202.665 116.755 202.835 ;
        RECT 117.045 202.665 117.215 202.835 ;
        RECT 117.505 202.665 117.675 202.835 ;
        RECT 117.965 202.665 118.135 202.835 ;
        RECT 118.425 202.665 118.595 202.835 ;
        RECT 118.885 202.665 119.055 202.835 ;
        RECT 119.345 202.665 119.515 202.835 ;
        RECT 119.805 202.665 119.975 202.835 ;
        RECT 120.265 202.665 120.435 202.835 ;
        RECT 120.725 202.665 120.895 202.835 ;
        RECT 121.185 202.665 121.355 202.835 ;
        RECT 121.645 202.665 121.815 202.835 ;
        RECT 67.825 199.945 67.995 200.115 ;
        RECT 68.285 199.945 68.455 200.115 ;
        RECT 68.745 199.945 68.915 200.115 ;
        RECT 69.205 199.945 69.375 200.115 ;
        RECT 69.665 199.945 69.835 200.115 ;
        RECT 70.125 199.945 70.295 200.115 ;
        RECT 70.585 199.945 70.755 200.115 ;
        RECT 71.045 199.945 71.215 200.115 ;
        RECT 71.505 199.945 71.675 200.115 ;
        RECT 71.965 199.945 72.135 200.115 ;
        RECT 72.425 199.945 72.595 200.115 ;
        RECT 72.885 199.945 73.055 200.115 ;
        RECT 73.345 199.945 73.515 200.115 ;
        RECT 73.805 199.945 73.975 200.115 ;
        RECT 74.265 199.945 74.435 200.115 ;
        RECT 74.725 199.945 74.895 200.115 ;
        RECT 75.185 199.945 75.355 200.115 ;
        RECT 75.645 199.945 75.815 200.115 ;
        RECT 76.105 199.945 76.275 200.115 ;
        RECT 76.565 199.945 76.735 200.115 ;
        RECT 77.025 199.945 77.195 200.115 ;
        RECT 77.485 199.945 77.655 200.115 ;
        RECT 77.945 199.945 78.115 200.115 ;
        RECT 78.405 199.945 78.575 200.115 ;
        RECT 78.865 199.945 79.035 200.115 ;
        RECT 79.325 199.945 79.495 200.115 ;
        RECT 79.785 199.945 79.955 200.115 ;
        RECT 80.245 199.945 80.415 200.115 ;
        RECT 80.705 199.945 80.875 200.115 ;
        RECT 81.165 199.945 81.335 200.115 ;
        RECT 81.625 199.945 81.795 200.115 ;
        RECT 82.085 199.945 82.255 200.115 ;
        RECT 82.545 199.945 82.715 200.115 ;
        RECT 83.005 199.945 83.175 200.115 ;
        RECT 83.465 199.945 83.635 200.115 ;
        RECT 83.925 199.945 84.095 200.115 ;
        RECT 84.385 199.945 84.555 200.115 ;
        RECT 84.845 199.945 85.015 200.115 ;
        RECT 85.305 199.945 85.475 200.115 ;
        RECT 85.765 199.945 85.935 200.115 ;
        RECT 86.225 199.945 86.395 200.115 ;
        RECT 86.685 199.945 86.855 200.115 ;
        RECT 87.145 199.945 87.315 200.115 ;
        RECT 87.605 199.945 87.775 200.115 ;
        RECT 88.065 199.945 88.235 200.115 ;
        RECT 88.525 199.945 88.695 200.115 ;
        RECT 88.985 199.945 89.155 200.115 ;
        RECT 89.445 199.945 89.615 200.115 ;
        RECT 89.905 199.945 90.075 200.115 ;
        RECT 90.365 199.945 90.535 200.115 ;
        RECT 90.825 199.945 90.995 200.115 ;
        RECT 91.285 199.945 91.455 200.115 ;
        RECT 91.745 199.945 91.915 200.115 ;
        RECT 92.205 199.945 92.375 200.115 ;
        RECT 92.665 199.945 92.835 200.115 ;
        RECT 93.125 199.945 93.295 200.115 ;
        RECT 93.585 199.945 93.755 200.115 ;
        RECT 94.045 199.945 94.215 200.115 ;
        RECT 94.505 199.945 94.675 200.115 ;
        RECT 94.965 199.945 95.135 200.115 ;
        RECT 95.425 199.945 95.595 200.115 ;
        RECT 95.885 199.945 96.055 200.115 ;
        RECT 96.345 199.945 96.515 200.115 ;
        RECT 96.805 199.945 96.975 200.115 ;
        RECT 97.265 199.945 97.435 200.115 ;
        RECT 97.725 199.945 97.895 200.115 ;
        RECT 98.185 199.945 98.355 200.115 ;
        RECT 98.645 199.945 98.815 200.115 ;
        RECT 99.105 199.945 99.275 200.115 ;
        RECT 99.565 199.945 99.735 200.115 ;
        RECT 100.025 199.945 100.195 200.115 ;
        RECT 100.485 199.945 100.655 200.115 ;
        RECT 100.945 199.945 101.115 200.115 ;
        RECT 101.405 199.945 101.575 200.115 ;
        RECT 101.865 199.945 102.035 200.115 ;
        RECT 102.325 199.945 102.495 200.115 ;
        RECT 102.785 199.945 102.955 200.115 ;
        RECT 103.245 199.945 103.415 200.115 ;
        RECT 103.705 199.945 103.875 200.115 ;
        RECT 104.165 199.945 104.335 200.115 ;
        RECT 104.625 199.945 104.795 200.115 ;
        RECT 105.085 199.945 105.255 200.115 ;
        RECT 105.545 199.945 105.715 200.115 ;
        RECT 106.005 199.945 106.175 200.115 ;
        RECT 106.465 199.945 106.635 200.115 ;
        RECT 106.925 199.945 107.095 200.115 ;
        RECT 107.385 199.945 107.555 200.115 ;
        RECT 107.845 199.945 108.015 200.115 ;
        RECT 108.305 199.945 108.475 200.115 ;
        RECT 108.765 199.945 108.935 200.115 ;
        RECT 109.225 199.945 109.395 200.115 ;
        RECT 109.685 199.945 109.855 200.115 ;
        RECT 110.145 199.945 110.315 200.115 ;
        RECT 110.605 199.945 110.775 200.115 ;
        RECT 111.065 199.945 111.235 200.115 ;
        RECT 111.525 199.945 111.695 200.115 ;
        RECT 111.985 199.945 112.155 200.115 ;
        RECT 112.445 199.945 112.615 200.115 ;
        RECT 112.905 199.945 113.075 200.115 ;
        RECT 113.365 199.945 113.535 200.115 ;
        RECT 113.825 199.945 113.995 200.115 ;
        RECT 114.285 199.945 114.455 200.115 ;
        RECT 114.745 199.945 114.915 200.115 ;
        RECT 115.205 199.945 115.375 200.115 ;
        RECT 115.665 199.945 115.835 200.115 ;
        RECT 116.125 199.945 116.295 200.115 ;
        RECT 116.585 199.945 116.755 200.115 ;
        RECT 117.045 199.945 117.215 200.115 ;
        RECT 117.505 199.945 117.675 200.115 ;
        RECT 117.965 199.945 118.135 200.115 ;
        RECT 118.425 199.945 118.595 200.115 ;
        RECT 118.885 199.945 119.055 200.115 ;
        RECT 119.345 199.945 119.515 200.115 ;
        RECT 119.805 199.945 119.975 200.115 ;
        RECT 120.265 199.945 120.435 200.115 ;
        RECT 120.725 199.945 120.895 200.115 ;
        RECT 121.185 199.945 121.355 200.115 ;
        RECT 121.645 199.945 121.815 200.115 ;
        RECT 67.825 197.225 67.995 197.395 ;
        RECT 68.285 197.225 68.455 197.395 ;
        RECT 68.745 197.225 68.915 197.395 ;
        RECT 69.205 197.225 69.375 197.395 ;
        RECT 69.665 197.225 69.835 197.395 ;
        RECT 70.125 197.225 70.295 197.395 ;
        RECT 70.585 197.225 70.755 197.395 ;
        RECT 71.045 197.225 71.215 197.395 ;
        RECT 71.505 197.225 71.675 197.395 ;
        RECT 71.965 197.225 72.135 197.395 ;
        RECT 72.425 197.225 72.595 197.395 ;
        RECT 72.885 197.225 73.055 197.395 ;
        RECT 73.345 197.225 73.515 197.395 ;
        RECT 73.805 197.225 73.975 197.395 ;
        RECT 74.265 197.225 74.435 197.395 ;
        RECT 74.725 197.225 74.895 197.395 ;
        RECT 75.185 197.225 75.355 197.395 ;
        RECT 75.645 197.225 75.815 197.395 ;
        RECT 76.105 197.225 76.275 197.395 ;
        RECT 76.565 197.225 76.735 197.395 ;
        RECT 77.025 197.225 77.195 197.395 ;
        RECT 77.485 197.225 77.655 197.395 ;
        RECT 77.945 197.225 78.115 197.395 ;
        RECT 78.405 197.225 78.575 197.395 ;
        RECT 78.865 197.225 79.035 197.395 ;
        RECT 79.325 197.225 79.495 197.395 ;
        RECT 79.785 197.225 79.955 197.395 ;
        RECT 80.245 197.225 80.415 197.395 ;
        RECT 80.705 197.225 80.875 197.395 ;
        RECT 81.165 197.225 81.335 197.395 ;
        RECT 81.625 197.225 81.795 197.395 ;
        RECT 82.085 197.225 82.255 197.395 ;
        RECT 82.545 197.225 82.715 197.395 ;
        RECT 83.005 197.225 83.175 197.395 ;
        RECT 83.465 197.225 83.635 197.395 ;
        RECT 83.925 197.225 84.095 197.395 ;
        RECT 84.385 197.225 84.555 197.395 ;
        RECT 84.845 197.225 85.015 197.395 ;
        RECT 85.305 197.225 85.475 197.395 ;
        RECT 85.765 197.225 85.935 197.395 ;
        RECT 86.225 197.225 86.395 197.395 ;
        RECT 86.685 197.225 86.855 197.395 ;
        RECT 87.145 197.225 87.315 197.395 ;
        RECT 87.605 197.225 87.775 197.395 ;
        RECT 88.065 197.225 88.235 197.395 ;
        RECT 88.525 197.225 88.695 197.395 ;
        RECT 88.985 197.225 89.155 197.395 ;
        RECT 89.445 197.225 89.615 197.395 ;
        RECT 89.905 197.225 90.075 197.395 ;
        RECT 90.365 197.225 90.535 197.395 ;
        RECT 90.825 197.225 90.995 197.395 ;
        RECT 91.285 197.225 91.455 197.395 ;
        RECT 91.745 197.225 91.915 197.395 ;
        RECT 92.205 197.225 92.375 197.395 ;
        RECT 92.665 197.225 92.835 197.395 ;
        RECT 93.125 197.225 93.295 197.395 ;
        RECT 93.585 197.225 93.755 197.395 ;
        RECT 94.045 197.225 94.215 197.395 ;
        RECT 94.505 197.225 94.675 197.395 ;
        RECT 94.965 197.225 95.135 197.395 ;
        RECT 95.425 197.225 95.595 197.395 ;
        RECT 95.885 197.225 96.055 197.395 ;
        RECT 96.345 197.225 96.515 197.395 ;
        RECT 96.805 197.225 96.975 197.395 ;
        RECT 97.265 197.225 97.435 197.395 ;
        RECT 97.725 197.225 97.895 197.395 ;
        RECT 98.185 197.225 98.355 197.395 ;
        RECT 98.645 197.225 98.815 197.395 ;
        RECT 99.105 197.225 99.275 197.395 ;
        RECT 99.565 197.225 99.735 197.395 ;
        RECT 100.025 197.225 100.195 197.395 ;
        RECT 100.485 197.225 100.655 197.395 ;
        RECT 100.945 197.225 101.115 197.395 ;
        RECT 101.405 197.225 101.575 197.395 ;
        RECT 101.865 197.225 102.035 197.395 ;
        RECT 102.325 197.225 102.495 197.395 ;
        RECT 102.785 197.225 102.955 197.395 ;
        RECT 103.245 197.225 103.415 197.395 ;
        RECT 103.705 197.225 103.875 197.395 ;
        RECT 104.165 197.225 104.335 197.395 ;
        RECT 104.625 197.225 104.795 197.395 ;
        RECT 105.085 197.225 105.255 197.395 ;
        RECT 105.545 197.225 105.715 197.395 ;
        RECT 106.005 197.225 106.175 197.395 ;
        RECT 106.465 197.225 106.635 197.395 ;
        RECT 106.925 197.225 107.095 197.395 ;
        RECT 107.385 197.225 107.555 197.395 ;
        RECT 107.845 197.225 108.015 197.395 ;
        RECT 108.305 197.225 108.475 197.395 ;
        RECT 108.765 197.225 108.935 197.395 ;
        RECT 109.225 197.225 109.395 197.395 ;
        RECT 109.685 197.225 109.855 197.395 ;
        RECT 110.145 197.225 110.315 197.395 ;
        RECT 110.605 197.225 110.775 197.395 ;
        RECT 111.065 197.225 111.235 197.395 ;
        RECT 111.525 197.225 111.695 197.395 ;
        RECT 111.985 197.225 112.155 197.395 ;
        RECT 112.445 197.225 112.615 197.395 ;
        RECT 112.905 197.225 113.075 197.395 ;
        RECT 113.365 197.225 113.535 197.395 ;
        RECT 113.825 197.225 113.995 197.395 ;
        RECT 114.285 197.225 114.455 197.395 ;
        RECT 114.745 197.225 114.915 197.395 ;
        RECT 115.205 197.225 115.375 197.395 ;
        RECT 115.665 197.225 115.835 197.395 ;
        RECT 116.125 197.225 116.295 197.395 ;
        RECT 116.585 197.225 116.755 197.395 ;
        RECT 117.045 197.225 117.215 197.395 ;
        RECT 117.505 197.225 117.675 197.395 ;
        RECT 117.965 197.225 118.135 197.395 ;
        RECT 118.425 197.225 118.595 197.395 ;
        RECT 118.885 197.225 119.055 197.395 ;
        RECT 119.345 197.225 119.515 197.395 ;
        RECT 119.805 197.225 119.975 197.395 ;
        RECT 120.265 197.225 120.435 197.395 ;
        RECT 120.725 197.225 120.895 197.395 ;
        RECT 121.185 197.225 121.355 197.395 ;
        RECT 121.645 197.225 121.815 197.395 ;
        RECT 67.825 194.505 67.995 194.675 ;
        RECT 68.285 194.505 68.455 194.675 ;
        RECT 68.745 194.505 68.915 194.675 ;
        RECT 69.205 194.505 69.375 194.675 ;
        RECT 69.665 194.505 69.835 194.675 ;
        RECT 70.125 194.505 70.295 194.675 ;
        RECT 70.585 194.505 70.755 194.675 ;
        RECT 71.045 194.505 71.215 194.675 ;
        RECT 71.505 194.505 71.675 194.675 ;
        RECT 71.965 194.505 72.135 194.675 ;
        RECT 72.425 194.505 72.595 194.675 ;
        RECT 72.885 194.505 73.055 194.675 ;
        RECT 73.345 194.505 73.515 194.675 ;
        RECT 73.805 194.505 73.975 194.675 ;
        RECT 74.265 194.505 74.435 194.675 ;
        RECT 74.725 194.505 74.895 194.675 ;
        RECT 75.185 194.505 75.355 194.675 ;
        RECT 75.645 194.505 75.815 194.675 ;
        RECT 76.105 194.505 76.275 194.675 ;
        RECT 76.565 194.505 76.735 194.675 ;
        RECT 77.025 194.505 77.195 194.675 ;
        RECT 77.485 194.505 77.655 194.675 ;
        RECT 77.945 194.505 78.115 194.675 ;
        RECT 78.405 194.505 78.575 194.675 ;
        RECT 78.865 194.505 79.035 194.675 ;
        RECT 79.325 194.505 79.495 194.675 ;
        RECT 79.785 194.505 79.955 194.675 ;
        RECT 80.245 194.505 80.415 194.675 ;
        RECT 80.705 194.505 80.875 194.675 ;
        RECT 81.165 194.505 81.335 194.675 ;
        RECT 81.625 194.505 81.795 194.675 ;
        RECT 82.085 194.505 82.255 194.675 ;
        RECT 82.545 194.505 82.715 194.675 ;
        RECT 83.005 194.505 83.175 194.675 ;
        RECT 83.465 194.505 83.635 194.675 ;
        RECT 83.925 194.505 84.095 194.675 ;
        RECT 84.385 194.505 84.555 194.675 ;
        RECT 84.845 194.505 85.015 194.675 ;
        RECT 85.305 194.505 85.475 194.675 ;
        RECT 85.765 194.505 85.935 194.675 ;
        RECT 86.225 194.505 86.395 194.675 ;
        RECT 86.685 194.505 86.855 194.675 ;
        RECT 87.145 194.505 87.315 194.675 ;
        RECT 87.605 194.505 87.775 194.675 ;
        RECT 88.065 194.505 88.235 194.675 ;
        RECT 88.525 194.505 88.695 194.675 ;
        RECT 88.985 194.505 89.155 194.675 ;
        RECT 89.445 194.505 89.615 194.675 ;
        RECT 89.905 194.505 90.075 194.675 ;
        RECT 90.365 194.505 90.535 194.675 ;
        RECT 90.825 194.505 90.995 194.675 ;
        RECT 91.285 194.505 91.455 194.675 ;
        RECT 91.745 194.505 91.915 194.675 ;
        RECT 92.205 194.505 92.375 194.675 ;
        RECT 92.665 194.505 92.835 194.675 ;
        RECT 93.125 194.505 93.295 194.675 ;
        RECT 93.585 194.505 93.755 194.675 ;
        RECT 94.045 194.505 94.215 194.675 ;
        RECT 94.505 194.505 94.675 194.675 ;
        RECT 94.965 194.505 95.135 194.675 ;
        RECT 95.425 194.505 95.595 194.675 ;
        RECT 95.885 194.505 96.055 194.675 ;
        RECT 96.345 194.505 96.515 194.675 ;
        RECT 96.805 194.505 96.975 194.675 ;
        RECT 97.265 194.505 97.435 194.675 ;
        RECT 97.725 194.505 97.895 194.675 ;
        RECT 98.185 194.505 98.355 194.675 ;
        RECT 98.645 194.505 98.815 194.675 ;
        RECT 99.105 194.505 99.275 194.675 ;
        RECT 99.565 194.505 99.735 194.675 ;
        RECT 100.025 194.505 100.195 194.675 ;
        RECT 100.485 194.505 100.655 194.675 ;
        RECT 100.945 194.505 101.115 194.675 ;
        RECT 101.405 194.505 101.575 194.675 ;
        RECT 101.865 194.505 102.035 194.675 ;
        RECT 102.325 194.505 102.495 194.675 ;
        RECT 102.785 194.505 102.955 194.675 ;
        RECT 103.245 194.505 103.415 194.675 ;
        RECT 103.705 194.505 103.875 194.675 ;
        RECT 104.165 194.505 104.335 194.675 ;
        RECT 104.625 194.505 104.795 194.675 ;
        RECT 105.085 194.505 105.255 194.675 ;
        RECT 105.545 194.505 105.715 194.675 ;
        RECT 106.005 194.505 106.175 194.675 ;
        RECT 106.465 194.505 106.635 194.675 ;
        RECT 106.925 194.505 107.095 194.675 ;
        RECT 107.385 194.505 107.555 194.675 ;
        RECT 107.845 194.505 108.015 194.675 ;
        RECT 108.305 194.505 108.475 194.675 ;
        RECT 108.765 194.505 108.935 194.675 ;
        RECT 109.225 194.505 109.395 194.675 ;
        RECT 109.685 194.505 109.855 194.675 ;
        RECT 110.145 194.505 110.315 194.675 ;
        RECT 110.605 194.505 110.775 194.675 ;
        RECT 111.065 194.505 111.235 194.675 ;
        RECT 111.525 194.505 111.695 194.675 ;
        RECT 111.985 194.505 112.155 194.675 ;
        RECT 112.445 194.505 112.615 194.675 ;
        RECT 112.905 194.505 113.075 194.675 ;
        RECT 113.365 194.505 113.535 194.675 ;
        RECT 113.825 194.505 113.995 194.675 ;
        RECT 114.285 194.505 114.455 194.675 ;
        RECT 114.745 194.505 114.915 194.675 ;
        RECT 115.205 194.505 115.375 194.675 ;
        RECT 115.665 194.505 115.835 194.675 ;
        RECT 116.125 194.505 116.295 194.675 ;
        RECT 116.585 194.505 116.755 194.675 ;
        RECT 117.045 194.505 117.215 194.675 ;
        RECT 117.505 194.505 117.675 194.675 ;
        RECT 117.965 194.505 118.135 194.675 ;
        RECT 118.425 194.505 118.595 194.675 ;
        RECT 118.885 194.505 119.055 194.675 ;
        RECT 119.345 194.505 119.515 194.675 ;
        RECT 119.805 194.505 119.975 194.675 ;
        RECT 120.265 194.505 120.435 194.675 ;
        RECT 120.725 194.505 120.895 194.675 ;
        RECT 121.185 194.505 121.355 194.675 ;
        RECT 121.645 194.505 121.815 194.675 ;
        RECT 67.825 191.785 67.995 191.955 ;
        RECT 68.285 191.785 68.455 191.955 ;
        RECT 68.745 191.785 68.915 191.955 ;
        RECT 69.205 191.785 69.375 191.955 ;
        RECT 69.665 191.785 69.835 191.955 ;
        RECT 70.125 191.785 70.295 191.955 ;
        RECT 70.585 191.785 70.755 191.955 ;
        RECT 71.045 191.785 71.215 191.955 ;
        RECT 71.505 191.785 71.675 191.955 ;
        RECT 71.965 191.785 72.135 191.955 ;
        RECT 72.425 191.785 72.595 191.955 ;
        RECT 72.885 191.785 73.055 191.955 ;
        RECT 73.345 191.785 73.515 191.955 ;
        RECT 73.805 191.785 73.975 191.955 ;
        RECT 74.265 191.785 74.435 191.955 ;
        RECT 74.725 191.785 74.895 191.955 ;
        RECT 75.185 191.785 75.355 191.955 ;
        RECT 75.645 191.785 75.815 191.955 ;
        RECT 76.105 191.785 76.275 191.955 ;
        RECT 76.565 191.785 76.735 191.955 ;
        RECT 77.025 191.785 77.195 191.955 ;
        RECT 77.485 191.785 77.655 191.955 ;
        RECT 77.945 191.785 78.115 191.955 ;
        RECT 78.405 191.785 78.575 191.955 ;
        RECT 78.865 191.785 79.035 191.955 ;
        RECT 79.325 191.785 79.495 191.955 ;
        RECT 79.785 191.785 79.955 191.955 ;
        RECT 80.245 191.785 80.415 191.955 ;
        RECT 80.705 191.785 80.875 191.955 ;
        RECT 81.165 191.785 81.335 191.955 ;
        RECT 81.625 191.785 81.795 191.955 ;
        RECT 82.085 191.785 82.255 191.955 ;
        RECT 82.545 191.785 82.715 191.955 ;
        RECT 83.005 191.785 83.175 191.955 ;
        RECT 83.465 191.785 83.635 191.955 ;
        RECT 83.925 191.785 84.095 191.955 ;
        RECT 84.385 191.785 84.555 191.955 ;
        RECT 84.845 191.785 85.015 191.955 ;
        RECT 85.305 191.785 85.475 191.955 ;
        RECT 85.765 191.785 85.935 191.955 ;
        RECT 86.225 191.785 86.395 191.955 ;
        RECT 86.685 191.785 86.855 191.955 ;
        RECT 87.145 191.785 87.315 191.955 ;
        RECT 87.605 191.785 87.775 191.955 ;
        RECT 88.065 191.785 88.235 191.955 ;
        RECT 88.525 191.785 88.695 191.955 ;
        RECT 88.985 191.785 89.155 191.955 ;
        RECT 89.445 191.785 89.615 191.955 ;
        RECT 89.905 191.785 90.075 191.955 ;
        RECT 90.365 191.785 90.535 191.955 ;
        RECT 90.825 191.785 90.995 191.955 ;
        RECT 91.285 191.785 91.455 191.955 ;
        RECT 91.745 191.785 91.915 191.955 ;
        RECT 92.205 191.785 92.375 191.955 ;
        RECT 92.665 191.785 92.835 191.955 ;
        RECT 93.125 191.785 93.295 191.955 ;
        RECT 93.585 191.785 93.755 191.955 ;
        RECT 94.045 191.785 94.215 191.955 ;
        RECT 94.505 191.785 94.675 191.955 ;
        RECT 94.965 191.785 95.135 191.955 ;
        RECT 95.425 191.785 95.595 191.955 ;
        RECT 95.885 191.785 96.055 191.955 ;
        RECT 96.345 191.785 96.515 191.955 ;
        RECT 96.805 191.785 96.975 191.955 ;
        RECT 97.265 191.785 97.435 191.955 ;
        RECT 97.725 191.785 97.895 191.955 ;
        RECT 98.185 191.785 98.355 191.955 ;
        RECT 98.645 191.785 98.815 191.955 ;
        RECT 99.105 191.785 99.275 191.955 ;
        RECT 99.565 191.785 99.735 191.955 ;
        RECT 100.025 191.785 100.195 191.955 ;
        RECT 100.485 191.785 100.655 191.955 ;
        RECT 100.945 191.785 101.115 191.955 ;
        RECT 101.405 191.785 101.575 191.955 ;
        RECT 101.865 191.785 102.035 191.955 ;
        RECT 102.325 191.785 102.495 191.955 ;
        RECT 102.785 191.785 102.955 191.955 ;
        RECT 103.245 191.785 103.415 191.955 ;
        RECT 103.705 191.785 103.875 191.955 ;
        RECT 104.165 191.785 104.335 191.955 ;
        RECT 104.625 191.785 104.795 191.955 ;
        RECT 105.085 191.785 105.255 191.955 ;
        RECT 105.545 191.785 105.715 191.955 ;
        RECT 106.005 191.785 106.175 191.955 ;
        RECT 106.465 191.785 106.635 191.955 ;
        RECT 106.925 191.785 107.095 191.955 ;
        RECT 107.385 191.785 107.555 191.955 ;
        RECT 107.845 191.785 108.015 191.955 ;
        RECT 108.305 191.785 108.475 191.955 ;
        RECT 108.765 191.785 108.935 191.955 ;
        RECT 109.225 191.785 109.395 191.955 ;
        RECT 109.685 191.785 109.855 191.955 ;
        RECT 110.145 191.785 110.315 191.955 ;
        RECT 110.605 191.785 110.775 191.955 ;
        RECT 111.065 191.785 111.235 191.955 ;
        RECT 111.525 191.785 111.695 191.955 ;
        RECT 111.985 191.785 112.155 191.955 ;
        RECT 112.445 191.785 112.615 191.955 ;
        RECT 112.905 191.785 113.075 191.955 ;
        RECT 113.365 191.785 113.535 191.955 ;
        RECT 113.825 191.785 113.995 191.955 ;
        RECT 114.285 191.785 114.455 191.955 ;
        RECT 114.745 191.785 114.915 191.955 ;
        RECT 115.205 191.785 115.375 191.955 ;
        RECT 115.665 191.785 115.835 191.955 ;
        RECT 116.125 191.785 116.295 191.955 ;
        RECT 116.585 191.785 116.755 191.955 ;
        RECT 117.045 191.785 117.215 191.955 ;
        RECT 117.505 191.785 117.675 191.955 ;
        RECT 117.965 191.785 118.135 191.955 ;
        RECT 118.425 191.785 118.595 191.955 ;
        RECT 118.885 191.785 119.055 191.955 ;
        RECT 119.345 191.785 119.515 191.955 ;
        RECT 119.805 191.785 119.975 191.955 ;
        RECT 120.265 191.785 120.435 191.955 ;
        RECT 120.725 191.785 120.895 191.955 ;
        RECT 121.185 191.785 121.355 191.955 ;
        RECT 121.645 191.785 121.815 191.955 ;
        RECT 67.825 189.065 67.995 189.235 ;
        RECT 68.285 189.065 68.455 189.235 ;
        RECT 68.745 189.065 68.915 189.235 ;
        RECT 69.205 189.065 69.375 189.235 ;
        RECT 69.665 189.065 69.835 189.235 ;
        RECT 70.125 189.065 70.295 189.235 ;
        RECT 70.585 189.065 70.755 189.235 ;
        RECT 71.045 189.065 71.215 189.235 ;
        RECT 71.505 189.065 71.675 189.235 ;
        RECT 71.965 189.065 72.135 189.235 ;
        RECT 72.425 189.065 72.595 189.235 ;
        RECT 72.885 189.065 73.055 189.235 ;
        RECT 73.345 189.065 73.515 189.235 ;
        RECT 73.805 189.065 73.975 189.235 ;
        RECT 74.265 189.065 74.435 189.235 ;
        RECT 74.725 189.065 74.895 189.235 ;
        RECT 75.185 189.065 75.355 189.235 ;
        RECT 75.645 189.065 75.815 189.235 ;
        RECT 76.105 189.065 76.275 189.235 ;
        RECT 76.565 189.065 76.735 189.235 ;
        RECT 77.025 189.065 77.195 189.235 ;
        RECT 77.485 189.065 77.655 189.235 ;
        RECT 77.945 189.065 78.115 189.235 ;
        RECT 78.405 189.065 78.575 189.235 ;
        RECT 78.865 189.065 79.035 189.235 ;
        RECT 79.325 189.065 79.495 189.235 ;
        RECT 79.785 189.065 79.955 189.235 ;
        RECT 80.245 189.065 80.415 189.235 ;
        RECT 80.705 189.065 80.875 189.235 ;
        RECT 81.165 189.065 81.335 189.235 ;
        RECT 81.625 189.065 81.795 189.235 ;
        RECT 82.085 189.065 82.255 189.235 ;
        RECT 82.545 189.065 82.715 189.235 ;
        RECT 83.005 189.065 83.175 189.235 ;
        RECT 83.465 189.065 83.635 189.235 ;
        RECT 83.925 189.065 84.095 189.235 ;
        RECT 84.385 189.065 84.555 189.235 ;
        RECT 84.845 189.065 85.015 189.235 ;
        RECT 85.305 189.065 85.475 189.235 ;
        RECT 85.765 189.065 85.935 189.235 ;
        RECT 86.225 189.065 86.395 189.235 ;
        RECT 86.685 189.065 86.855 189.235 ;
        RECT 87.145 189.065 87.315 189.235 ;
        RECT 87.605 189.065 87.775 189.235 ;
        RECT 88.065 189.065 88.235 189.235 ;
        RECT 88.525 189.065 88.695 189.235 ;
        RECT 88.985 189.065 89.155 189.235 ;
        RECT 89.445 189.065 89.615 189.235 ;
        RECT 89.905 189.065 90.075 189.235 ;
        RECT 90.365 189.065 90.535 189.235 ;
        RECT 90.825 189.065 90.995 189.235 ;
        RECT 91.285 189.065 91.455 189.235 ;
        RECT 91.745 189.065 91.915 189.235 ;
        RECT 92.205 189.065 92.375 189.235 ;
        RECT 92.665 189.065 92.835 189.235 ;
        RECT 93.125 189.065 93.295 189.235 ;
        RECT 93.585 189.065 93.755 189.235 ;
        RECT 94.045 189.065 94.215 189.235 ;
        RECT 94.505 189.065 94.675 189.235 ;
        RECT 94.965 189.065 95.135 189.235 ;
        RECT 95.425 189.065 95.595 189.235 ;
        RECT 95.885 189.065 96.055 189.235 ;
        RECT 96.345 189.065 96.515 189.235 ;
        RECT 96.805 189.065 96.975 189.235 ;
        RECT 97.265 189.065 97.435 189.235 ;
        RECT 97.725 189.065 97.895 189.235 ;
        RECT 98.185 189.065 98.355 189.235 ;
        RECT 98.645 189.065 98.815 189.235 ;
        RECT 99.105 189.065 99.275 189.235 ;
        RECT 99.565 189.065 99.735 189.235 ;
        RECT 100.025 189.065 100.195 189.235 ;
        RECT 100.485 189.065 100.655 189.235 ;
        RECT 100.945 189.065 101.115 189.235 ;
        RECT 101.405 189.065 101.575 189.235 ;
        RECT 101.865 189.065 102.035 189.235 ;
        RECT 102.325 189.065 102.495 189.235 ;
        RECT 102.785 189.065 102.955 189.235 ;
        RECT 103.245 189.065 103.415 189.235 ;
        RECT 103.705 189.065 103.875 189.235 ;
        RECT 104.165 189.065 104.335 189.235 ;
        RECT 104.625 189.065 104.795 189.235 ;
        RECT 105.085 189.065 105.255 189.235 ;
        RECT 105.545 189.065 105.715 189.235 ;
        RECT 106.005 189.065 106.175 189.235 ;
        RECT 106.465 189.065 106.635 189.235 ;
        RECT 106.925 189.065 107.095 189.235 ;
        RECT 107.385 189.065 107.555 189.235 ;
        RECT 107.845 189.065 108.015 189.235 ;
        RECT 108.305 189.065 108.475 189.235 ;
        RECT 108.765 189.065 108.935 189.235 ;
        RECT 109.225 189.065 109.395 189.235 ;
        RECT 109.685 189.065 109.855 189.235 ;
        RECT 110.145 189.065 110.315 189.235 ;
        RECT 110.605 189.065 110.775 189.235 ;
        RECT 111.065 189.065 111.235 189.235 ;
        RECT 111.525 189.065 111.695 189.235 ;
        RECT 111.985 189.065 112.155 189.235 ;
        RECT 112.445 189.065 112.615 189.235 ;
        RECT 112.905 189.065 113.075 189.235 ;
        RECT 113.365 189.065 113.535 189.235 ;
        RECT 113.825 189.065 113.995 189.235 ;
        RECT 114.285 189.065 114.455 189.235 ;
        RECT 114.745 189.065 114.915 189.235 ;
        RECT 115.205 189.065 115.375 189.235 ;
        RECT 115.665 189.065 115.835 189.235 ;
        RECT 116.125 189.065 116.295 189.235 ;
        RECT 116.585 189.065 116.755 189.235 ;
        RECT 117.045 189.065 117.215 189.235 ;
        RECT 117.505 189.065 117.675 189.235 ;
        RECT 117.965 189.065 118.135 189.235 ;
        RECT 118.425 189.065 118.595 189.235 ;
        RECT 118.885 189.065 119.055 189.235 ;
        RECT 119.345 189.065 119.515 189.235 ;
        RECT 119.805 189.065 119.975 189.235 ;
        RECT 120.265 189.065 120.435 189.235 ;
        RECT 120.725 189.065 120.895 189.235 ;
        RECT 121.185 189.065 121.355 189.235 ;
        RECT 121.645 189.065 121.815 189.235 ;
        RECT 67.825 186.345 67.995 186.515 ;
        RECT 68.285 186.345 68.455 186.515 ;
        RECT 68.745 186.345 68.915 186.515 ;
        RECT 69.205 186.345 69.375 186.515 ;
        RECT 69.665 186.345 69.835 186.515 ;
        RECT 70.125 186.345 70.295 186.515 ;
        RECT 70.585 186.345 70.755 186.515 ;
        RECT 71.045 186.345 71.215 186.515 ;
        RECT 71.505 186.345 71.675 186.515 ;
        RECT 71.965 186.345 72.135 186.515 ;
        RECT 72.425 186.345 72.595 186.515 ;
        RECT 72.885 186.345 73.055 186.515 ;
        RECT 73.345 186.345 73.515 186.515 ;
        RECT 73.805 186.345 73.975 186.515 ;
        RECT 74.265 186.345 74.435 186.515 ;
        RECT 74.725 186.345 74.895 186.515 ;
        RECT 75.185 186.345 75.355 186.515 ;
        RECT 75.645 186.345 75.815 186.515 ;
        RECT 76.105 186.345 76.275 186.515 ;
        RECT 76.565 186.345 76.735 186.515 ;
        RECT 77.025 186.345 77.195 186.515 ;
        RECT 77.485 186.345 77.655 186.515 ;
        RECT 77.945 186.345 78.115 186.515 ;
        RECT 78.405 186.345 78.575 186.515 ;
        RECT 78.865 186.345 79.035 186.515 ;
        RECT 79.325 186.345 79.495 186.515 ;
        RECT 79.785 186.345 79.955 186.515 ;
        RECT 80.245 186.345 80.415 186.515 ;
        RECT 80.705 186.345 80.875 186.515 ;
        RECT 81.165 186.345 81.335 186.515 ;
        RECT 81.625 186.345 81.795 186.515 ;
        RECT 82.085 186.345 82.255 186.515 ;
        RECT 82.545 186.345 82.715 186.515 ;
        RECT 83.005 186.345 83.175 186.515 ;
        RECT 83.465 186.345 83.635 186.515 ;
        RECT 83.925 186.345 84.095 186.515 ;
        RECT 84.385 186.345 84.555 186.515 ;
        RECT 84.845 186.345 85.015 186.515 ;
        RECT 85.305 186.345 85.475 186.515 ;
        RECT 85.765 186.345 85.935 186.515 ;
        RECT 86.225 186.345 86.395 186.515 ;
        RECT 86.685 186.345 86.855 186.515 ;
        RECT 87.145 186.345 87.315 186.515 ;
        RECT 87.605 186.345 87.775 186.515 ;
        RECT 88.065 186.345 88.235 186.515 ;
        RECT 88.525 186.345 88.695 186.515 ;
        RECT 88.985 186.345 89.155 186.515 ;
        RECT 89.445 186.345 89.615 186.515 ;
        RECT 89.905 186.345 90.075 186.515 ;
        RECT 90.365 186.345 90.535 186.515 ;
        RECT 90.825 186.345 90.995 186.515 ;
        RECT 91.285 186.345 91.455 186.515 ;
        RECT 91.745 186.345 91.915 186.515 ;
        RECT 92.205 186.345 92.375 186.515 ;
        RECT 92.665 186.345 92.835 186.515 ;
        RECT 93.125 186.345 93.295 186.515 ;
        RECT 93.585 186.345 93.755 186.515 ;
        RECT 94.045 186.345 94.215 186.515 ;
        RECT 94.505 186.345 94.675 186.515 ;
        RECT 94.965 186.345 95.135 186.515 ;
        RECT 95.425 186.345 95.595 186.515 ;
        RECT 95.885 186.345 96.055 186.515 ;
        RECT 96.345 186.345 96.515 186.515 ;
        RECT 96.805 186.345 96.975 186.515 ;
        RECT 97.265 186.345 97.435 186.515 ;
        RECT 97.725 186.345 97.895 186.515 ;
        RECT 98.185 186.345 98.355 186.515 ;
        RECT 98.645 186.345 98.815 186.515 ;
        RECT 99.105 186.345 99.275 186.515 ;
        RECT 99.565 186.345 99.735 186.515 ;
        RECT 100.025 186.345 100.195 186.515 ;
        RECT 100.485 186.345 100.655 186.515 ;
        RECT 100.945 186.345 101.115 186.515 ;
        RECT 101.405 186.345 101.575 186.515 ;
        RECT 101.865 186.345 102.035 186.515 ;
        RECT 102.325 186.345 102.495 186.515 ;
        RECT 102.785 186.345 102.955 186.515 ;
        RECT 103.245 186.345 103.415 186.515 ;
        RECT 103.705 186.345 103.875 186.515 ;
        RECT 104.165 186.345 104.335 186.515 ;
        RECT 104.625 186.345 104.795 186.515 ;
        RECT 105.085 186.345 105.255 186.515 ;
        RECT 105.545 186.345 105.715 186.515 ;
        RECT 106.005 186.345 106.175 186.515 ;
        RECT 106.465 186.345 106.635 186.515 ;
        RECT 106.925 186.345 107.095 186.515 ;
        RECT 107.385 186.345 107.555 186.515 ;
        RECT 107.845 186.345 108.015 186.515 ;
        RECT 108.305 186.345 108.475 186.515 ;
        RECT 108.765 186.345 108.935 186.515 ;
        RECT 109.225 186.345 109.395 186.515 ;
        RECT 109.685 186.345 109.855 186.515 ;
        RECT 110.145 186.345 110.315 186.515 ;
        RECT 110.605 186.345 110.775 186.515 ;
        RECT 111.065 186.345 111.235 186.515 ;
        RECT 111.525 186.345 111.695 186.515 ;
        RECT 111.985 186.345 112.155 186.515 ;
        RECT 112.445 186.345 112.615 186.515 ;
        RECT 112.905 186.345 113.075 186.515 ;
        RECT 113.365 186.345 113.535 186.515 ;
        RECT 113.825 186.345 113.995 186.515 ;
        RECT 114.285 186.345 114.455 186.515 ;
        RECT 114.745 186.345 114.915 186.515 ;
        RECT 115.205 186.345 115.375 186.515 ;
        RECT 115.665 186.345 115.835 186.515 ;
        RECT 116.125 186.345 116.295 186.515 ;
        RECT 116.585 186.345 116.755 186.515 ;
        RECT 117.045 186.345 117.215 186.515 ;
        RECT 117.505 186.345 117.675 186.515 ;
        RECT 117.965 186.345 118.135 186.515 ;
        RECT 118.425 186.345 118.595 186.515 ;
        RECT 118.885 186.345 119.055 186.515 ;
        RECT 119.345 186.345 119.515 186.515 ;
        RECT 119.805 186.345 119.975 186.515 ;
        RECT 120.265 186.345 120.435 186.515 ;
        RECT 120.725 186.345 120.895 186.515 ;
        RECT 121.185 186.345 121.355 186.515 ;
        RECT 121.645 186.345 121.815 186.515 ;
        RECT 67.825 183.625 67.995 183.795 ;
        RECT 68.285 183.625 68.455 183.795 ;
        RECT 68.745 183.625 68.915 183.795 ;
        RECT 69.205 183.625 69.375 183.795 ;
        RECT 69.665 183.625 69.835 183.795 ;
        RECT 70.125 183.625 70.295 183.795 ;
        RECT 70.585 183.625 70.755 183.795 ;
        RECT 71.045 183.625 71.215 183.795 ;
        RECT 71.505 183.625 71.675 183.795 ;
        RECT 71.965 183.625 72.135 183.795 ;
        RECT 72.425 183.625 72.595 183.795 ;
        RECT 72.885 183.625 73.055 183.795 ;
        RECT 73.345 183.625 73.515 183.795 ;
        RECT 73.805 183.625 73.975 183.795 ;
        RECT 74.265 183.625 74.435 183.795 ;
        RECT 74.725 183.625 74.895 183.795 ;
        RECT 75.185 183.625 75.355 183.795 ;
        RECT 75.645 183.625 75.815 183.795 ;
        RECT 76.105 183.625 76.275 183.795 ;
        RECT 76.565 183.625 76.735 183.795 ;
        RECT 77.025 183.625 77.195 183.795 ;
        RECT 77.485 183.625 77.655 183.795 ;
        RECT 77.945 183.625 78.115 183.795 ;
        RECT 78.405 183.625 78.575 183.795 ;
        RECT 78.865 183.625 79.035 183.795 ;
        RECT 79.325 183.625 79.495 183.795 ;
        RECT 79.785 183.625 79.955 183.795 ;
        RECT 80.245 183.625 80.415 183.795 ;
        RECT 80.705 183.625 80.875 183.795 ;
        RECT 81.165 183.625 81.335 183.795 ;
        RECT 81.625 183.625 81.795 183.795 ;
        RECT 82.085 183.625 82.255 183.795 ;
        RECT 82.545 183.625 82.715 183.795 ;
        RECT 83.005 183.625 83.175 183.795 ;
        RECT 83.465 183.625 83.635 183.795 ;
        RECT 83.925 183.625 84.095 183.795 ;
        RECT 84.385 183.625 84.555 183.795 ;
        RECT 84.845 183.625 85.015 183.795 ;
        RECT 85.305 183.625 85.475 183.795 ;
        RECT 85.765 183.625 85.935 183.795 ;
        RECT 86.225 183.625 86.395 183.795 ;
        RECT 86.685 183.625 86.855 183.795 ;
        RECT 87.145 183.625 87.315 183.795 ;
        RECT 87.605 183.625 87.775 183.795 ;
        RECT 88.065 183.625 88.235 183.795 ;
        RECT 88.525 183.625 88.695 183.795 ;
        RECT 88.985 183.625 89.155 183.795 ;
        RECT 89.445 183.625 89.615 183.795 ;
        RECT 89.905 183.625 90.075 183.795 ;
        RECT 90.365 183.625 90.535 183.795 ;
        RECT 90.825 183.625 90.995 183.795 ;
        RECT 91.285 183.625 91.455 183.795 ;
        RECT 91.745 183.625 91.915 183.795 ;
        RECT 92.205 183.625 92.375 183.795 ;
        RECT 92.665 183.625 92.835 183.795 ;
        RECT 93.125 183.625 93.295 183.795 ;
        RECT 93.585 183.625 93.755 183.795 ;
        RECT 94.045 183.625 94.215 183.795 ;
        RECT 94.505 183.625 94.675 183.795 ;
        RECT 94.965 183.625 95.135 183.795 ;
        RECT 95.425 183.625 95.595 183.795 ;
        RECT 95.885 183.625 96.055 183.795 ;
        RECT 96.345 183.625 96.515 183.795 ;
        RECT 96.805 183.625 96.975 183.795 ;
        RECT 97.265 183.625 97.435 183.795 ;
        RECT 97.725 183.625 97.895 183.795 ;
        RECT 98.185 183.625 98.355 183.795 ;
        RECT 98.645 183.625 98.815 183.795 ;
        RECT 99.105 183.625 99.275 183.795 ;
        RECT 99.565 183.625 99.735 183.795 ;
        RECT 100.025 183.625 100.195 183.795 ;
        RECT 100.485 183.625 100.655 183.795 ;
        RECT 100.945 183.625 101.115 183.795 ;
        RECT 101.405 183.625 101.575 183.795 ;
        RECT 101.865 183.625 102.035 183.795 ;
        RECT 102.325 183.625 102.495 183.795 ;
        RECT 102.785 183.625 102.955 183.795 ;
        RECT 103.245 183.625 103.415 183.795 ;
        RECT 103.705 183.625 103.875 183.795 ;
        RECT 104.165 183.625 104.335 183.795 ;
        RECT 104.625 183.625 104.795 183.795 ;
        RECT 105.085 183.625 105.255 183.795 ;
        RECT 105.545 183.625 105.715 183.795 ;
        RECT 106.005 183.625 106.175 183.795 ;
        RECT 106.465 183.625 106.635 183.795 ;
        RECT 106.925 183.625 107.095 183.795 ;
        RECT 107.385 183.625 107.555 183.795 ;
        RECT 107.845 183.625 108.015 183.795 ;
        RECT 108.305 183.625 108.475 183.795 ;
        RECT 108.765 183.625 108.935 183.795 ;
        RECT 109.225 183.625 109.395 183.795 ;
        RECT 109.685 183.625 109.855 183.795 ;
        RECT 110.145 183.625 110.315 183.795 ;
        RECT 110.605 183.625 110.775 183.795 ;
        RECT 111.065 183.625 111.235 183.795 ;
        RECT 111.525 183.625 111.695 183.795 ;
        RECT 111.985 183.625 112.155 183.795 ;
        RECT 112.445 183.625 112.615 183.795 ;
        RECT 112.905 183.625 113.075 183.795 ;
        RECT 113.365 183.625 113.535 183.795 ;
        RECT 113.825 183.625 113.995 183.795 ;
        RECT 114.285 183.625 114.455 183.795 ;
        RECT 114.745 183.625 114.915 183.795 ;
        RECT 115.205 183.625 115.375 183.795 ;
        RECT 115.665 183.625 115.835 183.795 ;
        RECT 116.125 183.625 116.295 183.795 ;
        RECT 116.585 183.625 116.755 183.795 ;
        RECT 117.045 183.625 117.215 183.795 ;
        RECT 117.505 183.625 117.675 183.795 ;
        RECT 117.965 183.625 118.135 183.795 ;
        RECT 118.425 183.625 118.595 183.795 ;
        RECT 118.885 183.625 119.055 183.795 ;
        RECT 119.345 183.625 119.515 183.795 ;
        RECT 119.805 183.625 119.975 183.795 ;
        RECT 120.265 183.625 120.435 183.795 ;
        RECT 120.725 183.625 120.895 183.795 ;
        RECT 121.185 183.625 121.355 183.795 ;
        RECT 121.645 183.625 121.815 183.795 ;
        RECT 67.825 180.905 67.995 181.075 ;
        RECT 68.285 180.905 68.455 181.075 ;
        RECT 68.745 180.905 68.915 181.075 ;
        RECT 69.205 180.905 69.375 181.075 ;
        RECT 69.665 180.905 69.835 181.075 ;
        RECT 70.125 180.905 70.295 181.075 ;
        RECT 70.585 180.905 70.755 181.075 ;
        RECT 71.045 180.905 71.215 181.075 ;
        RECT 71.505 180.905 71.675 181.075 ;
        RECT 71.965 180.905 72.135 181.075 ;
        RECT 72.425 180.905 72.595 181.075 ;
        RECT 72.885 180.905 73.055 181.075 ;
        RECT 73.345 180.905 73.515 181.075 ;
        RECT 73.805 180.905 73.975 181.075 ;
        RECT 74.265 180.905 74.435 181.075 ;
        RECT 74.725 180.905 74.895 181.075 ;
        RECT 75.185 180.905 75.355 181.075 ;
        RECT 75.645 180.905 75.815 181.075 ;
        RECT 76.105 180.905 76.275 181.075 ;
        RECT 76.565 180.905 76.735 181.075 ;
        RECT 77.025 180.905 77.195 181.075 ;
        RECT 77.485 180.905 77.655 181.075 ;
        RECT 77.945 180.905 78.115 181.075 ;
        RECT 78.405 180.905 78.575 181.075 ;
        RECT 78.865 180.905 79.035 181.075 ;
        RECT 79.325 180.905 79.495 181.075 ;
        RECT 79.785 180.905 79.955 181.075 ;
        RECT 80.245 180.905 80.415 181.075 ;
        RECT 80.705 180.905 80.875 181.075 ;
        RECT 81.165 180.905 81.335 181.075 ;
        RECT 81.625 180.905 81.795 181.075 ;
        RECT 82.085 180.905 82.255 181.075 ;
        RECT 82.545 180.905 82.715 181.075 ;
        RECT 83.005 180.905 83.175 181.075 ;
        RECT 83.465 180.905 83.635 181.075 ;
        RECT 83.925 180.905 84.095 181.075 ;
        RECT 84.385 180.905 84.555 181.075 ;
        RECT 84.845 180.905 85.015 181.075 ;
        RECT 85.305 180.905 85.475 181.075 ;
        RECT 85.765 180.905 85.935 181.075 ;
        RECT 86.225 180.905 86.395 181.075 ;
        RECT 86.685 180.905 86.855 181.075 ;
        RECT 87.145 180.905 87.315 181.075 ;
        RECT 87.605 180.905 87.775 181.075 ;
        RECT 88.065 180.905 88.235 181.075 ;
        RECT 88.525 180.905 88.695 181.075 ;
        RECT 88.985 180.905 89.155 181.075 ;
        RECT 89.445 180.905 89.615 181.075 ;
        RECT 89.905 180.905 90.075 181.075 ;
        RECT 90.365 180.905 90.535 181.075 ;
        RECT 90.825 180.905 90.995 181.075 ;
        RECT 91.285 180.905 91.455 181.075 ;
        RECT 91.745 180.905 91.915 181.075 ;
        RECT 92.205 180.905 92.375 181.075 ;
        RECT 92.665 180.905 92.835 181.075 ;
        RECT 93.125 180.905 93.295 181.075 ;
        RECT 93.585 180.905 93.755 181.075 ;
        RECT 94.045 180.905 94.215 181.075 ;
        RECT 94.505 180.905 94.675 181.075 ;
        RECT 94.965 180.905 95.135 181.075 ;
        RECT 95.425 180.905 95.595 181.075 ;
        RECT 95.885 180.905 96.055 181.075 ;
        RECT 96.345 180.905 96.515 181.075 ;
        RECT 96.805 180.905 96.975 181.075 ;
        RECT 97.265 180.905 97.435 181.075 ;
        RECT 97.725 180.905 97.895 181.075 ;
        RECT 98.185 180.905 98.355 181.075 ;
        RECT 98.645 180.905 98.815 181.075 ;
        RECT 99.105 180.905 99.275 181.075 ;
        RECT 99.565 180.905 99.735 181.075 ;
        RECT 100.025 180.905 100.195 181.075 ;
        RECT 100.485 180.905 100.655 181.075 ;
        RECT 100.945 180.905 101.115 181.075 ;
        RECT 101.405 180.905 101.575 181.075 ;
        RECT 101.865 180.905 102.035 181.075 ;
        RECT 102.325 180.905 102.495 181.075 ;
        RECT 102.785 180.905 102.955 181.075 ;
        RECT 103.245 180.905 103.415 181.075 ;
        RECT 103.705 180.905 103.875 181.075 ;
        RECT 104.165 180.905 104.335 181.075 ;
        RECT 104.625 180.905 104.795 181.075 ;
        RECT 105.085 180.905 105.255 181.075 ;
        RECT 105.545 180.905 105.715 181.075 ;
        RECT 106.005 180.905 106.175 181.075 ;
        RECT 106.465 180.905 106.635 181.075 ;
        RECT 106.925 180.905 107.095 181.075 ;
        RECT 107.385 180.905 107.555 181.075 ;
        RECT 107.845 180.905 108.015 181.075 ;
        RECT 108.305 180.905 108.475 181.075 ;
        RECT 108.765 180.905 108.935 181.075 ;
        RECT 109.225 180.905 109.395 181.075 ;
        RECT 109.685 180.905 109.855 181.075 ;
        RECT 110.145 180.905 110.315 181.075 ;
        RECT 110.605 180.905 110.775 181.075 ;
        RECT 111.065 180.905 111.235 181.075 ;
        RECT 111.525 180.905 111.695 181.075 ;
        RECT 111.985 180.905 112.155 181.075 ;
        RECT 112.445 180.905 112.615 181.075 ;
        RECT 112.905 180.905 113.075 181.075 ;
        RECT 113.365 180.905 113.535 181.075 ;
        RECT 113.825 180.905 113.995 181.075 ;
        RECT 114.285 180.905 114.455 181.075 ;
        RECT 114.745 180.905 114.915 181.075 ;
        RECT 115.205 180.905 115.375 181.075 ;
        RECT 115.665 180.905 115.835 181.075 ;
        RECT 116.125 180.905 116.295 181.075 ;
        RECT 116.585 180.905 116.755 181.075 ;
        RECT 117.045 180.905 117.215 181.075 ;
        RECT 117.505 180.905 117.675 181.075 ;
        RECT 117.965 180.905 118.135 181.075 ;
        RECT 118.425 180.905 118.595 181.075 ;
        RECT 118.885 180.905 119.055 181.075 ;
        RECT 119.345 180.905 119.515 181.075 ;
        RECT 119.805 180.905 119.975 181.075 ;
        RECT 120.265 180.905 120.435 181.075 ;
        RECT 120.725 180.905 120.895 181.075 ;
        RECT 121.185 180.905 121.355 181.075 ;
        RECT 121.645 180.905 121.815 181.075 ;
        RECT 67.825 178.185 67.995 178.355 ;
        RECT 68.285 178.185 68.455 178.355 ;
        RECT 68.745 178.185 68.915 178.355 ;
        RECT 69.205 178.185 69.375 178.355 ;
        RECT 69.665 178.185 69.835 178.355 ;
        RECT 70.125 178.185 70.295 178.355 ;
        RECT 70.585 178.185 70.755 178.355 ;
        RECT 71.045 178.185 71.215 178.355 ;
        RECT 71.505 178.185 71.675 178.355 ;
        RECT 71.965 178.185 72.135 178.355 ;
        RECT 72.425 178.185 72.595 178.355 ;
        RECT 72.885 178.185 73.055 178.355 ;
        RECT 73.345 178.185 73.515 178.355 ;
        RECT 73.805 178.185 73.975 178.355 ;
        RECT 74.265 178.185 74.435 178.355 ;
        RECT 74.725 178.185 74.895 178.355 ;
        RECT 75.185 178.185 75.355 178.355 ;
        RECT 75.645 178.185 75.815 178.355 ;
        RECT 76.105 178.185 76.275 178.355 ;
        RECT 76.565 178.185 76.735 178.355 ;
        RECT 77.025 178.185 77.195 178.355 ;
        RECT 77.485 178.185 77.655 178.355 ;
        RECT 77.945 178.185 78.115 178.355 ;
        RECT 78.405 178.185 78.575 178.355 ;
        RECT 78.865 178.185 79.035 178.355 ;
        RECT 79.325 178.185 79.495 178.355 ;
        RECT 79.785 178.185 79.955 178.355 ;
        RECT 80.245 178.185 80.415 178.355 ;
        RECT 80.705 178.185 80.875 178.355 ;
        RECT 81.165 178.185 81.335 178.355 ;
        RECT 81.625 178.185 81.795 178.355 ;
        RECT 82.085 178.185 82.255 178.355 ;
        RECT 82.545 178.185 82.715 178.355 ;
        RECT 83.005 178.185 83.175 178.355 ;
        RECT 83.465 178.185 83.635 178.355 ;
        RECT 83.925 178.185 84.095 178.355 ;
        RECT 84.385 178.185 84.555 178.355 ;
        RECT 84.845 178.185 85.015 178.355 ;
        RECT 85.305 178.185 85.475 178.355 ;
        RECT 85.765 178.185 85.935 178.355 ;
        RECT 86.225 178.185 86.395 178.355 ;
        RECT 86.685 178.185 86.855 178.355 ;
        RECT 87.145 178.185 87.315 178.355 ;
        RECT 87.605 178.185 87.775 178.355 ;
        RECT 88.065 178.185 88.235 178.355 ;
        RECT 88.525 178.185 88.695 178.355 ;
        RECT 88.985 178.185 89.155 178.355 ;
        RECT 89.445 178.185 89.615 178.355 ;
        RECT 89.905 178.185 90.075 178.355 ;
        RECT 90.365 178.185 90.535 178.355 ;
        RECT 90.825 178.185 90.995 178.355 ;
        RECT 91.285 178.185 91.455 178.355 ;
        RECT 91.745 178.185 91.915 178.355 ;
        RECT 92.205 178.185 92.375 178.355 ;
        RECT 92.665 178.185 92.835 178.355 ;
        RECT 93.125 178.185 93.295 178.355 ;
        RECT 93.585 178.185 93.755 178.355 ;
        RECT 94.045 178.185 94.215 178.355 ;
        RECT 94.505 178.185 94.675 178.355 ;
        RECT 94.965 178.185 95.135 178.355 ;
        RECT 95.425 178.185 95.595 178.355 ;
        RECT 95.885 178.185 96.055 178.355 ;
        RECT 96.345 178.185 96.515 178.355 ;
        RECT 96.805 178.185 96.975 178.355 ;
        RECT 97.265 178.185 97.435 178.355 ;
        RECT 97.725 178.185 97.895 178.355 ;
        RECT 98.185 178.185 98.355 178.355 ;
        RECT 98.645 178.185 98.815 178.355 ;
        RECT 99.105 178.185 99.275 178.355 ;
        RECT 99.565 178.185 99.735 178.355 ;
        RECT 100.025 178.185 100.195 178.355 ;
        RECT 100.485 178.185 100.655 178.355 ;
        RECT 100.945 178.185 101.115 178.355 ;
        RECT 101.405 178.185 101.575 178.355 ;
        RECT 101.865 178.185 102.035 178.355 ;
        RECT 102.325 178.185 102.495 178.355 ;
        RECT 102.785 178.185 102.955 178.355 ;
        RECT 103.245 178.185 103.415 178.355 ;
        RECT 103.705 178.185 103.875 178.355 ;
        RECT 104.165 178.185 104.335 178.355 ;
        RECT 104.625 178.185 104.795 178.355 ;
        RECT 105.085 178.185 105.255 178.355 ;
        RECT 105.545 178.185 105.715 178.355 ;
        RECT 106.005 178.185 106.175 178.355 ;
        RECT 106.465 178.185 106.635 178.355 ;
        RECT 106.925 178.185 107.095 178.355 ;
        RECT 107.385 178.185 107.555 178.355 ;
        RECT 107.845 178.185 108.015 178.355 ;
        RECT 108.305 178.185 108.475 178.355 ;
        RECT 108.765 178.185 108.935 178.355 ;
        RECT 109.225 178.185 109.395 178.355 ;
        RECT 109.685 178.185 109.855 178.355 ;
        RECT 110.145 178.185 110.315 178.355 ;
        RECT 110.605 178.185 110.775 178.355 ;
        RECT 111.065 178.185 111.235 178.355 ;
        RECT 111.525 178.185 111.695 178.355 ;
        RECT 111.985 178.185 112.155 178.355 ;
        RECT 112.445 178.185 112.615 178.355 ;
        RECT 112.905 178.185 113.075 178.355 ;
        RECT 113.365 178.185 113.535 178.355 ;
        RECT 113.825 178.185 113.995 178.355 ;
        RECT 114.285 178.185 114.455 178.355 ;
        RECT 114.745 178.185 114.915 178.355 ;
        RECT 115.205 178.185 115.375 178.355 ;
        RECT 115.665 178.185 115.835 178.355 ;
        RECT 116.125 178.185 116.295 178.355 ;
        RECT 116.585 178.185 116.755 178.355 ;
        RECT 117.045 178.185 117.215 178.355 ;
        RECT 117.505 178.185 117.675 178.355 ;
        RECT 117.965 178.185 118.135 178.355 ;
        RECT 118.425 178.185 118.595 178.355 ;
        RECT 118.885 178.185 119.055 178.355 ;
        RECT 119.345 178.185 119.515 178.355 ;
        RECT 119.805 178.185 119.975 178.355 ;
        RECT 120.265 178.185 120.435 178.355 ;
        RECT 120.725 178.185 120.895 178.355 ;
        RECT 121.185 178.185 121.355 178.355 ;
        RECT 121.645 178.185 121.815 178.355 ;
        RECT 67.825 175.465 67.995 175.635 ;
        RECT 68.285 175.465 68.455 175.635 ;
        RECT 68.745 175.465 68.915 175.635 ;
        RECT 69.205 175.465 69.375 175.635 ;
        RECT 69.665 175.465 69.835 175.635 ;
        RECT 70.125 175.465 70.295 175.635 ;
        RECT 70.585 175.465 70.755 175.635 ;
        RECT 71.045 175.465 71.215 175.635 ;
        RECT 71.505 175.465 71.675 175.635 ;
        RECT 71.965 175.465 72.135 175.635 ;
        RECT 72.425 175.465 72.595 175.635 ;
        RECT 72.885 175.465 73.055 175.635 ;
        RECT 73.345 175.465 73.515 175.635 ;
        RECT 73.805 175.465 73.975 175.635 ;
        RECT 74.265 175.465 74.435 175.635 ;
        RECT 74.725 175.465 74.895 175.635 ;
        RECT 75.185 175.465 75.355 175.635 ;
        RECT 75.645 175.465 75.815 175.635 ;
        RECT 76.105 175.465 76.275 175.635 ;
        RECT 76.565 175.465 76.735 175.635 ;
        RECT 77.025 175.465 77.195 175.635 ;
        RECT 77.485 175.465 77.655 175.635 ;
        RECT 77.945 175.465 78.115 175.635 ;
        RECT 78.405 175.465 78.575 175.635 ;
        RECT 78.865 175.465 79.035 175.635 ;
        RECT 79.325 175.465 79.495 175.635 ;
        RECT 79.785 175.465 79.955 175.635 ;
        RECT 80.245 175.465 80.415 175.635 ;
        RECT 80.705 175.465 80.875 175.635 ;
        RECT 81.165 175.465 81.335 175.635 ;
        RECT 81.625 175.465 81.795 175.635 ;
        RECT 82.085 175.465 82.255 175.635 ;
        RECT 82.545 175.465 82.715 175.635 ;
        RECT 83.005 175.465 83.175 175.635 ;
        RECT 83.465 175.465 83.635 175.635 ;
        RECT 83.925 175.465 84.095 175.635 ;
        RECT 84.385 175.465 84.555 175.635 ;
        RECT 84.845 175.465 85.015 175.635 ;
        RECT 85.305 175.465 85.475 175.635 ;
        RECT 85.765 175.465 85.935 175.635 ;
        RECT 86.225 175.465 86.395 175.635 ;
        RECT 86.685 175.465 86.855 175.635 ;
        RECT 87.145 175.465 87.315 175.635 ;
        RECT 87.605 175.465 87.775 175.635 ;
        RECT 88.065 175.465 88.235 175.635 ;
        RECT 88.525 175.465 88.695 175.635 ;
        RECT 88.985 175.465 89.155 175.635 ;
        RECT 89.445 175.465 89.615 175.635 ;
        RECT 89.905 175.465 90.075 175.635 ;
        RECT 90.365 175.465 90.535 175.635 ;
        RECT 90.825 175.465 90.995 175.635 ;
        RECT 91.285 175.465 91.455 175.635 ;
        RECT 91.745 175.465 91.915 175.635 ;
        RECT 92.205 175.465 92.375 175.635 ;
        RECT 92.665 175.465 92.835 175.635 ;
        RECT 93.125 175.465 93.295 175.635 ;
        RECT 93.585 175.465 93.755 175.635 ;
        RECT 94.045 175.465 94.215 175.635 ;
        RECT 94.505 175.465 94.675 175.635 ;
        RECT 94.965 175.465 95.135 175.635 ;
        RECT 95.425 175.465 95.595 175.635 ;
        RECT 95.885 175.465 96.055 175.635 ;
        RECT 96.345 175.465 96.515 175.635 ;
        RECT 96.805 175.465 96.975 175.635 ;
        RECT 97.265 175.465 97.435 175.635 ;
        RECT 97.725 175.465 97.895 175.635 ;
        RECT 98.185 175.465 98.355 175.635 ;
        RECT 98.645 175.465 98.815 175.635 ;
        RECT 99.105 175.465 99.275 175.635 ;
        RECT 99.565 175.465 99.735 175.635 ;
        RECT 100.025 175.465 100.195 175.635 ;
        RECT 100.485 175.465 100.655 175.635 ;
        RECT 100.945 175.465 101.115 175.635 ;
        RECT 101.405 175.465 101.575 175.635 ;
        RECT 101.865 175.465 102.035 175.635 ;
        RECT 102.325 175.465 102.495 175.635 ;
        RECT 102.785 175.465 102.955 175.635 ;
        RECT 103.245 175.465 103.415 175.635 ;
        RECT 103.705 175.465 103.875 175.635 ;
        RECT 104.165 175.465 104.335 175.635 ;
        RECT 104.625 175.465 104.795 175.635 ;
        RECT 105.085 175.465 105.255 175.635 ;
        RECT 105.545 175.465 105.715 175.635 ;
        RECT 106.005 175.465 106.175 175.635 ;
        RECT 106.465 175.465 106.635 175.635 ;
        RECT 106.925 175.465 107.095 175.635 ;
        RECT 107.385 175.465 107.555 175.635 ;
        RECT 107.845 175.465 108.015 175.635 ;
        RECT 108.305 175.465 108.475 175.635 ;
        RECT 108.765 175.465 108.935 175.635 ;
        RECT 109.225 175.465 109.395 175.635 ;
        RECT 109.685 175.465 109.855 175.635 ;
        RECT 110.145 175.465 110.315 175.635 ;
        RECT 110.605 175.465 110.775 175.635 ;
        RECT 111.065 175.465 111.235 175.635 ;
        RECT 111.525 175.465 111.695 175.635 ;
        RECT 111.985 175.465 112.155 175.635 ;
        RECT 112.445 175.465 112.615 175.635 ;
        RECT 112.905 175.465 113.075 175.635 ;
        RECT 113.365 175.465 113.535 175.635 ;
        RECT 113.825 175.465 113.995 175.635 ;
        RECT 114.285 175.465 114.455 175.635 ;
        RECT 114.745 175.465 114.915 175.635 ;
        RECT 115.205 175.465 115.375 175.635 ;
        RECT 115.665 175.465 115.835 175.635 ;
        RECT 116.125 175.465 116.295 175.635 ;
        RECT 116.585 175.465 116.755 175.635 ;
        RECT 117.045 175.465 117.215 175.635 ;
        RECT 117.505 175.465 117.675 175.635 ;
        RECT 117.965 175.465 118.135 175.635 ;
        RECT 118.425 175.465 118.595 175.635 ;
        RECT 118.885 175.465 119.055 175.635 ;
        RECT 119.345 175.465 119.515 175.635 ;
        RECT 119.805 175.465 119.975 175.635 ;
        RECT 120.265 175.465 120.435 175.635 ;
        RECT 120.725 175.465 120.895 175.635 ;
        RECT 121.185 175.465 121.355 175.635 ;
        RECT 121.645 175.465 121.815 175.635 ;
        RECT 99.105 174.955 99.275 175.125 ;
        RECT 95.425 173.255 95.595 173.425 ;
        RECT 96.345 173.935 96.515 174.105 ;
        RECT 96.805 174.275 96.975 174.445 ;
        RECT 97.265 173.935 97.435 174.105 ;
        RECT 97.725 174.275 97.895 174.445 ;
        RECT 102.760 174.615 102.930 174.785 ;
        RECT 102.760 173.595 102.930 173.765 ;
        RECT 104.600 174.615 104.770 174.785 ;
        RECT 104.140 173.595 104.310 173.765 ;
        RECT 106.000 174.615 106.170 174.785 ;
        RECT 105.545 173.935 105.715 174.105 ;
        RECT 106.925 173.935 107.095 174.105 ;
        RECT 106.460 173.595 106.630 173.765 ;
        RECT 118.885 174.275 119.055 174.445 ;
        RECT 117.965 173.255 118.135 173.425 ;
        RECT 67.825 172.745 67.995 172.915 ;
        RECT 68.285 172.745 68.455 172.915 ;
        RECT 68.745 172.745 68.915 172.915 ;
        RECT 69.205 172.745 69.375 172.915 ;
        RECT 69.665 172.745 69.835 172.915 ;
        RECT 70.125 172.745 70.295 172.915 ;
        RECT 70.585 172.745 70.755 172.915 ;
        RECT 71.045 172.745 71.215 172.915 ;
        RECT 71.505 172.745 71.675 172.915 ;
        RECT 71.965 172.745 72.135 172.915 ;
        RECT 72.425 172.745 72.595 172.915 ;
        RECT 72.885 172.745 73.055 172.915 ;
        RECT 73.345 172.745 73.515 172.915 ;
        RECT 73.805 172.745 73.975 172.915 ;
        RECT 74.265 172.745 74.435 172.915 ;
        RECT 74.725 172.745 74.895 172.915 ;
        RECT 75.185 172.745 75.355 172.915 ;
        RECT 75.645 172.745 75.815 172.915 ;
        RECT 76.105 172.745 76.275 172.915 ;
        RECT 76.565 172.745 76.735 172.915 ;
        RECT 77.025 172.745 77.195 172.915 ;
        RECT 77.485 172.745 77.655 172.915 ;
        RECT 77.945 172.745 78.115 172.915 ;
        RECT 78.405 172.745 78.575 172.915 ;
        RECT 78.865 172.745 79.035 172.915 ;
        RECT 79.325 172.745 79.495 172.915 ;
        RECT 79.785 172.745 79.955 172.915 ;
        RECT 80.245 172.745 80.415 172.915 ;
        RECT 80.705 172.745 80.875 172.915 ;
        RECT 81.165 172.745 81.335 172.915 ;
        RECT 81.625 172.745 81.795 172.915 ;
        RECT 82.085 172.745 82.255 172.915 ;
        RECT 82.545 172.745 82.715 172.915 ;
        RECT 83.005 172.745 83.175 172.915 ;
        RECT 83.465 172.745 83.635 172.915 ;
        RECT 83.925 172.745 84.095 172.915 ;
        RECT 84.385 172.745 84.555 172.915 ;
        RECT 84.845 172.745 85.015 172.915 ;
        RECT 85.305 172.745 85.475 172.915 ;
        RECT 85.765 172.745 85.935 172.915 ;
        RECT 86.225 172.745 86.395 172.915 ;
        RECT 86.685 172.745 86.855 172.915 ;
        RECT 87.145 172.745 87.315 172.915 ;
        RECT 87.605 172.745 87.775 172.915 ;
        RECT 88.065 172.745 88.235 172.915 ;
        RECT 88.525 172.745 88.695 172.915 ;
        RECT 88.985 172.745 89.155 172.915 ;
        RECT 89.445 172.745 89.615 172.915 ;
        RECT 89.905 172.745 90.075 172.915 ;
        RECT 90.365 172.745 90.535 172.915 ;
        RECT 90.825 172.745 90.995 172.915 ;
        RECT 91.285 172.745 91.455 172.915 ;
        RECT 91.745 172.745 91.915 172.915 ;
        RECT 92.205 172.745 92.375 172.915 ;
        RECT 92.665 172.745 92.835 172.915 ;
        RECT 93.125 172.745 93.295 172.915 ;
        RECT 93.585 172.745 93.755 172.915 ;
        RECT 94.045 172.745 94.215 172.915 ;
        RECT 94.505 172.745 94.675 172.915 ;
        RECT 94.965 172.745 95.135 172.915 ;
        RECT 95.425 172.745 95.595 172.915 ;
        RECT 95.885 172.745 96.055 172.915 ;
        RECT 96.345 172.745 96.515 172.915 ;
        RECT 96.805 172.745 96.975 172.915 ;
        RECT 97.265 172.745 97.435 172.915 ;
        RECT 97.725 172.745 97.895 172.915 ;
        RECT 98.185 172.745 98.355 172.915 ;
        RECT 98.645 172.745 98.815 172.915 ;
        RECT 99.105 172.745 99.275 172.915 ;
        RECT 99.565 172.745 99.735 172.915 ;
        RECT 100.025 172.745 100.195 172.915 ;
        RECT 100.485 172.745 100.655 172.915 ;
        RECT 100.945 172.745 101.115 172.915 ;
        RECT 101.405 172.745 101.575 172.915 ;
        RECT 101.865 172.745 102.035 172.915 ;
        RECT 102.325 172.745 102.495 172.915 ;
        RECT 102.785 172.745 102.955 172.915 ;
        RECT 103.245 172.745 103.415 172.915 ;
        RECT 103.705 172.745 103.875 172.915 ;
        RECT 104.165 172.745 104.335 172.915 ;
        RECT 104.625 172.745 104.795 172.915 ;
        RECT 105.085 172.745 105.255 172.915 ;
        RECT 105.545 172.745 105.715 172.915 ;
        RECT 106.005 172.745 106.175 172.915 ;
        RECT 106.465 172.745 106.635 172.915 ;
        RECT 106.925 172.745 107.095 172.915 ;
        RECT 107.385 172.745 107.555 172.915 ;
        RECT 107.845 172.745 108.015 172.915 ;
        RECT 108.305 172.745 108.475 172.915 ;
        RECT 108.765 172.745 108.935 172.915 ;
        RECT 109.225 172.745 109.395 172.915 ;
        RECT 109.685 172.745 109.855 172.915 ;
        RECT 110.145 172.745 110.315 172.915 ;
        RECT 110.605 172.745 110.775 172.915 ;
        RECT 111.065 172.745 111.235 172.915 ;
        RECT 111.525 172.745 111.695 172.915 ;
        RECT 111.985 172.745 112.155 172.915 ;
        RECT 112.445 172.745 112.615 172.915 ;
        RECT 112.905 172.745 113.075 172.915 ;
        RECT 113.365 172.745 113.535 172.915 ;
        RECT 113.825 172.745 113.995 172.915 ;
        RECT 114.285 172.745 114.455 172.915 ;
        RECT 114.745 172.745 114.915 172.915 ;
        RECT 115.205 172.745 115.375 172.915 ;
        RECT 115.665 172.745 115.835 172.915 ;
        RECT 116.125 172.745 116.295 172.915 ;
        RECT 116.585 172.745 116.755 172.915 ;
        RECT 117.045 172.745 117.215 172.915 ;
        RECT 117.505 172.745 117.675 172.915 ;
        RECT 117.965 172.745 118.135 172.915 ;
        RECT 118.425 172.745 118.595 172.915 ;
        RECT 118.885 172.745 119.055 172.915 ;
        RECT 119.345 172.745 119.515 172.915 ;
        RECT 119.805 172.745 119.975 172.915 ;
        RECT 120.265 172.745 120.435 172.915 ;
        RECT 120.725 172.745 120.895 172.915 ;
        RECT 121.185 172.745 121.355 172.915 ;
        RECT 121.645 172.745 121.815 172.915 ;
        RECT 85.770 171.895 85.940 172.065 ;
        RECT 85.305 171.215 85.475 171.385 ;
        RECT 86.685 171.215 86.855 171.385 ;
        RECT 86.230 170.875 86.400 171.045 ;
        RECT 88.090 171.895 88.260 172.065 ;
        RECT 87.630 170.875 87.800 171.045 ;
        RECT 89.470 171.895 89.640 172.065 ;
        RECT 89.470 170.875 89.640 171.045 ;
        RECT 104.165 172.235 104.335 172.405 ;
        RECT 94.045 171.215 94.215 171.385 ;
        RECT 93.125 170.535 93.295 170.705 ;
        RECT 103.245 171.215 103.415 171.385 ;
        RECT 100.485 170.535 100.655 170.705 ;
        RECT 105.545 170.535 105.715 170.705 ;
        RECT 110.145 171.215 110.315 171.385 ;
        RECT 109.685 170.535 109.855 170.705 ;
        RECT 67.825 170.025 67.995 170.195 ;
        RECT 68.285 170.025 68.455 170.195 ;
        RECT 68.745 170.025 68.915 170.195 ;
        RECT 69.205 170.025 69.375 170.195 ;
        RECT 69.665 170.025 69.835 170.195 ;
        RECT 70.125 170.025 70.295 170.195 ;
        RECT 70.585 170.025 70.755 170.195 ;
        RECT 71.045 170.025 71.215 170.195 ;
        RECT 71.505 170.025 71.675 170.195 ;
        RECT 71.965 170.025 72.135 170.195 ;
        RECT 72.425 170.025 72.595 170.195 ;
        RECT 72.885 170.025 73.055 170.195 ;
        RECT 73.345 170.025 73.515 170.195 ;
        RECT 73.805 170.025 73.975 170.195 ;
        RECT 74.265 170.025 74.435 170.195 ;
        RECT 74.725 170.025 74.895 170.195 ;
        RECT 75.185 170.025 75.355 170.195 ;
        RECT 75.645 170.025 75.815 170.195 ;
        RECT 76.105 170.025 76.275 170.195 ;
        RECT 76.565 170.025 76.735 170.195 ;
        RECT 77.025 170.025 77.195 170.195 ;
        RECT 77.485 170.025 77.655 170.195 ;
        RECT 77.945 170.025 78.115 170.195 ;
        RECT 78.405 170.025 78.575 170.195 ;
        RECT 78.865 170.025 79.035 170.195 ;
        RECT 79.325 170.025 79.495 170.195 ;
        RECT 79.785 170.025 79.955 170.195 ;
        RECT 80.245 170.025 80.415 170.195 ;
        RECT 80.705 170.025 80.875 170.195 ;
        RECT 81.165 170.025 81.335 170.195 ;
        RECT 81.625 170.025 81.795 170.195 ;
        RECT 82.085 170.025 82.255 170.195 ;
        RECT 82.545 170.025 82.715 170.195 ;
        RECT 83.005 170.025 83.175 170.195 ;
        RECT 83.465 170.025 83.635 170.195 ;
        RECT 83.925 170.025 84.095 170.195 ;
        RECT 84.385 170.025 84.555 170.195 ;
        RECT 84.845 170.025 85.015 170.195 ;
        RECT 85.305 170.025 85.475 170.195 ;
        RECT 85.765 170.025 85.935 170.195 ;
        RECT 86.225 170.025 86.395 170.195 ;
        RECT 86.685 170.025 86.855 170.195 ;
        RECT 87.145 170.025 87.315 170.195 ;
        RECT 87.605 170.025 87.775 170.195 ;
        RECT 88.065 170.025 88.235 170.195 ;
        RECT 88.525 170.025 88.695 170.195 ;
        RECT 88.985 170.025 89.155 170.195 ;
        RECT 89.445 170.025 89.615 170.195 ;
        RECT 89.905 170.025 90.075 170.195 ;
        RECT 90.365 170.025 90.535 170.195 ;
        RECT 90.825 170.025 90.995 170.195 ;
        RECT 91.285 170.025 91.455 170.195 ;
        RECT 91.745 170.025 91.915 170.195 ;
        RECT 92.205 170.025 92.375 170.195 ;
        RECT 92.665 170.025 92.835 170.195 ;
        RECT 93.125 170.025 93.295 170.195 ;
        RECT 93.585 170.025 93.755 170.195 ;
        RECT 94.045 170.025 94.215 170.195 ;
        RECT 94.505 170.025 94.675 170.195 ;
        RECT 94.965 170.025 95.135 170.195 ;
        RECT 95.425 170.025 95.595 170.195 ;
        RECT 95.885 170.025 96.055 170.195 ;
        RECT 96.345 170.025 96.515 170.195 ;
        RECT 96.805 170.025 96.975 170.195 ;
        RECT 97.265 170.025 97.435 170.195 ;
        RECT 97.725 170.025 97.895 170.195 ;
        RECT 98.185 170.025 98.355 170.195 ;
        RECT 98.645 170.025 98.815 170.195 ;
        RECT 99.105 170.025 99.275 170.195 ;
        RECT 99.565 170.025 99.735 170.195 ;
        RECT 100.025 170.025 100.195 170.195 ;
        RECT 100.485 170.025 100.655 170.195 ;
        RECT 100.945 170.025 101.115 170.195 ;
        RECT 101.405 170.025 101.575 170.195 ;
        RECT 101.865 170.025 102.035 170.195 ;
        RECT 102.325 170.025 102.495 170.195 ;
        RECT 102.785 170.025 102.955 170.195 ;
        RECT 103.245 170.025 103.415 170.195 ;
        RECT 103.705 170.025 103.875 170.195 ;
        RECT 104.165 170.025 104.335 170.195 ;
        RECT 104.625 170.025 104.795 170.195 ;
        RECT 105.085 170.025 105.255 170.195 ;
        RECT 105.545 170.025 105.715 170.195 ;
        RECT 106.005 170.025 106.175 170.195 ;
        RECT 106.465 170.025 106.635 170.195 ;
        RECT 106.925 170.025 107.095 170.195 ;
        RECT 107.385 170.025 107.555 170.195 ;
        RECT 107.845 170.025 108.015 170.195 ;
        RECT 108.305 170.025 108.475 170.195 ;
        RECT 108.765 170.025 108.935 170.195 ;
        RECT 109.225 170.025 109.395 170.195 ;
        RECT 109.685 170.025 109.855 170.195 ;
        RECT 110.145 170.025 110.315 170.195 ;
        RECT 110.605 170.025 110.775 170.195 ;
        RECT 111.065 170.025 111.235 170.195 ;
        RECT 111.525 170.025 111.695 170.195 ;
        RECT 111.985 170.025 112.155 170.195 ;
        RECT 112.445 170.025 112.615 170.195 ;
        RECT 112.905 170.025 113.075 170.195 ;
        RECT 113.365 170.025 113.535 170.195 ;
        RECT 113.825 170.025 113.995 170.195 ;
        RECT 114.285 170.025 114.455 170.195 ;
        RECT 114.745 170.025 114.915 170.195 ;
        RECT 115.205 170.025 115.375 170.195 ;
        RECT 115.665 170.025 115.835 170.195 ;
        RECT 116.125 170.025 116.295 170.195 ;
        RECT 116.585 170.025 116.755 170.195 ;
        RECT 117.045 170.025 117.215 170.195 ;
        RECT 117.505 170.025 117.675 170.195 ;
        RECT 117.965 170.025 118.135 170.195 ;
        RECT 118.425 170.025 118.595 170.195 ;
        RECT 118.885 170.025 119.055 170.195 ;
        RECT 119.345 170.025 119.515 170.195 ;
        RECT 119.805 170.025 119.975 170.195 ;
        RECT 120.265 170.025 120.435 170.195 ;
        RECT 120.725 170.025 120.895 170.195 ;
        RECT 121.185 170.025 121.355 170.195 ;
        RECT 121.645 170.025 121.815 170.195 ;
        RECT 83.925 168.495 84.095 168.665 ;
        RECT 84.385 168.835 84.555 169.005 ;
        RECT 84.845 168.495 85.015 168.665 ;
        RECT 85.305 168.835 85.475 169.005 ;
        RECT 86.685 168.495 86.855 168.665 ;
        RECT 86.225 167.815 86.395 167.985 ;
        RECT 88.525 169.515 88.695 169.685 ;
        RECT 89.445 168.155 89.615 168.325 ;
        RECT 88.525 167.815 88.695 167.985 ;
        RECT 89.905 168.835 90.075 169.005 ;
        RECT 92.665 168.835 92.835 169.005 ;
        RECT 94.505 167.815 94.675 167.985 ;
        RECT 98.645 169.515 98.815 169.685 ;
        RECT 100.485 169.515 100.655 169.685 ;
        RECT 98.185 168.835 98.355 169.005 ;
        RECT 99.200 168.835 99.370 169.005 ;
        RECT 100.025 168.495 100.195 168.665 ;
        RECT 101.965 169.175 102.135 169.345 ;
        RECT 102.265 168.860 102.435 169.030 ;
        RECT 98.645 168.155 98.815 168.325 ;
        RECT 103.345 168.835 103.515 169.005 ;
        RECT 105.205 169.175 105.375 169.345 ;
        RECT 105.565 169.175 105.735 169.345 ;
        RECT 103.345 168.155 103.515 168.325 ;
        RECT 106.925 168.835 107.095 169.005 ;
        RECT 106.465 168.155 106.635 168.325 ;
        RECT 107.845 169.175 108.015 169.345 ;
        RECT 108.355 168.155 108.525 168.325 ;
        RECT 108.760 168.835 108.930 169.005 ;
        RECT 109.225 168.495 109.395 168.665 ;
        RECT 67.825 167.305 67.995 167.475 ;
        RECT 68.285 167.305 68.455 167.475 ;
        RECT 68.745 167.305 68.915 167.475 ;
        RECT 69.205 167.305 69.375 167.475 ;
        RECT 69.665 167.305 69.835 167.475 ;
        RECT 70.125 167.305 70.295 167.475 ;
        RECT 70.585 167.305 70.755 167.475 ;
        RECT 71.045 167.305 71.215 167.475 ;
        RECT 71.505 167.305 71.675 167.475 ;
        RECT 71.965 167.305 72.135 167.475 ;
        RECT 72.425 167.305 72.595 167.475 ;
        RECT 72.885 167.305 73.055 167.475 ;
        RECT 73.345 167.305 73.515 167.475 ;
        RECT 73.805 167.305 73.975 167.475 ;
        RECT 74.265 167.305 74.435 167.475 ;
        RECT 74.725 167.305 74.895 167.475 ;
        RECT 75.185 167.305 75.355 167.475 ;
        RECT 75.645 167.305 75.815 167.475 ;
        RECT 76.105 167.305 76.275 167.475 ;
        RECT 76.565 167.305 76.735 167.475 ;
        RECT 77.025 167.305 77.195 167.475 ;
        RECT 77.485 167.305 77.655 167.475 ;
        RECT 77.945 167.305 78.115 167.475 ;
        RECT 78.405 167.305 78.575 167.475 ;
        RECT 78.865 167.305 79.035 167.475 ;
        RECT 79.325 167.305 79.495 167.475 ;
        RECT 79.785 167.305 79.955 167.475 ;
        RECT 80.245 167.305 80.415 167.475 ;
        RECT 80.705 167.305 80.875 167.475 ;
        RECT 81.165 167.305 81.335 167.475 ;
        RECT 81.625 167.305 81.795 167.475 ;
        RECT 82.085 167.305 82.255 167.475 ;
        RECT 82.545 167.305 82.715 167.475 ;
        RECT 83.005 167.305 83.175 167.475 ;
        RECT 83.465 167.305 83.635 167.475 ;
        RECT 83.925 167.305 84.095 167.475 ;
        RECT 84.385 167.305 84.555 167.475 ;
        RECT 84.845 167.305 85.015 167.475 ;
        RECT 85.305 167.305 85.475 167.475 ;
        RECT 85.765 167.305 85.935 167.475 ;
        RECT 86.225 167.305 86.395 167.475 ;
        RECT 86.685 167.305 86.855 167.475 ;
        RECT 87.145 167.305 87.315 167.475 ;
        RECT 87.605 167.305 87.775 167.475 ;
        RECT 88.065 167.305 88.235 167.475 ;
        RECT 88.525 167.305 88.695 167.475 ;
        RECT 88.985 167.305 89.155 167.475 ;
        RECT 89.445 167.305 89.615 167.475 ;
        RECT 89.905 167.305 90.075 167.475 ;
        RECT 90.365 167.305 90.535 167.475 ;
        RECT 90.825 167.305 90.995 167.475 ;
        RECT 91.285 167.305 91.455 167.475 ;
        RECT 91.745 167.305 91.915 167.475 ;
        RECT 92.205 167.305 92.375 167.475 ;
        RECT 92.665 167.305 92.835 167.475 ;
        RECT 93.125 167.305 93.295 167.475 ;
        RECT 93.585 167.305 93.755 167.475 ;
        RECT 94.045 167.305 94.215 167.475 ;
        RECT 94.505 167.305 94.675 167.475 ;
        RECT 94.965 167.305 95.135 167.475 ;
        RECT 95.425 167.305 95.595 167.475 ;
        RECT 95.885 167.305 96.055 167.475 ;
        RECT 96.345 167.305 96.515 167.475 ;
        RECT 96.805 167.305 96.975 167.475 ;
        RECT 97.265 167.305 97.435 167.475 ;
        RECT 97.725 167.305 97.895 167.475 ;
        RECT 98.185 167.305 98.355 167.475 ;
        RECT 98.645 167.305 98.815 167.475 ;
        RECT 99.105 167.305 99.275 167.475 ;
        RECT 99.565 167.305 99.735 167.475 ;
        RECT 100.025 167.305 100.195 167.475 ;
        RECT 100.485 167.305 100.655 167.475 ;
        RECT 100.945 167.305 101.115 167.475 ;
        RECT 101.405 167.305 101.575 167.475 ;
        RECT 101.865 167.305 102.035 167.475 ;
        RECT 102.325 167.305 102.495 167.475 ;
        RECT 102.785 167.305 102.955 167.475 ;
        RECT 103.245 167.305 103.415 167.475 ;
        RECT 103.705 167.305 103.875 167.475 ;
        RECT 104.165 167.305 104.335 167.475 ;
        RECT 104.625 167.305 104.795 167.475 ;
        RECT 105.085 167.305 105.255 167.475 ;
        RECT 105.545 167.305 105.715 167.475 ;
        RECT 106.005 167.305 106.175 167.475 ;
        RECT 106.465 167.305 106.635 167.475 ;
        RECT 106.925 167.305 107.095 167.475 ;
        RECT 107.385 167.305 107.555 167.475 ;
        RECT 107.845 167.305 108.015 167.475 ;
        RECT 108.305 167.305 108.475 167.475 ;
        RECT 108.765 167.305 108.935 167.475 ;
        RECT 109.225 167.305 109.395 167.475 ;
        RECT 109.685 167.305 109.855 167.475 ;
        RECT 110.145 167.305 110.315 167.475 ;
        RECT 110.605 167.305 110.775 167.475 ;
        RECT 111.065 167.305 111.235 167.475 ;
        RECT 111.525 167.305 111.695 167.475 ;
        RECT 111.985 167.305 112.155 167.475 ;
        RECT 112.445 167.305 112.615 167.475 ;
        RECT 112.905 167.305 113.075 167.475 ;
        RECT 113.365 167.305 113.535 167.475 ;
        RECT 113.825 167.305 113.995 167.475 ;
        RECT 114.285 167.305 114.455 167.475 ;
        RECT 114.745 167.305 114.915 167.475 ;
        RECT 115.205 167.305 115.375 167.475 ;
        RECT 115.665 167.305 115.835 167.475 ;
        RECT 116.125 167.305 116.295 167.475 ;
        RECT 116.585 167.305 116.755 167.475 ;
        RECT 117.045 167.305 117.215 167.475 ;
        RECT 117.505 167.305 117.675 167.475 ;
        RECT 117.965 167.305 118.135 167.475 ;
        RECT 118.425 167.305 118.595 167.475 ;
        RECT 118.885 167.305 119.055 167.475 ;
        RECT 119.345 167.305 119.515 167.475 ;
        RECT 119.805 167.305 119.975 167.475 ;
        RECT 120.265 167.305 120.435 167.475 ;
        RECT 120.725 167.305 120.895 167.475 ;
        RECT 121.185 167.305 121.355 167.475 ;
        RECT 121.645 167.305 121.815 167.475 ;
        RECT 86.685 166.455 86.855 166.625 ;
        RECT 85.305 165.775 85.475 165.945 ;
        RECT 87.605 166.115 87.775 166.285 ;
        RECT 88.990 166.455 89.160 166.625 ;
        RECT 85.765 165.095 85.935 165.265 ;
        RECT 87.145 165.775 87.315 165.945 ;
        RECT 86.685 165.435 86.855 165.605 ;
        RECT 88.525 166.115 88.695 166.285 ;
        RECT 88.065 165.775 88.235 165.945 ;
        RECT 89.905 165.775 90.075 165.945 ;
        RECT 89.450 165.435 89.620 165.605 ;
        RECT 91.310 166.455 91.480 166.625 ;
        RECT 90.850 165.435 91.020 165.605 ;
        RECT 92.690 166.455 92.860 166.625 ;
        RECT 92.690 165.435 92.860 165.605 ;
        RECT 95.425 165.095 95.595 165.265 ;
        RECT 102.325 165.775 102.495 165.945 ;
        RECT 101.405 165.095 101.575 165.265 ;
        RECT 67.825 164.585 67.995 164.755 ;
        RECT 68.285 164.585 68.455 164.755 ;
        RECT 68.745 164.585 68.915 164.755 ;
        RECT 69.205 164.585 69.375 164.755 ;
        RECT 69.665 164.585 69.835 164.755 ;
        RECT 70.125 164.585 70.295 164.755 ;
        RECT 70.585 164.585 70.755 164.755 ;
        RECT 71.045 164.585 71.215 164.755 ;
        RECT 71.505 164.585 71.675 164.755 ;
        RECT 71.965 164.585 72.135 164.755 ;
        RECT 72.425 164.585 72.595 164.755 ;
        RECT 72.885 164.585 73.055 164.755 ;
        RECT 73.345 164.585 73.515 164.755 ;
        RECT 73.805 164.585 73.975 164.755 ;
        RECT 74.265 164.585 74.435 164.755 ;
        RECT 74.725 164.585 74.895 164.755 ;
        RECT 75.185 164.585 75.355 164.755 ;
        RECT 75.645 164.585 75.815 164.755 ;
        RECT 76.105 164.585 76.275 164.755 ;
        RECT 76.565 164.585 76.735 164.755 ;
        RECT 77.025 164.585 77.195 164.755 ;
        RECT 77.485 164.585 77.655 164.755 ;
        RECT 77.945 164.585 78.115 164.755 ;
        RECT 78.405 164.585 78.575 164.755 ;
        RECT 78.865 164.585 79.035 164.755 ;
        RECT 79.325 164.585 79.495 164.755 ;
        RECT 79.785 164.585 79.955 164.755 ;
        RECT 80.245 164.585 80.415 164.755 ;
        RECT 80.705 164.585 80.875 164.755 ;
        RECT 81.165 164.585 81.335 164.755 ;
        RECT 81.625 164.585 81.795 164.755 ;
        RECT 82.085 164.585 82.255 164.755 ;
        RECT 82.545 164.585 82.715 164.755 ;
        RECT 83.005 164.585 83.175 164.755 ;
        RECT 83.465 164.585 83.635 164.755 ;
        RECT 83.925 164.585 84.095 164.755 ;
        RECT 84.385 164.585 84.555 164.755 ;
        RECT 84.845 164.585 85.015 164.755 ;
        RECT 85.305 164.585 85.475 164.755 ;
        RECT 85.765 164.585 85.935 164.755 ;
        RECT 86.225 164.585 86.395 164.755 ;
        RECT 86.685 164.585 86.855 164.755 ;
        RECT 87.145 164.585 87.315 164.755 ;
        RECT 87.605 164.585 87.775 164.755 ;
        RECT 88.065 164.585 88.235 164.755 ;
        RECT 88.525 164.585 88.695 164.755 ;
        RECT 88.985 164.585 89.155 164.755 ;
        RECT 89.445 164.585 89.615 164.755 ;
        RECT 89.905 164.585 90.075 164.755 ;
        RECT 90.365 164.585 90.535 164.755 ;
        RECT 90.825 164.585 90.995 164.755 ;
        RECT 91.285 164.585 91.455 164.755 ;
        RECT 91.745 164.585 91.915 164.755 ;
        RECT 92.205 164.585 92.375 164.755 ;
        RECT 92.665 164.585 92.835 164.755 ;
        RECT 93.125 164.585 93.295 164.755 ;
        RECT 93.585 164.585 93.755 164.755 ;
        RECT 94.045 164.585 94.215 164.755 ;
        RECT 94.505 164.585 94.675 164.755 ;
        RECT 94.965 164.585 95.135 164.755 ;
        RECT 95.425 164.585 95.595 164.755 ;
        RECT 95.885 164.585 96.055 164.755 ;
        RECT 96.345 164.585 96.515 164.755 ;
        RECT 96.805 164.585 96.975 164.755 ;
        RECT 97.265 164.585 97.435 164.755 ;
        RECT 97.725 164.585 97.895 164.755 ;
        RECT 98.185 164.585 98.355 164.755 ;
        RECT 98.645 164.585 98.815 164.755 ;
        RECT 99.105 164.585 99.275 164.755 ;
        RECT 99.565 164.585 99.735 164.755 ;
        RECT 100.025 164.585 100.195 164.755 ;
        RECT 100.485 164.585 100.655 164.755 ;
        RECT 100.945 164.585 101.115 164.755 ;
        RECT 101.405 164.585 101.575 164.755 ;
        RECT 101.865 164.585 102.035 164.755 ;
        RECT 102.325 164.585 102.495 164.755 ;
        RECT 102.785 164.585 102.955 164.755 ;
        RECT 103.245 164.585 103.415 164.755 ;
        RECT 103.705 164.585 103.875 164.755 ;
        RECT 104.165 164.585 104.335 164.755 ;
        RECT 104.625 164.585 104.795 164.755 ;
        RECT 105.085 164.585 105.255 164.755 ;
        RECT 105.545 164.585 105.715 164.755 ;
        RECT 106.005 164.585 106.175 164.755 ;
        RECT 106.465 164.585 106.635 164.755 ;
        RECT 106.925 164.585 107.095 164.755 ;
        RECT 107.385 164.585 107.555 164.755 ;
        RECT 107.845 164.585 108.015 164.755 ;
        RECT 108.305 164.585 108.475 164.755 ;
        RECT 108.765 164.585 108.935 164.755 ;
        RECT 109.225 164.585 109.395 164.755 ;
        RECT 109.685 164.585 109.855 164.755 ;
        RECT 110.145 164.585 110.315 164.755 ;
        RECT 110.605 164.585 110.775 164.755 ;
        RECT 111.065 164.585 111.235 164.755 ;
        RECT 111.525 164.585 111.695 164.755 ;
        RECT 111.985 164.585 112.155 164.755 ;
        RECT 112.445 164.585 112.615 164.755 ;
        RECT 112.905 164.585 113.075 164.755 ;
        RECT 113.365 164.585 113.535 164.755 ;
        RECT 113.825 164.585 113.995 164.755 ;
        RECT 114.285 164.585 114.455 164.755 ;
        RECT 114.745 164.585 114.915 164.755 ;
        RECT 115.205 164.585 115.375 164.755 ;
        RECT 115.665 164.585 115.835 164.755 ;
        RECT 116.125 164.585 116.295 164.755 ;
        RECT 116.585 164.585 116.755 164.755 ;
        RECT 117.045 164.585 117.215 164.755 ;
        RECT 117.505 164.585 117.675 164.755 ;
        RECT 117.965 164.585 118.135 164.755 ;
        RECT 118.425 164.585 118.595 164.755 ;
        RECT 118.885 164.585 119.055 164.755 ;
        RECT 119.345 164.585 119.515 164.755 ;
        RECT 119.805 164.585 119.975 164.755 ;
        RECT 120.265 164.585 120.435 164.755 ;
        RECT 120.725 164.585 120.895 164.755 ;
        RECT 121.185 164.585 121.355 164.755 ;
        RECT 121.645 164.585 121.815 164.755 ;
        RECT 90.825 164.075 90.995 164.245 ;
        RECT 94.045 163.735 94.215 163.905 ;
        RECT 91.745 163.395 91.915 163.565 ;
        RECT 92.665 163.055 92.835 163.225 ;
        RECT 94.965 163.395 95.135 163.565 ;
        RECT 95.425 163.395 95.595 163.565 ;
        RECT 94.045 162.715 94.215 162.885 ;
        RECT 97.725 162.375 97.895 162.545 ;
        RECT 100.460 163.735 100.630 163.905 ;
        RECT 100.460 162.715 100.630 162.885 ;
        RECT 102.300 163.735 102.470 163.905 ;
        RECT 101.840 162.715 102.010 162.885 ;
        RECT 103.700 163.735 103.870 163.905 ;
        RECT 103.245 163.055 103.415 163.225 ;
        RECT 104.625 163.055 104.795 163.225 ;
        RECT 104.160 162.715 104.330 162.885 ;
        RECT 67.825 161.865 67.995 162.035 ;
        RECT 68.285 161.865 68.455 162.035 ;
        RECT 68.745 161.865 68.915 162.035 ;
        RECT 69.205 161.865 69.375 162.035 ;
        RECT 69.665 161.865 69.835 162.035 ;
        RECT 70.125 161.865 70.295 162.035 ;
        RECT 70.585 161.865 70.755 162.035 ;
        RECT 71.045 161.865 71.215 162.035 ;
        RECT 71.505 161.865 71.675 162.035 ;
        RECT 71.965 161.865 72.135 162.035 ;
        RECT 72.425 161.865 72.595 162.035 ;
        RECT 72.885 161.865 73.055 162.035 ;
        RECT 73.345 161.865 73.515 162.035 ;
        RECT 73.805 161.865 73.975 162.035 ;
        RECT 74.265 161.865 74.435 162.035 ;
        RECT 74.725 161.865 74.895 162.035 ;
        RECT 75.185 161.865 75.355 162.035 ;
        RECT 75.645 161.865 75.815 162.035 ;
        RECT 76.105 161.865 76.275 162.035 ;
        RECT 76.565 161.865 76.735 162.035 ;
        RECT 77.025 161.865 77.195 162.035 ;
        RECT 77.485 161.865 77.655 162.035 ;
        RECT 77.945 161.865 78.115 162.035 ;
        RECT 78.405 161.865 78.575 162.035 ;
        RECT 78.865 161.865 79.035 162.035 ;
        RECT 79.325 161.865 79.495 162.035 ;
        RECT 79.785 161.865 79.955 162.035 ;
        RECT 80.245 161.865 80.415 162.035 ;
        RECT 80.705 161.865 80.875 162.035 ;
        RECT 81.165 161.865 81.335 162.035 ;
        RECT 81.625 161.865 81.795 162.035 ;
        RECT 82.085 161.865 82.255 162.035 ;
        RECT 82.545 161.865 82.715 162.035 ;
        RECT 83.005 161.865 83.175 162.035 ;
        RECT 83.465 161.865 83.635 162.035 ;
        RECT 83.925 161.865 84.095 162.035 ;
        RECT 84.385 161.865 84.555 162.035 ;
        RECT 84.845 161.865 85.015 162.035 ;
        RECT 85.305 161.865 85.475 162.035 ;
        RECT 85.765 161.865 85.935 162.035 ;
        RECT 86.225 161.865 86.395 162.035 ;
        RECT 86.685 161.865 86.855 162.035 ;
        RECT 87.145 161.865 87.315 162.035 ;
        RECT 87.605 161.865 87.775 162.035 ;
        RECT 88.065 161.865 88.235 162.035 ;
        RECT 88.525 161.865 88.695 162.035 ;
        RECT 88.985 161.865 89.155 162.035 ;
        RECT 89.445 161.865 89.615 162.035 ;
        RECT 89.905 161.865 90.075 162.035 ;
        RECT 90.365 161.865 90.535 162.035 ;
        RECT 90.825 161.865 90.995 162.035 ;
        RECT 91.285 161.865 91.455 162.035 ;
        RECT 91.745 161.865 91.915 162.035 ;
        RECT 92.205 161.865 92.375 162.035 ;
        RECT 92.665 161.865 92.835 162.035 ;
        RECT 93.125 161.865 93.295 162.035 ;
        RECT 93.585 161.865 93.755 162.035 ;
        RECT 94.045 161.865 94.215 162.035 ;
        RECT 94.505 161.865 94.675 162.035 ;
        RECT 94.965 161.865 95.135 162.035 ;
        RECT 95.425 161.865 95.595 162.035 ;
        RECT 95.885 161.865 96.055 162.035 ;
        RECT 96.345 161.865 96.515 162.035 ;
        RECT 96.805 161.865 96.975 162.035 ;
        RECT 97.265 161.865 97.435 162.035 ;
        RECT 97.725 161.865 97.895 162.035 ;
        RECT 98.185 161.865 98.355 162.035 ;
        RECT 98.645 161.865 98.815 162.035 ;
        RECT 99.105 161.865 99.275 162.035 ;
        RECT 99.565 161.865 99.735 162.035 ;
        RECT 100.025 161.865 100.195 162.035 ;
        RECT 100.485 161.865 100.655 162.035 ;
        RECT 100.945 161.865 101.115 162.035 ;
        RECT 101.405 161.865 101.575 162.035 ;
        RECT 101.865 161.865 102.035 162.035 ;
        RECT 102.325 161.865 102.495 162.035 ;
        RECT 102.785 161.865 102.955 162.035 ;
        RECT 103.245 161.865 103.415 162.035 ;
        RECT 103.705 161.865 103.875 162.035 ;
        RECT 104.165 161.865 104.335 162.035 ;
        RECT 104.625 161.865 104.795 162.035 ;
        RECT 105.085 161.865 105.255 162.035 ;
        RECT 105.545 161.865 105.715 162.035 ;
        RECT 106.005 161.865 106.175 162.035 ;
        RECT 106.465 161.865 106.635 162.035 ;
        RECT 106.925 161.865 107.095 162.035 ;
        RECT 107.385 161.865 107.555 162.035 ;
        RECT 107.845 161.865 108.015 162.035 ;
        RECT 108.305 161.865 108.475 162.035 ;
        RECT 108.765 161.865 108.935 162.035 ;
        RECT 109.225 161.865 109.395 162.035 ;
        RECT 109.685 161.865 109.855 162.035 ;
        RECT 110.145 161.865 110.315 162.035 ;
        RECT 110.605 161.865 110.775 162.035 ;
        RECT 111.065 161.865 111.235 162.035 ;
        RECT 111.525 161.865 111.695 162.035 ;
        RECT 111.985 161.865 112.155 162.035 ;
        RECT 112.445 161.865 112.615 162.035 ;
        RECT 112.905 161.865 113.075 162.035 ;
        RECT 113.365 161.865 113.535 162.035 ;
        RECT 113.825 161.865 113.995 162.035 ;
        RECT 114.285 161.865 114.455 162.035 ;
        RECT 114.745 161.865 114.915 162.035 ;
        RECT 115.205 161.865 115.375 162.035 ;
        RECT 115.665 161.865 115.835 162.035 ;
        RECT 116.125 161.865 116.295 162.035 ;
        RECT 116.585 161.865 116.755 162.035 ;
        RECT 117.045 161.865 117.215 162.035 ;
        RECT 117.505 161.865 117.675 162.035 ;
        RECT 117.965 161.865 118.135 162.035 ;
        RECT 118.425 161.865 118.595 162.035 ;
        RECT 118.885 161.865 119.055 162.035 ;
        RECT 119.345 161.865 119.515 162.035 ;
        RECT 119.805 161.865 119.975 162.035 ;
        RECT 120.265 161.865 120.435 162.035 ;
        RECT 120.725 161.865 120.895 162.035 ;
        RECT 121.185 161.865 121.355 162.035 ;
        RECT 121.645 161.865 121.815 162.035 ;
        RECT 83.465 161.355 83.635 161.525 ;
        RECT 89.905 159.995 90.075 160.165 ;
        RECT 98.185 160.675 98.355 160.845 ;
        RECT 100.945 161.355 101.115 161.525 ;
        RECT 101.865 160.675 102.035 160.845 ;
        RECT 101.405 160.335 101.575 160.505 ;
        RECT 102.325 160.335 102.495 160.505 ;
        RECT 113.365 161.355 113.535 161.525 ;
        RECT 106.925 159.995 107.095 160.165 ;
        RECT 67.825 159.145 67.995 159.315 ;
        RECT 68.285 159.145 68.455 159.315 ;
        RECT 68.745 159.145 68.915 159.315 ;
        RECT 69.205 159.145 69.375 159.315 ;
        RECT 69.665 159.145 69.835 159.315 ;
        RECT 70.125 159.145 70.295 159.315 ;
        RECT 70.585 159.145 70.755 159.315 ;
        RECT 71.045 159.145 71.215 159.315 ;
        RECT 71.505 159.145 71.675 159.315 ;
        RECT 71.965 159.145 72.135 159.315 ;
        RECT 72.425 159.145 72.595 159.315 ;
        RECT 72.885 159.145 73.055 159.315 ;
        RECT 73.345 159.145 73.515 159.315 ;
        RECT 73.805 159.145 73.975 159.315 ;
        RECT 74.265 159.145 74.435 159.315 ;
        RECT 74.725 159.145 74.895 159.315 ;
        RECT 75.185 159.145 75.355 159.315 ;
        RECT 75.645 159.145 75.815 159.315 ;
        RECT 76.105 159.145 76.275 159.315 ;
        RECT 76.565 159.145 76.735 159.315 ;
        RECT 77.025 159.145 77.195 159.315 ;
        RECT 77.485 159.145 77.655 159.315 ;
        RECT 77.945 159.145 78.115 159.315 ;
        RECT 78.405 159.145 78.575 159.315 ;
        RECT 78.865 159.145 79.035 159.315 ;
        RECT 79.325 159.145 79.495 159.315 ;
        RECT 79.785 159.145 79.955 159.315 ;
        RECT 80.245 159.145 80.415 159.315 ;
        RECT 80.705 159.145 80.875 159.315 ;
        RECT 81.165 159.145 81.335 159.315 ;
        RECT 81.625 159.145 81.795 159.315 ;
        RECT 82.085 159.145 82.255 159.315 ;
        RECT 82.545 159.145 82.715 159.315 ;
        RECT 83.005 159.145 83.175 159.315 ;
        RECT 83.465 159.145 83.635 159.315 ;
        RECT 83.925 159.145 84.095 159.315 ;
        RECT 84.385 159.145 84.555 159.315 ;
        RECT 84.845 159.145 85.015 159.315 ;
        RECT 85.305 159.145 85.475 159.315 ;
        RECT 85.765 159.145 85.935 159.315 ;
        RECT 86.225 159.145 86.395 159.315 ;
        RECT 86.685 159.145 86.855 159.315 ;
        RECT 87.145 159.145 87.315 159.315 ;
        RECT 87.605 159.145 87.775 159.315 ;
        RECT 88.065 159.145 88.235 159.315 ;
        RECT 88.525 159.145 88.695 159.315 ;
        RECT 88.985 159.145 89.155 159.315 ;
        RECT 89.445 159.145 89.615 159.315 ;
        RECT 89.905 159.145 90.075 159.315 ;
        RECT 90.365 159.145 90.535 159.315 ;
        RECT 90.825 159.145 90.995 159.315 ;
        RECT 91.285 159.145 91.455 159.315 ;
        RECT 91.745 159.145 91.915 159.315 ;
        RECT 92.205 159.145 92.375 159.315 ;
        RECT 92.665 159.145 92.835 159.315 ;
        RECT 93.125 159.145 93.295 159.315 ;
        RECT 93.585 159.145 93.755 159.315 ;
        RECT 94.045 159.145 94.215 159.315 ;
        RECT 94.505 159.145 94.675 159.315 ;
        RECT 94.965 159.145 95.135 159.315 ;
        RECT 95.425 159.145 95.595 159.315 ;
        RECT 95.885 159.145 96.055 159.315 ;
        RECT 96.345 159.145 96.515 159.315 ;
        RECT 96.805 159.145 96.975 159.315 ;
        RECT 97.265 159.145 97.435 159.315 ;
        RECT 97.725 159.145 97.895 159.315 ;
        RECT 98.185 159.145 98.355 159.315 ;
        RECT 98.645 159.145 98.815 159.315 ;
        RECT 99.105 159.145 99.275 159.315 ;
        RECT 99.565 159.145 99.735 159.315 ;
        RECT 100.025 159.145 100.195 159.315 ;
        RECT 100.485 159.145 100.655 159.315 ;
        RECT 100.945 159.145 101.115 159.315 ;
        RECT 101.405 159.145 101.575 159.315 ;
        RECT 101.865 159.145 102.035 159.315 ;
        RECT 102.325 159.145 102.495 159.315 ;
        RECT 102.785 159.145 102.955 159.315 ;
        RECT 103.245 159.145 103.415 159.315 ;
        RECT 103.705 159.145 103.875 159.315 ;
        RECT 104.165 159.145 104.335 159.315 ;
        RECT 104.625 159.145 104.795 159.315 ;
        RECT 105.085 159.145 105.255 159.315 ;
        RECT 105.545 159.145 105.715 159.315 ;
        RECT 106.005 159.145 106.175 159.315 ;
        RECT 106.465 159.145 106.635 159.315 ;
        RECT 106.925 159.145 107.095 159.315 ;
        RECT 107.385 159.145 107.555 159.315 ;
        RECT 107.845 159.145 108.015 159.315 ;
        RECT 108.305 159.145 108.475 159.315 ;
        RECT 108.765 159.145 108.935 159.315 ;
        RECT 109.225 159.145 109.395 159.315 ;
        RECT 109.685 159.145 109.855 159.315 ;
        RECT 110.145 159.145 110.315 159.315 ;
        RECT 110.605 159.145 110.775 159.315 ;
        RECT 111.065 159.145 111.235 159.315 ;
        RECT 111.525 159.145 111.695 159.315 ;
        RECT 111.985 159.145 112.155 159.315 ;
        RECT 112.445 159.145 112.615 159.315 ;
        RECT 112.905 159.145 113.075 159.315 ;
        RECT 113.365 159.145 113.535 159.315 ;
        RECT 113.825 159.145 113.995 159.315 ;
        RECT 114.285 159.145 114.455 159.315 ;
        RECT 114.745 159.145 114.915 159.315 ;
        RECT 115.205 159.145 115.375 159.315 ;
        RECT 115.665 159.145 115.835 159.315 ;
        RECT 116.125 159.145 116.295 159.315 ;
        RECT 116.585 159.145 116.755 159.315 ;
        RECT 117.045 159.145 117.215 159.315 ;
        RECT 117.505 159.145 117.675 159.315 ;
        RECT 117.965 159.145 118.135 159.315 ;
        RECT 118.425 159.145 118.595 159.315 ;
        RECT 118.885 159.145 119.055 159.315 ;
        RECT 119.345 159.145 119.515 159.315 ;
        RECT 119.805 159.145 119.975 159.315 ;
        RECT 120.265 159.145 120.435 159.315 ;
        RECT 120.725 159.145 120.895 159.315 ;
        RECT 121.185 159.145 121.355 159.315 ;
        RECT 121.645 159.145 121.815 159.315 ;
        RECT 86.630 74.280 86.800 76.265 ;
        RECT 88.720 74.240 88.890 76.225 ;
        RECT 90.840 74.090 91.010 76.075 ;
        RECT 93.110 74.090 93.280 76.075 ;
        RECT 95.480 74.340 95.650 76.325 ;
        RECT 90.840 60.410 91.010 62.395 ;
        RECT 93.210 60.560 93.380 62.545 ;
        RECT 95.580 60.310 95.750 62.295 ;
      LAYER met1 ;
        RECT 67.680 213.390 122.760 213.870 ;
        RECT 67.680 210.670 121.960 211.150 ;
        RECT 67.680 207.950 122.760 208.430 ;
        RECT 67.680 205.230 121.960 205.710 ;
        RECT 67.680 202.510 122.760 202.990 ;
        RECT 67.680 199.790 121.960 200.270 ;
        RECT 67.680 197.070 122.760 197.550 ;
        RECT 67.680 194.350 121.960 194.830 ;
        RECT 78.790 194.150 79.110 194.210 ;
        RECT 92.590 194.150 92.910 194.210 ;
        RECT 78.790 194.010 92.910 194.150 ;
        RECT 78.790 193.950 79.110 194.010 ;
        RECT 92.590 193.950 92.910 194.010 ;
        RECT 67.680 191.630 122.760 192.110 ;
        RECT 67.680 188.910 121.960 189.390 ;
        RECT 67.680 186.190 122.760 186.670 ;
        RECT 67.680 183.470 121.960 183.950 ;
        RECT 67.680 180.750 122.760 181.230 ;
        RECT 67.680 178.030 121.960 178.510 ;
        RECT 99.030 177.150 99.350 177.210 ;
        RECT 122.950 177.150 123.270 177.210 ;
        RECT 99.030 177.010 123.270 177.150 ;
        RECT 99.030 176.950 99.350 177.010 ;
        RECT 122.950 176.950 123.270 177.010 ;
        RECT 67.680 175.310 122.760 175.790 ;
        RECT 99.030 174.910 99.350 175.170 ;
        RECT 96.270 174.570 96.590 174.830 ;
        RECT 96.360 174.430 96.500 174.570 ;
        RECT 96.745 174.430 97.035 174.475 ;
        RECT 96.360 174.290 97.035 174.430 ;
        RECT 96.745 174.245 97.035 174.290 ;
        RECT 97.665 174.430 97.955 174.475 ;
        RECT 99.120 174.430 99.260 174.910 ;
        RECT 102.700 174.770 102.990 174.815 ;
        RECT 104.540 174.770 104.830 174.815 ;
        RECT 105.940 174.770 106.230 174.815 ;
        RECT 102.700 174.630 106.230 174.770 ;
        RECT 102.700 174.585 102.990 174.630 ;
        RECT 104.540 174.585 104.830 174.630 ;
        RECT 105.940 174.585 106.230 174.630 ;
        RECT 97.665 174.290 99.260 174.430 ;
        RECT 97.665 174.245 97.955 174.290 ;
        RECT 118.825 174.245 119.115 174.475 ;
        RECT 93.510 174.090 93.830 174.150 ;
        RECT 96.285 174.090 96.575 174.135 ;
        RECT 93.510 173.950 96.575 174.090 ;
        RECT 93.510 173.890 93.830 173.950 ;
        RECT 96.285 173.905 96.575 173.950 ;
        RECT 97.205 173.905 97.495 174.135 ;
        RECT 97.280 173.750 97.420 173.905 ;
        RECT 105.470 173.890 105.790 174.150 ;
        RECT 106.865 174.090 107.155 174.135 ;
        RECT 109.610 174.090 109.930 174.150 ;
        RECT 106.865 173.950 109.930 174.090 ;
        RECT 118.900 174.090 119.040 174.245 ;
        RECT 121.110 174.090 121.430 174.150 ;
        RECT 118.900 173.950 121.430 174.090 ;
        RECT 106.865 173.905 107.155 173.950 ;
        RECT 109.610 173.890 109.930 173.950 ;
        RECT 121.110 173.890 121.430 173.950 ;
        RECT 96.820 173.610 97.420 173.750 ;
        RECT 102.700 173.750 102.990 173.795 ;
        RECT 104.080 173.750 104.370 173.795 ;
        RECT 106.400 173.750 106.690 173.795 ;
        RECT 102.700 173.610 106.690 173.750 ;
        RECT 96.820 173.470 96.960 173.610 ;
        RECT 102.700 173.565 102.990 173.610 ;
        RECT 104.080 173.565 104.370 173.610 ;
        RECT 106.400 173.565 106.690 173.610 ;
        RECT 93.050 173.410 93.370 173.470 ;
        RECT 95.365 173.410 95.655 173.455 ;
        RECT 93.050 173.270 95.655 173.410 ;
        RECT 93.050 173.210 93.370 173.270 ;
        RECT 95.365 173.225 95.655 173.270 ;
        RECT 96.730 173.210 97.050 173.470 ;
        RECT 117.890 173.210 118.210 173.470 ;
        RECT 67.680 172.590 121.960 173.070 ;
        RECT 104.105 172.390 104.395 172.435 ;
        RECT 105.470 172.390 105.790 172.450 ;
        RECT 104.105 172.250 105.790 172.390 ;
        RECT 104.105 172.205 104.395 172.250 ;
        RECT 105.470 172.190 105.790 172.250 ;
        RECT 117.890 172.190 118.210 172.450 ;
        RECT 85.710 172.050 86.000 172.095 ;
        RECT 88.030 172.050 88.320 172.095 ;
        RECT 89.410 172.050 89.700 172.095 ;
        RECT 85.710 171.910 89.700 172.050 ;
        RECT 85.710 171.865 86.000 171.910 ;
        RECT 88.030 171.865 88.320 171.910 ;
        RECT 89.410 171.865 89.700 171.910 ;
        RECT 85.245 171.370 85.535 171.415 ;
        RECT 83.480 171.230 85.535 171.370 ;
        RECT 83.480 170.750 83.620 171.230 ;
        RECT 85.245 171.185 85.535 171.230 ;
        RECT 86.610 171.170 86.930 171.430 ;
        RECT 92.590 171.370 92.910 171.430 ;
        RECT 93.985 171.370 94.275 171.415 ;
        RECT 92.590 171.230 94.275 171.370 ;
        RECT 92.590 171.170 92.910 171.230 ;
        RECT 93.985 171.185 94.275 171.230 ;
        RECT 95.810 171.370 96.130 171.430 ;
        RECT 103.185 171.370 103.475 171.415 ;
        RECT 95.810 171.230 103.475 171.370 ;
        RECT 95.810 171.170 96.130 171.230 ;
        RECT 103.185 171.185 103.475 171.230 ;
        RECT 110.085 171.370 110.375 171.415 ;
        RECT 117.980 171.370 118.120 172.190 ;
        RECT 110.085 171.230 118.120 171.370 ;
        RECT 110.085 171.185 110.375 171.230 ;
        RECT 86.170 171.030 86.460 171.075 ;
        RECT 87.570 171.030 87.860 171.075 ;
        RECT 89.410 171.030 89.700 171.075 ;
        RECT 86.170 170.890 89.700 171.030 ;
        RECT 86.170 170.845 86.460 170.890 ;
        RECT 87.570 170.845 87.860 170.890 ;
        RECT 89.410 170.845 89.700 170.890 ;
        RECT 83.390 170.490 83.710 170.750 ;
        RECT 92.590 170.690 92.910 170.750 ;
        RECT 93.065 170.690 93.355 170.735 ;
        RECT 93.510 170.690 93.830 170.750 ;
        RECT 98.570 170.690 98.890 170.750 ;
        RECT 92.590 170.550 98.890 170.690 ;
        RECT 92.590 170.490 92.910 170.550 ;
        RECT 93.065 170.505 93.355 170.550 ;
        RECT 93.510 170.490 93.830 170.550 ;
        RECT 98.570 170.490 98.890 170.550 ;
        RECT 100.410 170.490 100.730 170.750 ;
        RECT 105.485 170.690 105.775 170.735 ;
        RECT 106.390 170.690 106.710 170.750 ;
        RECT 105.485 170.550 106.710 170.690 ;
        RECT 105.485 170.505 105.775 170.550 ;
        RECT 106.390 170.490 106.710 170.550 ;
        RECT 106.850 170.690 107.170 170.750 ;
        RECT 109.625 170.690 109.915 170.735 ;
        RECT 106.850 170.550 109.915 170.690 ;
        RECT 106.850 170.490 107.170 170.550 ;
        RECT 109.625 170.505 109.915 170.550 ;
        RECT 67.680 169.870 122.760 170.350 ;
        RECT 88.465 169.670 88.755 169.715 ;
        RECT 93.050 169.670 93.370 169.730 ;
        RECT 88.465 169.530 93.370 169.670 ;
        RECT 88.465 169.485 88.755 169.530 ;
        RECT 93.050 169.470 93.370 169.530 ;
        RECT 98.570 169.470 98.890 169.730 ;
        RECT 100.425 169.485 100.715 169.715 ;
        RECT 106.850 169.670 107.170 169.730 ;
        RECT 106.020 169.530 107.170 169.670 ;
        RECT 99.950 169.330 100.270 169.390 ;
        RECT 100.500 169.330 100.640 169.485 ;
        RECT 84.400 169.190 85.920 169.330 ;
        RECT 84.400 169.035 84.540 169.190 ;
        RECT 84.325 168.805 84.615 169.035 ;
        RECT 85.230 168.790 85.550 169.050 ;
        RECT 83.850 168.450 84.170 168.710 ;
        RECT 84.785 168.650 85.075 168.695 ;
        RECT 84.785 168.510 85.460 168.650 ;
        RECT 84.785 168.465 85.075 168.510 ;
        RECT 85.320 168.030 85.460 168.510 ;
        RECT 85.780 168.030 85.920 169.190 ;
        RECT 86.700 169.190 100.640 169.330 ;
        RECT 101.905 169.330 102.195 169.375 ;
        RECT 105.145 169.330 105.795 169.375 ;
        RECT 106.020 169.330 106.160 169.530 ;
        RECT 106.850 169.470 107.170 169.530 ;
        RECT 101.905 169.190 106.160 169.330 ;
        RECT 106.390 169.330 106.710 169.390 ;
        RECT 107.785 169.330 108.075 169.375 ;
        RECT 106.390 169.190 108.075 169.330 ;
        RECT 86.700 168.695 86.840 169.190 ;
        RECT 99.950 169.130 100.270 169.190 ;
        RECT 101.905 169.145 102.495 169.190 ;
        RECT 105.145 169.145 105.795 169.190 ;
        RECT 89.370 168.990 89.690 169.050 ;
        RECT 89.845 168.990 90.135 169.035 ;
        RECT 89.370 168.850 90.135 168.990 ;
        RECT 89.370 168.790 89.690 168.850 ;
        RECT 89.845 168.805 90.135 168.850 ;
        RECT 92.590 168.790 92.910 169.050 ;
        RECT 95.810 168.790 96.130 169.050 ;
        RECT 98.110 168.790 98.430 169.050 ;
        RECT 99.140 168.990 99.430 169.035 ;
        RECT 99.120 168.805 99.430 168.990 ;
        RECT 102.205 168.830 102.495 169.145 ;
        RECT 106.390 169.130 106.710 169.190 ;
        RECT 107.785 169.145 108.075 169.190 ;
        RECT 103.285 168.990 103.575 169.035 ;
        RECT 106.865 168.990 107.155 169.035 ;
        RECT 108.700 168.990 108.990 169.035 ;
        RECT 103.285 168.850 108.990 168.990 ;
        RECT 103.285 168.805 103.575 168.850 ;
        RECT 106.865 168.805 107.155 168.850 ;
        RECT 108.700 168.805 108.990 168.850 ;
        RECT 86.625 168.465 86.915 168.695 ;
        RECT 95.900 168.650 96.040 168.790 ;
        RECT 89.460 168.510 96.040 168.650 ;
        RECT 96.270 168.650 96.590 168.710 ;
        RECT 97.205 168.650 97.495 168.695 ;
        RECT 99.120 168.650 99.260 168.805 ;
        RECT 96.270 168.510 99.260 168.650 ;
        RECT 89.460 168.355 89.600 168.510 ;
        RECT 96.270 168.450 96.590 168.510 ;
        RECT 97.205 168.465 97.495 168.510 ;
        RECT 99.965 168.465 100.255 168.695 ;
        RECT 109.165 168.650 109.455 168.695 ;
        RECT 109.610 168.650 109.930 168.710 ;
        RECT 109.165 168.510 109.930 168.650 ;
        RECT 109.165 168.465 109.455 168.510 ;
        RECT 89.385 168.125 89.675 168.355 ;
        RECT 98.585 168.310 98.875 168.355 ;
        RECT 100.040 168.310 100.180 168.465 ;
        RECT 109.610 168.450 109.930 168.510 ;
        RECT 92.220 168.170 98.875 168.310 ;
        RECT 85.230 167.770 85.550 168.030 ;
        RECT 85.690 167.770 86.010 168.030 ;
        RECT 86.150 167.770 86.470 168.030 ;
        RECT 88.465 167.970 88.755 168.015 ;
        RECT 92.220 167.970 92.360 168.170 ;
        RECT 98.585 168.125 98.875 168.170 ;
        RECT 99.120 168.170 100.180 168.310 ;
        RECT 103.285 168.310 103.575 168.355 ;
        RECT 106.405 168.310 106.695 168.355 ;
        RECT 108.295 168.310 108.585 168.355 ;
        RECT 103.285 168.170 108.585 168.310 ;
        RECT 99.120 168.030 99.260 168.170 ;
        RECT 103.285 168.125 103.575 168.170 ;
        RECT 106.405 168.125 106.695 168.170 ;
        RECT 108.295 168.125 108.585 168.170 ;
        RECT 88.465 167.830 92.360 167.970 ;
        RECT 92.590 167.970 92.910 168.030 ;
        RECT 94.445 167.970 94.735 168.015 ;
        RECT 92.590 167.830 94.735 167.970 ;
        RECT 88.465 167.785 88.755 167.830 ;
        RECT 92.590 167.770 92.910 167.830 ;
        RECT 94.445 167.785 94.735 167.830 ;
        RECT 96.730 167.970 97.050 168.030 ;
        RECT 99.030 167.970 99.350 168.030 ;
        RECT 96.730 167.830 99.350 167.970 ;
        RECT 96.730 167.770 97.050 167.830 ;
        RECT 99.030 167.770 99.350 167.830 ;
        RECT 67.680 167.150 121.960 167.630 ;
        RECT 83.480 166.810 88.680 166.950 ;
        RECT 83.480 166.670 83.620 166.810 ;
        RECT 83.390 166.410 83.710 166.670 ;
        RECT 86.625 166.610 86.915 166.655 ;
        RECT 86.625 166.470 88.220 166.610 ;
        RECT 86.625 166.425 86.915 166.470 ;
        RECT 87.530 166.070 87.850 166.330 ;
        RECT 85.230 165.730 85.550 165.990 ;
        RECT 86.150 165.930 86.470 165.990 ;
        RECT 88.080 165.975 88.220 166.470 ;
        RECT 88.540 166.315 88.680 166.810 ;
        RECT 99.950 166.750 100.270 167.010 ;
        RECT 88.930 166.610 89.220 166.655 ;
        RECT 91.250 166.610 91.540 166.655 ;
        RECT 92.630 166.610 92.920 166.655 ;
        RECT 88.930 166.470 92.920 166.610 ;
        RECT 88.930 166.425 89.220 166.470 ;
        RECT 91.250 166.425 91.540 166.470 ;
        RECT 92.630 166.425 92.920 166.470 ;
        RECT 88.465 166.085 88.755 166.315 ;
        RECT 89.370 166.070 89.690 166.330 ;
        RECT 87.085 165.930 87.375 165.975 ;
        RECT 86.150 165.790 87.375 165.930 ;
        RECT 86.150 165.730 86.470 165.790 ;
        RECT 87.085 165.745 87.375 165.790 ;
        RECT 88.005 165.745 88.295 165.975 ;
        RECT 89.460 165.930 89.600 166.070 ;
        RECT 88.540 165.790 89.600 165.930 ;
        RECT 64.990 165.590 65.310 165.650 ;
        RECT 85.320 165.590 85.460 165.730 ;
        RECT 86.625 165.590 86.915 165.635 ;
        RECT 88.540 165.590 88.680 165.790 ;
        RECT 89.830 165.730 90.150 165.990 ;
        RECT 100.040 165.930 100.180 166.750 ;
        RECT 102.265 165.930 102.555 165.975 ;
        RECT 100.040 165.790 102.555 165.930 ;
        RECT 102.265 165.745 102.555 165.790 ;
        RECT 64.990 165.450 86.380 165.590 ;
        RECT 64.990 165.390 65.310 165.450 ;
        RECT 85.690 165.050 86.010 165.310 ;
        RECT 86.240 165.250 86.380 165.450 ;
        RECT 86.625 165.450 88.680 165.590 ;
        RECT 89.390 165.590 89.680 165.635 ;
        RECT 90.790 165.590 91.080 165.635 ;
        RECT 92.630 165.590 92.920 165.635 ;
        RECT 89.390 165.450 92.920 165.590 ;
        RECT 86.625 165.405 86.915 165.450 ;
        RECT 89.390 165.405 89.680 165.450 ;
        RECT 90.790 165.405 91.080 165.450 ;
        RECT 92.630 165.405 92.920 165.450 ;
        RECT 95.365 165.250 95.655 165.295 ;
        RECT 95.810 165.250 96.130 165.310 ;
        RECT 86.240 165.110 96.130 165.250 ;
        RECT 95.365 165.065 95.655 165.110 ;
        RECT 95.810 165.050 96.130 165.110 ;
        RECT 99.490 165.250 99.810 165.310 ;
        RECT 101.345 165.250 101.635 165.295 ;
        RECT 99.490 165.110 101.635 165.250 ;
        RECT 99.490 165.050 99.810 165.110 ;
        RECT 101.345 165.065 101.635 165.110 ;
        RECT 67.680 164.430 122.760 164.910 ;
        RECT 83.850 164.030 84.170 164.290 ;
        RECT 89.830 164.230 90.150 164.290 ;
        RECT 90.765 164.230 91.055 164.275 ;
        RECT 89.830 164.090 91.055 164.230 ;
        RECT 89.830 164.030 90.150 164.090 ;
        RECT 90.765 164.045 91.055 164.090 ;
        RECT 83.940 163.890 84.080 164.030 ;
        RECT 93.985 163.890 94.275 163.935 ;
        RECT 99.490 163.890 99.810 163.950 ;
        RECT 83.940 163.750 99.810 163.890 ;
        RECT 93.985 163.705 94.275 163.750 ;
        RECT 99.490 163.690 99.810 163.750 ;
        RECT 100.400 163.890 100.690 163.935 ;
        RECT 102.240 163.890 102.530 163.935 ;
        RECT 103.640 163.890 103.930 163.935 ;
        RECT 100.400 163.750 103.930 163.890 ;
        RECT 100.400 163.705 100.690 163.750 ;
        RECT 102.240 163.705 102.530 163.750 ;
        RECT 103.640 163.705 103.930 163.750 ;
        RECT 85.690 163.550 86.010 163.610 ;
        RECT 91.685 163.550 91.975 163.595 ;
        RECT 85.690 163.410 91.440 163.550 ;
        RECT 85.690 163.350 86.010 163.410 ;
        RECT 91.300 163.210 91.440 163.410 ;
        RECT 91.685 163.410 94.660 163.550 ;
        RECT 91.685 163.365 91.975 163.410 ;
        RECT 91.300 163.070 92.360 163.210 ;
        RECT 92.220 162.870 92.360 163.070 ;
        RECT 92.590 163.010 92.910 163.270 ;
        RECT 93.065 163.025 93.355 163.255 ;
        RECT 93.140 162.870 93.280 163.025 ;
        RECT 92.220 162.730 93.280 162.870 ;
        RECT 93.140 162.530 93.280 162.730 ;
        RECT 93.985 162.870 94.275 162.915 ;
        RECT 94.520 162.870 94.660 163.410 ;
        RECT 94.905 163.365 95.195 163.595 ;
        RECT 95.365 163.550 95.655 163.595 ;
        RECT 95.810 163.550 96.130 163.610 ;
        RECT 95.365 163.410 96.130 163.550 ;
        RECT 95.365 163.365 95.655 163.410 ;
        RECT 93.985 162.730 94.660 162.870 ;
        RECT 94.980 163.210 95.120 163.365 ;
        RECT 95.810 163.350 96.130 163.410 ;
        RECT 94.980 163.070 97.880 163.210 ;
        RECT 93.985 162.685 94.275 162.730 ;
        RECT 94.980 162.530 95.120 163.070 ;
        RECT 97.740 162.575 97.880 163.070 ;
        RECT 103.170 163.010 103.490 163.270 ;
        RECT 104.565 163.210 104.855 163.255 ;
        RECT 109.150 163.210 109.470 163.270 ;
        RECT 104.565 163.070 109.470 163.210 ;
        RECT 104.565 163.025 104.855 163.070 ;
        RECT 109.150 163.010 109.470 163.070 ;
        RECT 100.400 162.870 100.690 162.915 ;
        RECT 101.780 162.870 102.070 162.915 ;
        RECT 104.100 162.870 104.390 162.915 ;
        RECT 100.400 162.730 104.390 162.870 ;
        RECT 100.400 162.685 100.690 162.730 ;
        RECT 101.780 162.685 102.070 162.730 ;
        RECT 104.100 162.685 104.390 162.730 ;
        RECT 93.140 162.390 95.120 162.530 ;
        RECT 97.665 162.530 97.955 162.575 ;
        RECT 99.030 162.530 99.350 162.590 ;
        RECT 103.630 162.530 103.950 162.590 ;
        RECT 97.665 162.390 103.950 162.530 ;
        RECT 97.665 162.345 97.955 162.390 ;
        RECT 99.030 162.330 99.350 162.390 ;
        RECT 103.630 162.330 103.950 162.390 ;
        RECT 67.680 161.710 121.960 162.190 ;
        RECT 83.390 161.310 83.710 161.570 ;
        RECT 100.885 161.510 101.175 161.555 ;
        RECT 103.170 161.510 103.490 161.570 ;
        RECT 100.885 161.370 103.490 161.510 ;
        RECT 100.885 161.325 101.175 161.370 ;
        RECT 103.170 161.310 103.490 161.370 ;
        RECT 109.150 161.510 109.470 161.570 ;
        RECT 113.305 161.510 113.595 161.555 ;
        RECT 109.150 161.370 113.595 161.510 ;
        RECT 109.150 161.310 109.470 161.370 ;
        RECT 113.305 161.325 113.595 161.370 ;
        RECT 98.125 160.830 98.415 160.875 ;
        RECT 101.805 160.830 102.095 160.875 ;
        RECT 98.125 160.690 102.095 160.830 ;
        RECT 98.125 160.645 98.415 160.690 ;
        RECT 101.805 160.645 102.095 160.690 ;
        RECT 99.490 160.490 99.810 160.550 ;
        RECT 101.345 160.490 101.635 160.535 ;
        RECT 99.490 160.350 101.635 160.490 ;
        RECT 99.490 160.290 99.810 160.350 ;
        RECT 101.345 160.305 101.635 160.350 ;
        RECT 102.265 160.490 102.555 160.535 ;
        RECT 103.630 160.490 103.950 160.550 ;
        RECT 102.265 160.350 103.950 160.490 ;
        RECT 102.265 160.305 102.555 160.350 ;
        RECT 103.630 160.290 103.950 160.350 ;
        RECT 89.845 160.150 90.135 160.195 ;
        RECT 100.410 160.150 100.730 160.210 ;
        RECT 106.865 160.150 107.155 160.195 ;
        RECT 89.845 160.010 107.155 160.150 ;
        RECT 89.845 159.965 90.135 160.010 ;
        RECT 100.410 159.950 100.730 160.010 ;
        RECT 106.865 159.965 107.155 160.010 ;
        RECT 67.680 158.990 122.760 159.470 ;
        RECT 85.690 102.970 86.230 103.390 ;
        RECT 85.830 101.540 86.050 102.970 ;
        RECT 89.360 102.890 90.030 103.450 ;
        RECT 85.835 94.075 86.045 101.540 ;
        RECT 89.525 97.305 89.735 102.890 ;
        RECT 92.760 102.880 93.430 103.440 ;
        RECT 96.520 103.255 97.190 103.470 ;
        RECT 95.430 103.045 97.190 103.255 ;
        RECT 89.525 97.095 91.040 97.305 ;
        RECT 85.835 93.865 88.935 94.075 ;
        RECT 81.780 91.380 83.060 91.800 ;
        RECT 86.450 91.380 86.970 92.240 ;
        RECT 88.725 92.130 88.935 93.865 ;
        RECT 81.780 90.860 86.970 91.380 ;
        RECT 81.780 90.650 83.060 90.860 ;
        RECT 86.450 90.540 86.970 90.860 ;
        RECT 88.690 90.775 88.935 92.130 ;
        RECT 90.830 91.980 91.040 97.095 ;
        RECT 93.120 91.980 93.330 102.880 ;
        RECT 86.600 90.065 86.830 90.540 ;
        RECT 88.690 90.025 88.920 90.775 ;
        RECT 90.810 89.875 91.040 91.980 ;
        RECT 93.080 90.640 93.330 91.980 ;
        RECT 95.430 92.230 95.640 103.045 ;
        RECT 96.520 102.910 97.190 103.045 ;
        RECT 93.080 89.875 93.310 90.640 ;
        RECT 95.430 90.610 95.680 92.230 ;
        RECT 95.450 90.125 95.680 90.610 ;
        RECT 86.600 75.700 86.830 76.325 ;
        RECT 88.690 75.700 88.920 76.285 ;
        RECT 86.280 74.850 89.180 75.700 ;
        RECT 90.810 75.530 91.040 76.135 ;
        RECT 93.080 75.730 93.310 76.135 ;
        RECT 95.450 75.790 95.680 76.385 ;
        RECT 86.600 74.220 86.830 74.850 ;
        RECT 87.275 63.455 88.105 74.850 ;
        RECT 88.690 74.180 88.920 74.850 ;
        RECT 90.560 71.020 91.260 75.530 ;
        RECT 92.920 72.550 93.620 75.730 ;
        RECT 95.340 73.440 96.040 75.790 ;
        RECT 95.340 72.740 106.000 73.440 ;
        RECT 92.920 71.850 94.720 72.550 ;
        RECT 90.560 70.320 92.440 71.020 ;
        RECT 92.920 70.520 93.620 71.850 ;
        RECT 90.810 69.355 91.040 70.320 ;
        RECT 87.280 61.620 88.100 63.455 ;
        RECT 90.810 61.620 91.040 62.455 ;
        RECT 87.280 60.800 91.360 61.620 ;
        RECT 91.750 61.450 92.430 70.320 ;
        RECT 93.180 69.505 93.410 70.520 ;
        RECT 93.180 61.450 93.410 62.605 ;
        RECT 94.030 61.520 94.710 71.850 ;
        RECT 95.340 70.580 96.040 72.740 ;
        RECT 95.550 69.255 95.780 70.580 ;
        RECT 95.550 61.520 95.780 62.355 ;
        RECT 90.810 60.350 91.040 60.800 ;
        RECT 91.750 60.770 93.700 61.450 ;
        RECT 94.030 60.840 96.020 61.520 ;
        RECT 93.180 60.500 93.410 60.770 ;
        RECT 95.550 60.250 95.780 60.840 ;
      LAYER via ;
        RECT 80.480 213.500 80.740 213.760 ;
        RECT 80.800 213.500 81.060 213.760 ;
        RECT 81.120 213.500 81.380 213.760 ;
        RECT 81.440 213.500 81.700 213.760 ;
        RECT 81.760 213.500 82.020 213.760 ;
        RECT 94.050 213.500 94.310 213.760 ;
        RECT 94.370 213.500 94.630 213.760 ;
        RECT 94.690 213.500 94.950 213.760 ;
        RECT 95.010 213.500 95.270 213.760 ;
        RECT 95.330 213.500 95.590 213.760 ;
        RECT 107.620 213.500 107.880 213.760 ;
        RECT 107.940 213.500 108.200 213.760 ;
        RECT 108.260 213.500 108.520 213.760 ;
        RECT 108.580 213.500 108.840 213.760 ;
        RECT 108.900 213.500 109.160 213.760 ;
        RECT 121.190 213.500 121.450 213.760 ;
        RECT 121.510 213.500 121.770 213.760 ;
        RECT 121.830 213.500 122.090 213.760 ;
        RECT 122.150 213.500 122.410 213.760 ;
        RECT 122.470 213.500 122.730 213.760 ;
        RECT 73.695 210.780 73.955 211.040 ;
        RECT 74.015 210.780 74.275 211.040 ;
        RECT 74.335 210.780 74.595 211.040 ;
        RECT 74.655 210.780 74.915 211.040 ;
        RECT 74.975 210.780 75.235 211.040 ;
        RECT 87.265 210.780 87.525 211.040 ;
        RECT 87.585 210.780 87.845 211.040 ;
        RECT 87.905 210.780 88.165 211.040 ;
        RECT 88.225 210.780 88.485 211.040 ;
        RECT 88.545 210.780 88.805 211.040 ;
        RECT 100.835 210.780 101.095 211.040 ;
        RECT 101.155 210.780 101.415 211.040 ;
        RECT 101.475 210.780 101.735 211.040 ;
        RECT 101.795 210.780 102.055 211.040 ;
        RECT 102.115 210.780 102.375 211.040 ;
        RECT 114.405 210.780 114.665 211.040 ;
        RECT 114.725 210.780 114.985 211.040 ;
        RECT 115.045 210.780 115.305 211.040 ;
        RECT 115.365 210.780 115.625 211.040 ;
        RECT 115.685 210.780 115.945 211.040 ;
        RECT 80.480 208.060 80.740 208.320 ;
        RECT 80.800 208.060 81.060 208.320 ;
        RECT 81.120 208.060 81.380 208.320 ;
        RECT 81.440 208.060 81.700 208.320 ;
        RECT 81.760 208.060 82.020 208.320 ;
        RECT 94.050 208.060 94.310 208.320 ;
        RECT 94.370 208.060 94.630 208.320 ;
        RECT 94.690 208.060 94.950 208.320 ;
        RECT 95.010 208.060 95.270 208.320 ;
        RECT 95.330 208.060 95.590 208.320 ;
        RECT 107.620 208.060 107.880 208.320 ;
        RECT 107.940 208.060 108.200 208.320 ;
        RECT 108.260 208.060 108.520 208.320 ;
        RECT 108.580 208.060 108.840 208.320 ;
        RECT 108.900 208.060 109.160 208.320 ;
        RECT 121.190 208.060 121.450 208.320 ;
        RECT 121.510 208.060 121.770 208.320 ;
        RECT 121.830 208.060 122.090 208.320 ;
        RECT 122.150 208.060 122.410 208.320 ;
        RECT 122.470 208.060 122.730 208.320 ;
        RECT 73.695 205.340 73.955 205.600 ;
        RECT 74.015 205.340 74.275 205.600 ;
        RECT 74.335 205.340 74.595 205.600 ;
        RECT 74.655 205.340 74.915 205.600 ;
        RECT 74.975 205.340 75.235 205.600 ;
        RECT 87.265 205.340 87.525 205.600 ;
        RECT 87.585 205.340 87.845 205.600 ;
        RECT 87.905 205.340 88.165 205.600 ;
        RECT 88.225 205.340 88.485 205.600 ;
        RECT 88.545 205.340 88.805 205.600 ;
        RECT 100.835 205.340 101.095 205.600 ;
        RECT 101.155 205.340 101.415 205.600 ;
        RECT 101.475 205.340 101.735 205.600 ;
        RECT 101.795 205.340 102.055 205.600 ;
        RECT 102.115 205.340 102.375 205.600 ;
        RECT 114.405 205.340 114.665 205.600 ;
        RECT 114.725 205.340 114.985 205.600 ;
        RECT 115.045 205.340 115.305 205.600 ;
        RECT 115.365 205.340 115.625 205.600 ;
        RECT 115.685 205.340 115.945 205.600 ;
        RECT 80.480 202.620 80.740 202.880 ;
        RECT 80.800 202.620 81.060 202.880 ;
        RECT 81.120 202.620 81.380 202.880 ;
        RECT 81.440 202.620 81.700 202.880 ;
        RECT 81.760 202.620 82.020 202.880 ;
        RECT 94.050 202.620 94.310 202.880 ;
        RECT 94.370 202.620 94.630 202.880 ;
        RECT 94.690 202.620 94.950 202.880 ;
        RECT 95.010 202.620 95.270 202.880 ;
        RECT 95.330 202.620 95.590 202.880 ;
        RECT 107.620 202.620 107.880 202.880 ;
        RECT 107.940 202.620 108.200 202.880 ;
        RECT 108.260 202.620 108.520 202.880 ;
        RECT 108.580 202.620 108.840 202.880 ;
        RECT 108.900 202.620 109.160 202.880 ;
        RECT 121.190 202.620 121.450 202.880 ;
        RECT 121.510 202.620 121.770 202.880 ;
        RECT 121.830 202.620 122.090 202.880 ;
        RECT 122.150 202.620 122.410 202.880 ;
        RECT 122.470 202.620 122.730 202.880 ;
        RECT 73.695 199.900 73.955 200.160 ;
        RECT 74.015 199.900 74.275 200.160 ;
        RECT 74.335 199.900 74.595 200.160 ;
        RECT 74.655 199.900 74.915 200.160 ;
        RECT 74.975 199.900 75.235 200.160 ;
        RECT 87.265 199.900 87.525 200.160 ;
        RECT 87.585 199.900 87.845 200.160 ;
        RECT 87.905 199.900 88.165 200.160 ;
        RECT 88.225 199.900 88.485 200.160 ;
        RECT 88.545 199.900 88.805 200.160 ;
        RECT 100.835 199.900 101.095 200.160 ;
        RECT 101.155 199.900 101.415 200.160 ;
        RECT 101.475 199.900 101.735 200.160 ;
        RECT 101.795 199.900 102.055 200.160 ;
        RECT 102.115 199.900 102.375 200.160 ;
        RECT 114.405 199.900 114.665 200.160 ;
        RECT 114.725 199.900 114.985 200.160 ;
        RECT 115.045 199.900 115.305 200.160 ;
        RECT 115.365 199.900 115.625 200.160 ;
        RECT 115.685 199.900 115.945 200.160 ;
        RECT 80.480 197.180 80.740 197.440 ;
        RECT 80.800 197.180 81.060 197.440 ;
        RECT 81.120 197.180 81.380 197.440 ;
        RECT 81.440 197.180 81.700 197.440 ;
        RECT 81.760 197.180 82.020 197.440 ;
        RECT 94.050 197.180 94.310 197.440 ;
        RECT 94.370 197.180 94.630 197.440 ;
        RECT 94.690 197.180 94.950 197.440 ;
        RECT 95.010 197.180 95.270 197.440 ;
        RECT 95.330 197.180 95.590 197.440 ;
        RECT 107.620 197.180 107.880 197.440 ;
        RECT 107.940 197.180 108.200 197.440 ;
        RECT 108.260 197.180 108.520 197.440 ;
        RECT 108.580 197.180 108.840 197.440 ;
        RECT 108.900 197.180 109.160 197.440 ;
        RECT 121.190 197.180 121.450 197.440 ;
        RECT 121.510 197.180 121.770 197.440 ;
        RECT 121.830 197.180 122.090 197.440 ;
        RECT 122.150 197.180 122.410 197.440 ;
        RECT 122.470 197.180 122.730 197.440 ;
        RECT 73.695 194.460 73.955 194.720 ;
        RECT 74.015 194.460 74.275 194.720 ;
        RECT 74.335 194.460 74.595 194.720 ;
        RECT 74.655 194.460 74.915 194.720 ;
        RECT 74.975 194.460 75.235 194.720 ;
        RECT 87.265 194.460 87.525 194.720 ;
        RECT 87.585 194.460 87.845 194.720 ;
        RECT 87.905 194.460 88.165 194.720 ;
        RECT 88.225 194.460 88.485 194.720 ;
        RECT 88.545 194.460 88.805 194.720 ;
        RECT 100.835 194.460 101.095 194.720 ;
        RECT 101.155 194.460 101.415 194.720 ;
        RECT 101.475 194.460 101.735 194.720 ;
        RECT 101.795 194.460 102.055 194.720 ;
        RECT 102.115 194.460 102.375 194.720 ;
        RECT 114.405 194.460 114.665 194.720 ;
        RECT 114.725 194.460 114.985 194.720 ;
        RECT 115.045 194.460 115.305 194.720 ;
        RECT 115.365 194.460 115.625 194.720 ;
        RECT 115.685 194.460 115.945 194.720 ;
        RECT 78.820 193.950 79.080 194.210 ;
        RECT 92.620 193.950 92.880 194.210 ;
        RECT 80.480 191.740 80.740 192.000 ;
        RECT 80.800 191.740 81.060 192.000 ;
        RECT 81.120 191.740 81.380 192.000 ;
        RECT 81.440 191.740 81.700 192.000 ;
        RECT 81.760 191.740 82.020 192.000 ;
        RECT 94.050 191.740 94.310 192.000 ;
        RECT 94.370 191.740 94.630 192.000 ;
        RECT 94.690 191.740 94.950 192.000 ;
        RECT 95.010 191.740 95.270 192.000 ;
        RECT 95.330 191.740 95.590 192.000 ;
        RECT 107.620 191.740 107.880 192.000 ;
        RECT 107.940 191.740 108.200 192.000 ;
        RECT 108.260 191.740 108.520 192.000 ;
        RECT 108.580 191.740 108.840 192.000 ;
        RECT 108.900 191.740 109.160 192.000 ;
        RECT 121.190 191.740 121.450 192.000 ;
        RECT 121.510 191.740 121.770 192.000 ;
        RECT 121.830 191.740 122.090 192.000 ;
        RECT 122.150 191.740 122.410 192.000 ;
        RECT 122.470 191.740 122.730 192.000 ;
        RECT 73.695 189.020 73.955 189.280 ;
        RECT 74.015 189.020 74.275 189.280 ;
        RECT 74.335 189.020 74.595 189.280 ;
        RECT 74.655 189.020 74.915 189.280 ;
        RECT 74.975 189.020 75.235 189.280 ;
        RECT 87.265 189.020 87.525 189.280 ;
        RECT 87.585 189.020 87.845 189.280 ;
        RECT 87.905 189.020 88.165 189.280 ;
        RECT 88.225 189.020 88.485 189.280 ;
        RECT 88.545 189.020 88.805 189.280 ;
        RECT 100.835 189.020 101.095 189.280 ;
        RECT 101.155 189.020 101.415 189.280 ;
        RECT 101.475 189.020 101.735 189.280 ;
        RECT 101.795 189.020 102.055 189.280 ;
        RECT 102.115 189.020 102.375 189.280 ;
        RECT 114.405 189.020 114.665 189.280 ;
        RECT 114.725 189.020 114.985 189.280 ;
        RECT 115.045 189.020 115.305 189.280 ;
        RECT 115.365 189.020 115.625 189.280 ;
        RECT 115.685 189.020 115.945 189.280 ;
        RECT 80.480 186.300 80.740 186.560 ;
        RECT 80.800 186.300 81.060 186.560 ;
        RECT 81.120 186.300 81.380 186.560 ;
        RECT 81.440 186.300 81.700 186.560 ;
        RECT 81.760 186.300 82.020 186.560 ;
        RECT 94.050 186.300 94.310 186.560 ;
        RECT 94.370 186.300 94.630 186.560 ;
        RECT 94.690 186.300 94.950 186.560 ;
        RECT 95.010 186.300 95.270 186.560 ;
        RECT 95.330 186.300 95.590 186.560 ;
        RECT 107.620 186.300 107.880 186.560 ;
        RECT 107.940 186.300 108.200 186.560 ;
        RECT 108.260 186.300 108.520 186.560 ;
        RECT 108.580 186.300 108.840 186.560 ;
        RECT 108.900 186.300 109.160 186.560 ;
        RECT 121.190 186.300 121.450 186.560 ;
        RECT 121.510 186.300 121.770 186.560 ;
        RECT 121.830 186.300 122.090 186.560 ;
        RECT 122.150 186.300 122.410 186.560 ;
        RECT 122.470 186.300 122.730 186.560 ;
        RECT 73.695 183.580 73.955 183.840 ;
        RECT 74.015 183.580 74.275 183.840 ;
        RECT 74.335 183.580 74.595 183.840 ;
        RECT 74.655 183.580 74.915 183.840 ;
        RECT 74.975 183.580 75.235 183.840 ;
        RECT 87.265 183.580 87.525 183.840 ;
        RECT 87.585 183.580 87.845 183.840 ;
        RECT 87.905 183.580 88.165 183.840 ;
        RECT 88.225 183.580 88.485 183.840 ;
        RECT 88.545 183.580 88.805 183.840 ;
        RECT 100.835 183.580 101.095 183.840 ;
        RECT 101.155 183.580 101.415 183.840 ;
        RECT 101.475 183.580 101.735 183.840 ;
        RECT 101.795 183.580 102.055 183.840 ;
        RECT 102.115 183.580 102.375 183.840 ;
        RECT 114.405 183.580 114.665 183.840 ;
        RECT 114.725 183.580 114.985 183.840 ;
        RECT 115.045 183.580 115.305 183.840 ;
        RECT 115.365 183.580 115.625 183.840 ;
        RECT 115.685 183.580 115.945 183.840 ;
        RECT 80.480 180.860 80.740 181.120 ;
        RECT 80.800 180.860 81.060 181.120 ;
        RECT 81.120 180.860 81.380 181.120 ;
        RECT 81.440 180.860 81.700 181.120 ;
        RECT 81.760 180.860 82.020 181.120 ;
        RECT 94.050 180.860 94.310 181.120 ;
        RECT 94.370 180.860 94.630 181.120 ;
        RECT 94.690 180.860 94.950 181.120 ;
        RECT 95.010 180.860 95.270 181.120 ;
        RECT 95.330 180.860 95.590 181.120 ;
        RECT 107.620 180.860 107.880 181.120 ;
        RECT 107.940 180.860 108.200 181.120 ;
        RECT 108.260 180.860 108.520 181.120 ;
        RECT 108.580 180.860 108.840 181.120 ;
        RECT 108.900 180.860 109.160 181.120 ;
        RECT 121.190 180.860 121.450 181.120 ;
        RECT 121.510 180.860 121.770 181.120 ;
        RECT 121.830 180.860 122.090 181.120 ;
        RECT 122.150 180.860 122.410 181.120 ;
        RECT 122.470 180.860 122.730 181.120 ;
        RECT 73.695 178.140 73.955 178.400 ;
        RECT 74.015 178.140 74.275 178.400 ;
        RECT 74.335 178.140 74.595 178.400 ;
        RECT 74.655 178.140 74.915 178.400 ;
        RECT 74.975 178.140 75.235 178.400 ;
        RECT 87.265 178.140 87.525 178.400 ;
        RECT 87.585 178.140 87.845 178.400 ;
        RECT 87.905 178.140 88.165 178.400 ;
        RECT 88.225 178.140 88.485 178.400 ;
        RECT 88.545 178.140 88.805 178.400 ;
        RECT 100.835 178.140 101.095 178.400 ;
        RECT 101.155 178.140 101.415 178.400 ;
        RECT 101.475 178.140 101.735 178.400 ;
        RECT 101.795 178.140 102.055 178.400 ;
        RECT 102.115 178.140 102.375 178.400 ;
        RECT 114.405 178.140 114.665 178.400 ;
        RECT 114.725 178.140 114.985 178.400 ;
        RECT 115.045 178.140 115.305 178.400 ;
        RECT 115.365 178.140 115.625 178.400 ;
        RECT 115.685 178.140 115.945 178.400 ;
        RECT 99.060 176.950 99.320 177.210 ;
        RECT 122.980 176.950 123.240 177.210 ;
        RECT 80.480 175.420 80.740 175.680 ;
        RECT 80.800 175.420 81.060 175.680 ;
        RECT 81.120 175.420 81.380 175.680 ;
        RECT 81.440 175.420 81.700 175.680 ;
        RECT 81.760 175.420 82.020 175.680 ;
        RECT 94.050 175.420 94.310 175.680 ;
        RECT 94.370 175.420 94.630 175.680 ;
        RECT 94.690 175.420 94.950 175.680 ;
        RECT 95.010 175.420 95.270 175.680 ;
        RECT 95.330 175.420 95.590 175.680 ;
        RECT 107.620 175.420 107.880 175.680 ;
        RECT 107.940 175.420 108.200 175.680 ;
        RECT 108.260 175.420 108.520 175.680 ;
        RECT 108.580 175.420 108.840 175.680 ;
        RECT 108.900 175.420 109.160 175.680 ;
        RECT 121.190 175.420 121.450 175.680 ;
        RECT 121.510 175.420 121.770 175.680 ;
        RECT 121.830 175.420 122.090 175.680 ;
        RECT 122.150 175.420 122.410 175.680 ;
        RECT 122.470 175.420 122.730 175.680 ;
        RECT 99.060 174.910 99.320 175.170 ;
        RECT 96.300 174.570 96.560 174.830 ;
        RECT 93.540 173.890 93.800 174.150 ;
        RECT 105.500 173.890 105.760 174.150 ;
        RECT 109.640 173.890 109.900 174.150 ;
        RECT 121.140 173.890 121.400 174.150 ;
        RECT 93.080 173.210 93.340 173.470 ;
        RECT 96.760 173.210 97.020 173.470 ;
        RECT 117.920 173.210 118.180 173.470 ;
        RECT 73.695 172.700 73.955 172.960 ;
        RECT 74.015 172.700 74.275 172.960 ;
        RECT 74.335 172.700 74.595 172.960 ;
        RECT 74.655 172.700 74.915 172.960 ;
        RECT 74.975 172.700 75.235 172.960 ;
        RECT 87.265 172.700 87.525 172.960 ;
        RECT 87.585 172.700 87.845 172.960 ;
        RECT 87.905 172.700 88.165 172.960 ;
        RECT 88.225 172.700 88.485 172.960 ;
        RECT 88.545 172.700 88.805 172.960 ;
        RECT 100.835 172.700 101.095 172.960 ;
        RECT 101.155 172.700 101.415 172.960 ;
        RECT 101.475 172.700 101.735 172.960 ;
        RECT 101.795 172.700 102.055 172.960 ;
        RECT 102.115 172.700 102.375 172.960 ;
        RECT 114.405 172.700 114.665 172.960 ;
        RECT 114.725 172.700 114.985 172.960 ;
        RECT 115.045 172.700 115.305 172.960 ;
        RECT 115.365 172.700 115.625 172.960 ;
        RECT 115.685 172.700 115.945 172.960 ;
        RECT 105.500 172.190 105.760 172.450 ;
        RECT 117.920 172.190 118.180 172.450 ;
        RECT 86.640 171.170 86.900 171.430 ;
        RECT 92.620 171.170 92.880 171.430 ;
        RECT 95.840 171.170 96.100 171.430 ;
        RECT 83.420 170.490 83.680 170.750 ;
        RECT 92.620 170.490 92.880 170.750 ;
        RECT 93.540 170.490 93.800 170.750 ;
        RECT 98.600 170.490 98.860 170.750 ;
        RECT 100.440 170.490 100.700 170.750 ;
        RECT 106.420 170.490 106.680 170.750 ;
        RECT 106.880 170.490 107.140 170.750 ;
        RECT 80.480 169.980 80.740 170.240 ;
        RECT 80.800 169.980 81.060 170.240 ;
        RECT 81.120 169.980 81.380 170.240 ;
        RECT 81.440 169.980 81.700 170.240 ;
        RECT 81.760 169.980 82.020 170.240 ;
        RECT 94.050 169.980 94.310 170.240 ;
        RECT 94.370 169.980 94.630 170.240 ;
        RECT 94.690 169.980 94.950 170.240 ;
        RECT 95.010 169.980 95.270 170.240 ;
        RECT 95.330 169.980 95.590 170.240 ;
        RECT 107.620 169.980 107.880 170.240 ;
        RECT 107.940 169.980 108.200 170.240 ;
        RECT 108.260 169.980 108.520 170.240 ;
        RECT 108.580 169.980 108.840 170.240 ;
        RECT 108.900 169.980 109.160 170.240 ;
        RECT 121.190 169.980 121.450 170.240 ;
        RECT 121.510 169.980 121.770 170.240 ;
        RECT 121.830 169.980 122.090 170.240 ;
        RECT 122.150 169.980 122.410 170.240 ;
        RECT 122.470 169.980 122.730 170.240 ;
        RECT 93.080 169.470 93.340 169.730 ;
        RECT 98.600 169.470 98.860 169.730 ;
        RECT 85.260 168.790 85.520 169.050 ;
        RECT 83.880 168.450 84.140 168.710 ;
        RECT 99.980 169.130 100.240 169.390 ;
        RECT 106.880 169.470 107.140 169.730 ;
        RECT 89.400 168.790 89.660 169.050 ;
        RECT 92.620 168.790 92.880 169.050 ;
        RECT 95.840 168.790 96.100 169.050 ;
        RECT 98.140 168.790 98.400 169.050 ;
        RECT 106.420 169.130 106.680 169.390 ;
        RECT 96.300 168.450 96.560 168.710 ;
        RECT 109.640 168.450 109.900 168.710 ;
        RECT 85.260 167.770 85.520 168.030 ;
        RECT 85.720 167.770 85.980 168.030 ;
        RECT 86.180 167.770 86.440 168.030 ;
        RECT 92.620 167.770 92.880 168.030 ;
        RECT 96.760 167.770 97.020 168.030 ;
        RECT 99.060 167.770 99.320 168.030 ;
        RECT 73.695 167.260 73.955 167.520 ;
        RECT 74.015 167.260 74.275 167.520 ;
        RECT 74.335 167.260 74.595 167.520 ;
        RECT 74.655 167.260 74.915 167.520 ;
        RECT 74.975 167.260 75.235 167.520 ;
        RECT 87.265 167.260 87.525 167.520 ;
        RECT 87.585 167.260 87.845 167.520 ;
        RECT 87.905 167.260 88.165 167.520 ;
        RECT 88.225 167.260 88.485 167.520 ;
        RECT 88.545 167.260 88.805 167.520 ;
        RECT 100.835 167.260 101.095 167.520 ;
        RECT 101.155 167.260 101.415 167.520 ;
        RECT 101.475 167.260 101.735 167.520 ;
        RECT 101.795 167.260 102.055 167.520 ;
        RECT 102.115 167.260 102.375 167.520 ;
        RECT 114.405 167.260 114.665 167.520 ;
        RECT 114.725 167.260 114.985 167.520 ;
        RECT 115.045 167.260 115.305 167.520 ;
        RECT 115.365 167.260 115.625 167.520 ;
        RECT 115.685 167.260 115.945 167.520 ;
        RECT 83.420 166.410 83.680 166.670 ;
        RECT 87.560 166.070 87.820 166.330 ;
        RECT 85.260 165.730 85.520 165.990 ;
        RECT 86.180 165.730 86.440 165.990 ;
        RECT 99.980 166.750 100.240 167.010 ;
        RECT 89.400 166.070 89.660 166.330 ;
        RECT 65.020 165.390 65.280 165.650 ;
        RECT 89.860 165.730 90.120 165.990 ;
        RECT 85.720 165.050 85.980 165.310 ;
        RECT 95.840 165.050 96.100 165.310 ;
        RECT 99.520 165.050 99.780 165.310 ;
        RECT 80.480 164.540 80.740 164.800 ;
        RECT 80.800 164.540 81.060 164.800 ;
        RECT 81.120 164.540 81.380 164.800 ;
        RECT 81.440 164.540 81.700 164.800 ;
        RECT 81.760 164.540 82.020 164.800 ;
        RECT 94.050 164.540 94.310 164.800 ;
        RECT 94.370 164.540 94.630 164.800 ;
        RECT 94.690 164.540 94.950 164.800 ;
        RECT 95.010 164.540 95.270 164.800 ;
        RECT 95.330 164.540 95.590 164.800 ;
        RECT 107.620 164.540 107.880 164.800 ;
        RECT 107.940 164.540 108.200 164.800 ;
        RECT 108.260 164.540 108.520 164.800 ;
        RECT 108.580 164.540 108.840 164.800 ;
        RECT 108.900 164.540 109.160 164.800 ;
        RECT 121.190 164.540 121.450 164.800 ;
        RECT 121.510 164.540 121.770 164.800 ;
        RECT 121.830 164.540 122.090 164.800 ;
        RECT 122.150 164.540 122.410 164.800 ;
        RECT 122.470 164.540 122.730 164.800 ;
        RECT 83.880 164.030 84.140 164.290 ;
        RECT 89.860 164.030 90.120 164.290 ;
        RECT 99.520 163.690 99.780 163.950 ;
        RECT 85.720 163.350 85.980 163.610 ;
        RECT 92.620 163.010 92.880 163.270 ;
        RECT 95.840 163.350 96.100 163.610 ;
        RECT 103.200 163.010 103.460 163.270 ;
        RECT 109.180 163.010 109.440 163.270 ;
        RECT 99.060 162.330 99.320 162.590 ;
        RECT 103.660 162.330 103.920 162.590 ;
        RECT 73.695 161.820 73.955 162.080 ;
        RECT 74.015 161.820 74.275 162.080 ;
        RECT 74.335 161.820 74.595 162.080 ;
        RECT 74.655 161.820 74.915 162.080 ;
        RECT 74.975 161.820 75.235 162.080 ;
        RECT 87.265 161.820 87.525 162.080 ;
        RECT 87.585 161.820 87.845 162.080 ;
        RECT 87.905 161.820 88.165 162.080 ;
        RECT 88.225 161.820 88.485 162.080 ;
        RECT 88.545 161.820 88.805 162.080 ;
        RECT 100.835 161.820 101.095 162.080 ;
        RECT 101.155 161.820 101.415 162.080 ;
        RECT 101.475 161.820 101.735 162.080 ;
        RECT 101.795 161.820 102.055 162.080 ;
        RECT 102.115 161.820 102.375 162.080 ;
        RECT 114.405 161.820 114.665 162.080 ;
        RECT 114.725 161.820 114.985 162.080 ;
        RECT 115.045 161.820 115.305 162.080 ;
        RECT 115.365 161.820 115.625 162.080 ;
        RECT 115.685 161.820 115.945 162.080 ;
        RECT 83.420 161.310 83.680 161.570 ;
        RECT 103.200 161.310 103.460 161.570 ;
        RECT 109.180 161.310 109.440 161.570 ;
        RECT 99.520 160.290 99.780 160.550 ;
        RECT 103.660 160.290 103.920 160.550 ;
        RECT 100.440 159.950 100.700 160.210 ;
        RECT 80.480 159.100 80.740 159.360 ;
        RECT 80.800 159.100 81.060 159.360 ;
        RECT 81.120 159.100 81.380 159.360 ;
        RECT 81.440 159.100 81.700 159.360 ;
        RECT 81.760 159.100 82.020 159.360 ;
        RECT 94.050 159.100 94.310 159.360 ;
        RECT 94.370 159.100 94.630 159.360 ;
        RECT 94.690 159.100 94.950 159.360 ;
        RECT 95.010 159.100 95.270 159.360 ;
        RECT 95.330 159.100 95.590 159.360 ;
        RECT 107.620 159.100 107.880 159.360 ;
        RECT 107.940 159.100 108.200 159.360 ;
        RECT 108.260 159.100 108.520 159.360 ;
        RECT 108.580 159.100 108.840 159.360 ;
        RECT 108.900 159.100 109.160 159.360 ;
        RECT 121.190 159.100 121.450 159.360 ;
        RECT 121.510 159.100 121.770 159.360 ;
        RECT 121.830 159.100 122.090 159.360 ;
        RECT 122.150 159.100 122.410 159.360 ;
        RECT 122.470 159.100 122.730 159.360 ;
        RECT 85.740 102.970 86.180 103.390 ;
        RECT 89.410 102.890 89.980 103.450 ;
        RECT 92.810 102.880 93.380 103.440 ;
        RECT 81.830 90.650 83.010 91.800 ;
        RECT 96.570 102.910 97.140 103.470 ;
        RECT 105.360 72.810 105.810 73.210 ;
      LAYER met2 ;
        RECT 84.330 214.510 84.610 216.510 ;
        RECT 122.970 214.510 123.250 216.510 ;
        RECT 80.480 213.445 82.020 213.815 ;
        RECT 73.695 210.725 75.235 211.095 ;
        RECT 80.480 208.005 82.020 208.375 ;
        RECT 73.695 205.285 75.235 205.655 ;
        RECT 80.480 202.565 82.020 202.935 ;
        RECT 73.695 199.845 75.235 200.215 ;
        RECT 78.810 197.465 79.090 197.835 ;
        RECT 73.695 194.405 75.235 194.775 ;
        RECT 78.880 194.240 79.020 197.465 ;
        RECT 80.480 197.125 82.020 197.495 ;
        RECT 78.820 193.920 79.080 194.240 ;
        RECT 80.480 191.685 82.020 192.055 ;
        RECT 84.400 191.080 84.540 214.510 ;
        RECT 94.050 213.445 95.590 213.815 ;
        RECT 107.620 213.445 109.160 213.815 ;
        RECT 121.190 213.445 122.730 213.815 ;
        RECT 87.265 210.725 88.805 211.095 ;
        RECT 100.835 210.725 102.375 211.095 ;
        RECT 114.405 210.725 115.945 211.095 ;
        RECT 94.050 208.005 95.590 208.375 ;
        RECT 107.620 208.005 109.160 208.375 ;
        RECT 121.190 208.005 122.730 208.375 ;
        RECT 87.265 205.285 88.805 205.655 ;
        RECT 100.835 205.285 102.375 205.655 ;
        RECT 114.405 205.285 115.945 205.655 ;
        RECT 94.050 202.565 95.590 202.935 ;
        RECT 107.620 202.565 109.160 202.935 ;
        RECT 121.190 202.565 122.730 202.935 ;
        RECT 87.265 199.845 88.805 200.215 ;
        RECT 100.835 199.845 102.375 200.215 ;
        RECT 114.405 199.845 115.945 200.215 ;
        RECT 94.050 197.125 95.590 197.495 ;
        RECT 107.620 197.125 109.160 197.495 ;
        RECT 121.190 197.125 122.730 197.495 ;
        RECT 87.265 194.405 88.805 194.775 ;
        RECT 100.835 194.405 102.375 194.775 ;
        RECT 114.405 194.405 115.945 194.775 ;
        RECT 92.620 193.920 92.880 194.240 ;
        RECT 84.400 190.940 85.000 191.080 ;
        RECT 73.695 188.965 75.235 189.335 ;
        RECT 80.480 186.245 82.020 186.615 ;
        RECT 73.695 183.525 75.235 183.895 ;
        RECT 80.480 180.805 82.020 181.175 ;
        RECT 73.695 178.085 75.235 178.455 ;
        RECT 80.480 175.365 82.020 175.735 ;
        RECT 73.695 172.645 75.235 173.015 ;
        RECT 83.420 170.460 83.680 170.780 ;
        RECT 80.480 169.925 82.020 170.295 ;
        RECT 73.695 167.205 75.235 167.575 ;
        RECT 83.480 166.700 83.620 170.460 ;
        RECT 84.860 170.380 85.000 190.940 ;
        RECT 87.265 188.965 88.805 189.335 ;
        RECT 87.265 183.525 88.805 183.895 ;
        RECT 87.265 178.085 88.805 178.455 ;
        RECT 87.265 172.645 88.805 173.015 ;
        RECT 92.680 171.460 92.820 193.920 ;
        RECT 94.050 191.685 95.590 192.055 ;
        RECT 107.620 191.685 109.160 192.055 ;
        RECT 121.190 191.685 122.730 192.055 ;
        RECT 100.835 188.965 102.375 189.335 ;
        RECT 114.405 188.965 115.945 189.335 ;
        RECT 94.050 186.245 95.590 186.615 ;
        RECT 107.620 186.245 109.160 186.615 ;
        RECT 121.190 186.245 122.730 186.615 ;
        RECT 100.835 183.525 102.375 183.895 ;
        RECT 114.405 183.525 115.945 183.895 ;
        RECT 94.050 180.805 95.590 181.175 ;
        RECT 107.620 180.805 109.160 181.175 ;
        RECT 121.190 180.805 122.730 181.175 ;
        RECT 100.835 178.085 102.375 178.455 ;
        RECT 114.405 178.085 115.945 178.455 ;
        RECT 123.040 177.240 123.180 214.510 ;
        RECT 99.060 176.920 99.320 177.240 ;
        RECT 122.980 176.920 123.240 177.240 ;
        RECT 94.050 175.365 95.590 175.735 ;
        RECT 99.120 175.200 99.260 176.920 ;
        RECT 107.620 175.365 109.160 175.735 ;
        RECT 121.190 175.365 122.730 175.735 ;
        RECT 99.060 174.880 99.320 175.200 ;
        RECT 96.300 174.540 96.560 174.860 ;
        RECT 93.540 173.860 93.800 174.180 ;
        RECT 93.080 173.180 93.340 173.500 ;
        RECT 86.640 171.140 86.900 171.460 ;
        RECT 92.620 171.140 92.880 171.460 ;
        RECT 84.860 170.240 85.460 170.380 ;
        RECT 85.320 169.275 85.460 170.240 ;
        RECT 85.250 168.905 85.530 169.275 ;
        RECT 85.260 168.760 85.520 168.905 ;
        RECT 83.880 168.420 84.140 168.740 ;
        RECT 83.420 166.380 83.680 166.700 ;
        RECT 65.020 165.360 65.280 165.680 ;
        RECT 65.080 158.510 65.220 165.360 ;
        RECT 80.480 164.485 82.020 164.855 ;
        RECT 73.695 161.765 75.235 162.135 ;
        RECT 83.480 161.600 83.620 166.380 ;
        RECT 83.940 164.320 84.080 168.420 ;
        RECT 85.260 167.740 85.520 168.060 ;
        RECT 85.720 167.740 85.980 168.060 ;
        RECT 86.180 167.740 86.440 168.060 ;
        RECT 85.320 166.020 85.460 167.740 ;
        RECT 85.260 165.700 85.520 166.020 ;
        RECT 85.780 165.340 85.920 167.740 ;
        RECT 86.240 166.020 86.380 167.740 ;
        RECT 86.700 166.440 86.840 171.140 ;
        RECT 92.620 170.460 92.880 170.780 ;
        RECT 92.680 169.275 92.820 170.460 ;
        RECT 93.140 169.760 93.280 173.180 ;
        RECT 93.600 170.780 93.740 173.860 ;
        RECT 95.840 171.140 96.100 171.460 ;
        RECT 93.540 170.460 93.800 170.780 ;
        RECT 94.050 169.925 95.590 170.295 ;
        RECT 93.080 169.440 93.340 169.760 ;
        RECT 89.400 168.760 89.660 169.080 ;
        RECT 92.610 168.905 92.890 169.275 ;
        RECT 95.900 169.080 96.040 171.140 ;
        RECT 92.620 168.760 92.880 168.905 ;
        RECT 95.840 168.760 96.100 169.080 ;
        RECT 87.265 167.205 88.805 167.575 ;
        RECT 86.700 166.360 87.760 166.440 ;
        RECT 89.460 166.360 89.600 168.760 ;
        RECT 96.360 168.740 96.500 174.540 ;
        RECT 96.760 173.180 97.020 173.500 ;
        RECT 96.300 168.420 96.560 168.740 ;
        RECT 92.620 167.740 92.880 168.060 ;
        RECT 96.360 167.800 96.500 168.420 ;
        RECT 96.820 168.060 96.960 173.180 ;
        RECT 98.600 170.460 98.860 170.780 ;
        RECT 98.660 169.760 98.800 170.460 ;
        RECT 98.600 169.440 98.860 169.760 ;
        RECT 99.120 169.160 99.260 174.880 ;
        RECT 105.500 173.860 105.760 174.180 ;
        RECT 109.640 173.860 109.900 174.180 ;
        RECT 121.140 174.035 121.400 174.180 ;
        RECT 100.835 172.645 102.375 173.015 ;
        RECT 105.560 172.480 105.700 173.860 ;
        RECT 105.500 172.160 105.760 172.480 ;
        RECT 100.440 170.460 100.700 170.780 ;
        RECT 106.420 170.460 106.680 170.780 ;
        RECT 106.880 170.460 107.140 170.780 ;
        RECT 98.200 169.080 99.260 169.160 ;
        RECT 99.980 169.100 100.240 169.420 ;
        RECT 98.140 169.020 99.260 169.080 ;
        RECT 98.140 168.760 98.400 169.020 ;
        RECT 86.700 166.300 87.820 166.360 ;
        RECT 87.560 166.040 87.820 166.300 ;
        RECT 89.400 166.040 89.660 166.360 ;
        RECT 86.180 165.700 86.440 166.020 ;
        RECT 89.860 165.700 90.120 166.020 ;
        RECT 85.720 165.020 85.980 165.340 ;
        RECT 83.880 164.000 84.140 164.320 ;
        RECT 85.780 163.640 85.920 165.020 ;
        RECT 89.920 164.320 90.060 165.700 ;
        RECT 89.860 164.000 90.120 164.320 ;
        RECT 85.720 163.320 85.980 163.640 ;
        RECT 92.680 163.300 92.820 167.740 ;
        RECT 95.900 167.660 96.500 167.800 ;
        RECT 96.760 167.740 97.020 168.060 ;
        RECT 99.060 167.740 99.320 168.060 ;
        RECT 95.900 165.340 96.040 167.660 ;
        RECT 95.840 165.020 96.100 165.340 ;
        RECT 94.050 164.485 95.590 164.855 ;
        RECT 95.900 163.640 96.040 165.020 ;
        RECT 95.840 163.320 96.100 163.640 ;
        RECT 92.620 162.980 92.880 163.300 ;
        RECT 99.120 162.620 99.260 167.740 ;
        RECT 100.040 167.040 100.180 169.100 ;
        RECT 99.980 166.720 100.240 167.040 ;
        RECT 99.520 165.020 99.780 165.340 ;
        RECT 99.580 163.980 99.720 165.020 ;
        RECT 99.520 163.660 99.780 163.980 ;
        RECT 99.060 162.300 99.320 162.620 ;
        RECT 87.265 161.765 88.805 162.135 ;
        RECT 83.420 161.280 83.680 161.600 ;
        RECT 99.580 160.580 99.720 163.660 ;
        RECT 99.520 160.260 99.780 160.580 ;
        RECT 100.500 160.240 100.640 170.460 ;
        RECT 106.480 169.420 106.620 170.460 ;
        RECT 106.940 169.760 107.080 170.460 ;
        RECT 107.620 169.925 109.160 170.295 ;
        RECT 106.880 169.440 107.140 169.760 ;
        RECT 106.420 169.100 106.680 169.420 ;
        RECT 109.700 168.740 109.840 173.860 ;
        RECT 121.130 173.665 121.410 174.035 ;
        RECT 117.920 173.180 118.180 173.500 ;
        RECT 114.405 172.645 115.945 173.015 ;
        RECT 117.980 172.480 118.120 173.180 ;
        RECT 117.920 172.160 118.180 172.480 ;
        RECT 121.190 169.925 122.730 170.295 ;
        RECT 109.640 168.420 109.900 168.740 ;
        RECT 100.835 167.205 102.375 167.575 ;
        RECT 107.620 164.485 109.160 164.855 ;
        RECT 109.700 163.720 109.840 168.420 ;
        RECT 114.405 167.205 115.945 167.575 ;
        RECT 121.190 164.485 122.730 164.855 ;
        RECT 109.240 163.580 109.840 163.720 ;
        RECT 109.240 163.300 109.380 163.580 ;
        RECT 103.200 162.980 103.460 163.300 ;
        RECT 109.180 162.980 109.440 163.300 ;
        RECT 100.835 161.765 102.375 162.135 ;
        RECT 103.260 161.600 103.400 162.980 ;
        RECT 103.660 162.300 103.920 162.620 ;
        RECT 103.200 161.280 103.460 161.600 ;
        RECT 103.720 160.580 103.860 162.300 ;
        RECT 109.240 161.600 109.380 162.980 ;
        RECT 114.405 161.765 115.945 162.135 ;
        RECT 109.180 161.280 109.440 161.600 ;
        RECT 103.660 160.260 103.920 160.580 ;
        RECT 100.440 159.920 100.700 160.240 ;
        RECT 80.480 159.045 82.020 159.415 ;
        RECT 94.050 159.045 95.590 159.415 ;
        RECT 103.720 158.510 103.860 160.260 ;
        RECT 107.620 159.045 109.160 159.415 ;
        RECT 121.190 159.045 122.730 159.415 ;
        RECT 65.010 156.510 65.290 158.510 ;
        RECT 103.650 156.510 103.930 158.510 ;
        RECT 85.740 102.920 86.180 103.440 ;
        RECT 89.410 102.840 89.980 103.500 ;
        RECT 92.810 102.830 93.380 103.490 ;
        RECT 96.570 102.860 97.140 103.520 ;
        RECT 81.830 90.600 83.010 91.850 ;
        RECT 105.360 72.760 105.810 73.260 ;
      LAYER via2 ;
        RECT 80.510 213.490 80.790 213.770 ;
        RECT 80.910 213.490 81.190 213.770 ;
        RECT 81.310 213.490 81.590 213.770 ;
        RECT 81.710 213.490 81.990 213.770 ;
        RECT 73.725 210.770 74.005 211.050 ;
        RECT 74.125 210.770 74.405 211.050 ;
        RECT 74.525 210.770 74.805 211.050 ;
        RECT 74.925 210.770 75.205 211.050 ;
        RECT 80.510 208.050 80.790 208.330 ;
        RECT 80.910 208.050 81.190 208.330 ;
        RECT 81.310 208.050 81.590 208.330 ;
        RECT 81.710 208.050 81.990 208.330 ;
        RECT 73.725 205.330 74.005 205.610 ;
        RECT 74.125 205.330 74.405 205.610 ;
        RECT 74.525 205.330 74.805 205.610 ;
        RECT 74.925 205.330 75.205 205.610 ;
        RECT 80.510 202.610 80.790 202.890 ;
        RECT 80.910 202.610 81.190 202.890 ;
        RECT 81.310 202.610 81.590 202.890 ;
        RECT 81.710 202.610 81.990 202.890 ;
        RECT 73.725 199.890 74.005 200.170 ;
        RECT 74.125 199.890 74.405 200.170 ;
        RECT 74.525 199.890 74.805 200.170 ;
        RECT 74.925 199.890 75.205 200.170 ;
        RECT 78.810 197.510 79.090 197.790 ;
        RECT 73.725 194.450 74.005 194.730 ;
        RECT 74.125 194.450 74.405 194.730 ;
        RECT 74.525 194.450 74.805 194.730 ;
        RECT 74.925 194.450 75.205 194.730 ;
        RECT 80.510 197.170 80.790 197.450 ;
        RECT 80.910 197.170 81.190 197.450 ;
        RECT 81.310 197.170 81.590 197.450 ;
        RECT 81.710 197.170 81.990 197.450 ;
        RECT 80.510 191.730 80.790 192.010 ;
        RECT 80.910 191.730 81.190 192.010 ;
        RECT 81.310 191.730 81.590 192.010 ;
        RECT 81.710 191.730 81.990 192.010 ;
        RECT 94.080 213.490 94.360 213.770 ;
        RECT 94.480 213.490 94.760 213.770 ;
        RECT 94.880 213.490 95.160 213.770 ;
        RECT 95.280 213.490 95.560 213.770 ;
        RECT 107.650 213.490 107.930 213.770 ;
        RECT 108.050 213.490 108.330 213.770 ;
        RECT 108.450 213.490 108.730 213.770 ;
        RECT 108.850 213.490 109.130 213.770 ;
        RECT 121.220 213.490 121.500 213.770 ;
        RECT 121.620 213.490 121.900 213.770 ;
        RECT 122.020 213.490 122.300 213.770 ;
        RECT 122.420 213.490 122.700 213.770 ;
        RECT 87.295 210.770 87.575 211.050 ;
        RECT 87.695 210.770 87.975 211.050 ;
        RECT 88.095 210.770 88.375 211.050 ;
        RECT 88.495 210.770 88.775 211.050 ;
        RECT 100.865 210.770 101.145 211.050 ;
        RECT 101.265 210.770 101.545 211.050 ;
        RECT 101.665 210.770 101.945 211.050 ;
        RECT 102.065 210.770 102.345 211.050 ;
        RECT 114.435 210.770 114.715 211.050 ;
        RECT 114.835 210.770 115.115 211.050 ;
        RECT 115.235 210.770 115.515 211.050 ;
        RECT 115.635 210.770 115.915 211.050 ;
        RECT 94.080 208.050 94.360 208.330 ;
        RECT 94.480 208.050 94.760 208.330 ;
        RECT 94.880 208.050 95.160 208.330 ;
        RECT 95.280 208.050 95.560 208.330 ;
        RECT 107.650 208.050 107.930 208.330 ;
        RECT 108.050 208.050 108.330 208.330 ;
        RECT 108.450 208.050 108.730 208.330 ;
        RECT 108.850 208.050 109.130 208.330 ;
        RECT 121.220 208.050 121.500 208.330 ;
        RECT 121.620 208.050 121.900 208.330 ;
        RECT 122.020 208.050 122.300 208.330 ;
        RECT 122.420 208.050 122.700 208.330 ;
        RECT 87.295 205.330 87.575 205.610 ;
        RECT 87.695 205.330 87.975 205.610 ;
        RECT 88.095 205.330 88.375 205.610 ;
        RECT 88.495 205.330 88.775 205.610 ;
        RECT 100.865 205.330 101.145 205.610 ;
        RECT 101.265 205.330 101.545 205.610 ;
        RECT 101.665 205.330 101.945 205.610 ;
        RECT 102.065 205.330 102.345 205.610 ;
        RECT 114.435 205.330 114.715 205.610 ;
        RECT 114.835 205.330 115.115 205.610 ;
        RECT 115.235 205.330 115.515 205.610 ;
        RECT 115.635 205.330 115.915 205.610 ;
        RECT 94.080 202.610 94.360 202.890 ;
        RECT 94.480 202.610 94.760 202.890 ;
        RECT 94.880 202.610 95.160 202.890 ;
        RECT 95.280 202.610 95.560 202.890 ;
        RECT 107.650 202.610 107.930 202.890 ;
        RECT 108.050 202.610 108.330 202.890 ;
        RECT 108.450 202.610 108.730 202.890 ;
        RECT 108.850 202.610 109.130 202.890 ;
        RECT 121.220 202.610 121.500 202.890 ;
        RECT 121.620 202.610 121.900 202.890 ;
        RECT 122.020 202.610 122.300 202.890 ;
        RECT 122.420 202.610 122.700 202.890 ;
        RECT 87.295 199.890 87.575 200.170 ;
        RECT 87.695 199.890 87.975 200.170 ;
        RECT 88.095 199.890 88.375 200.170 ;
        RECT 88.495 199.890 88.775 200.170 ;
        RECT 100.865 199.890 101.145 200.170 ;
        RECT 101.265 199.890 101.545 200.170 ;
        RECT 101.665 199.890 101.945 200.170 ;
        RECT 102.065 199.890 102.345 200.170 ;
        RECT 114.435 199.890 114.715 200.170 ;
        RECT 114.835 199.890 115.115 200.170 ;
        RECT 115.235 199.890 115.515 200.170 ;
        RECT 115.635 199.890 115.915 200.170 ;
        RECT 94.080 197.170 94.360 197.450 ;
        RECT 94.480 197.170 94.760 197.450 ;
        RECT 94.880 197.170 95.160 197.450 ;
        RECT 95.280 197.170 95.560 197.450 ;
        RECT 107.650 197.170 107.930 197.450 ;
        RECT 108.050 197.170 108.330 197.450 ;
        RECT 108.450 197.170 108.730 197.450 ;
        RECT 108.850 197.170 109.130 197.450 ;
        RECT 121.220 197.170 121.500 197.450 ;
        RECT 121.620 197.170 121.900 197.450 ;
        RECT 122.020 197.170 122.300 197.450 ;
        RECT 122.420 197.170 122.700 197.450 ;
        RECT 87.295 194.450 87.575 194.730 ;
        RECT 87.695 194.450 87.975 194.730 ;
        RECT 88.095 194.450 88.375 194.730 ;
        RECT 88.495 194.450 88.775 194.730 ;
        RECT 100.865 194.450 101.145 194.730 ;
        RECT 101.265 194.450 101.545 194.730 ;
        RECT 101.665 194.450 101.945 194.730 ;
        RECT 102.065 194.450 102.345 194.730 ;
        RECT 114.435 194.450 114.715 194.730 ;
        RECT 114.835 194.450 115.115 194.730 ;
        RECT 115.235 194.450 115.515 194.730 ;
        RECT 115.635 194.450 115.915 194.730 ;
        RECT 73.725 189.010 74.005 189.290 ;
        RECT 74.125 189.010 74.405 189.290 ;
        RECT 74.525 189.010 74.805 189.290 ;
        RECT 74.925 189.010 75.205 189.290 ;
        RECT 80.510 186.290 80.790 186.570 ;
        RECT 80.910 186.290 81.190 186.570 ;
        RECT 81.310 186.290 81.590 186.570 ;
        RECT 81.710 186.290 81.990 186.570 ;
        RECT 73.725 183.570 74.005 183.850 ;
        RECT 74.125 183.570 74.405 183.850 ;
        RECT 74.525 183.570 74.805 183.850 ;
        RECT 74.925 183.570 75.205 183.850 ;
        RECT 80.510 180.850 80.790 181.130 ;
        RECT 80.910 180.850 81.190 181.130 ;
        RECT 81.310 180.850 81.590 181.130 ;
        RECT 81.710 180.850 81.990 181.130 ;
        RECT 73.725 178.130 74.005 178.410 ;
        RECT 74.125 178.130 74.405 178.410 ;
        RECT 74.525 178.130 74.805 178.410 ;
        RECT 74.925 178.130 75.205 178.410 ;
        RECT 80.510 175.410 80.790 175.690 ;
        RECT 80.910 175.410 81.190 175.690 ;
        RECT 81.310 175.410 81.590 175.690 ;
        RECT 81.710 175.410 81.990 175.690 ;
        RECT 73.725 172.690 74.005 172.970 ;
        RECT 74.125 172.690 74.405 172.970 ;
        RECT 74.525 172.690 74.805 172.970 ;
        RECT 74.925 172.690 75.205 172.970 ;
        RECT 80.510 169.970 80.790 170.250 ;
        RECT 80.910 169.970 81.190 170.250 ;
        RECT 81.310 169.970 81.590 170.250 ;
        RECT 81.710 169.970 81.990 170.250 ;
        RECT 73.725 167.250 74.005 167.530 ;
        RECT 74.125 167.250 74.405 167.530 ;
        RECT 74.525 167.250 74.805 167.530 ;
        RECT 74.925 167.250 75.205 167.530 ;
        RECT 87.295 189.010 87.575 189.290 ;
        RECT 87.695 189.010 87.975 189.290 ;
        RECT 88.095 189.010 88.375 189.290 ;
        RECT 88.495 189.010 88.775 189.290 ;
        RECT 87.295 183.570 87.575 183.850 ;
        RECT 87.695 183.570 87.975 183.850 ;
        RECT 88.095 183.570 88.375 183.850 ;
        RECT 88.495 183.570 88.775 183.850 ;
        RECT 87.295 178.130 87.575 178.410 ;
        RECT 87.695 178.130 87.975 178.410 ;
        RECT 88.095 178.130 88.375 178.410 ;
        RECT 88.495 178.130 88.775 178.410 ;
        RECT 87.295 172.690 87.575 172.970 ;
        RECT 87.695 172.690 87.975 172.970 ;
        RECT 88.095 172.690 88.375 172.970 ;
        RECT 88.495 172.690 88.775 172.970 ;
        RECT 94.080 191.730 94.360 192.010 ;
        RECT 94.480 191.730 94.760 192.010 ;
        RECT 94.880 191.730 95.160 192.010 ;
        RECT 95.280 191.730 95.560 192.010 ;
        RECT 107.650 191.730 107.930 192.010 ;
        RECT 108.050 191.730 108.330 192.010 ;
        RECT 108.450 191.730 108.730 192.010 ;
        RECT 108.850 191.730 109.130 192.010 ;
        RECT 121.220 191.730 121.500 192.010 ;
        RECT 121.620 191.730 121.900 192.010 ;
        RECT 122.020 191.730 122.300 192.010 ;
        RECT 122.420 191.730 122.700 192.010 ;
        RECT 100.865 189.010 101.145 189.290 ;
        RECT 101.265 189.010 101.545 189.290 ;
        RECT 101.665 189.010 101.945 189.290 ;
        RECT 102.065 189.010 102.345 189.290 ;
        RECT 114.435 189.010 114.715 189.290 ;
        RECT 114.835 189.010 115.115 189.290 ;
        RECT 115.235 189.010 115.515 189.290 ;
        RECT 115.635 189.010 115.915 189.290 ;
        RECT 94.080 186.290 94.360 186.570 ;
        RECT 94.480 186.290 94.760 186.570 ;
        RECT 94.880 186.290 95.160 186.570 ;
        RECT 95.280 186.290 95.560 186.570 ;
        RECT 107.650 186.290 107.930 186.570 ;
        RECT 108.050 186.290 108.330 186.570 ;
        RECT 108.450 186.290 108.730 186.570 ;
        RECT 108.850 186.290 109.130 186.570 ;
        RECT 121.220 186.290 121.500 186.570 ;
        RECT 121.620 186.290 121.900 186.570 ;
        RECT 122.020 186.290 122.300 186.570 ;
        RECT 122.420 186.290 122.700 186.570 ;
        RECT 100.865 183.570 101.145 183.850 ;
        RECT 101.265 183.570 101.545 183.850 ;
        RECT 101.665 183.570 101.945 183.850 ;
        RECT 102.065 183.570 102.345 183.850 ;
        RECT 114.435 183.570 114.715 183.850 ;
        RECT 114.835 183.570 115.115 183.850 ;
        RECT 115.235 183.570 115.515 183.850 ;
        RECT 115.635 183.570 115.915 183.850 ;
        RECT 94.080 180.850 94.360 181.130 ;
        RECT 94.480 180.850 94.760 181.130 ;
        RECT 94.880 180.850 95.160 181.130 ;
        RECT 95.280 180.850 95.560 181.130 ;
        RECT 107.650 180.850 107.930 181.130 ;
        RECT 108.050 180.850 108.330 181.130 ;
        RECT 108.450 180.850 108.730 181.130 ;
        RECT 108.850 180.850 109.130 181.130 ;
        RECT 121.220 180.850 121.500 181.130 ;
        RECT 121.620 180.850 121.900 181.130 ;
        RECT 122.020 180.850 122.300 181.130 ;
        RECT 122.420 180.850 122.700 181.130 ;
        RECT 100.865 178.130 101.145 178.410 ;
        RECT 101.265 178.130 101.545 178.410 ;
        RECT 101.665 178.130 101.945 178.410 ;
        RECT 102.065 178.130 102.345 178.410 ;
        RECT 114.435 178.130 114.715 178.410 ;
        RECT 114.835 178.130 115.115 178.410 ;
        RECT 115.235 178.130 115.515 178.410 ;
        RECT 115.635 178.130 115.915 178.410 ;
        RECT 94.080 175.410 94.360 175.690 ;
        RECT 94.480 175.410 94.760 175.690 ;
        RECT 94.880 175.410 95.160 175.690 ;
        RECT 95.280 175.410 95.560 175.690 ;
        RECT 107.650 175.410 107.930 175.690 ;
        RECT 108.050 175.410 108.330 175.690 ;
        RECT 108.450 175.410 108.730 175.690 ;
        RECT 108.850 175.410 109.130 175.690 ;
        RECT 121.220 175.410 121.500 175.690 ;
        RECT 121.620 175.410 121.900 175.690 ;
        RECT 122.020 175.410 122.300 175.690 ;
        RECT 122.420 175.410 122.700 175.690 ;
        RECT 85.250 168.950 85.530 169.230 ;
        RECT 80.510 164.530 80.790 164.810 ;
        RECT 80.910 164.530 81.190 164.810 ;
        RECT 81.310 164.530 81.590 164.810 ;
        RECT 81.710 164.530 81.990 164.810 ;
        RECT 73.725 161.810 74.005 162.090 ;
        RECT 74.125 161.810 74.405 162.090 ;
        RECT 74.525 161.810 74.805 162.090 ;
        RECT 74.925 161.810 75.205 162.090 ;
        RECT 94.080 169.970 94.360 170.250 ;
        RECT 94.480 169.970 94.760 170.250 ;
        RECT 94.880 169.970 95.160 170.250 ;
        RECT 95.280 169.970 95.560 170.250 ;
        RECT 92.610 168.950 92.890 169.230 ;
        RECT 87.295 167.250 87.575 167.530 ;
        RECT 87.695 167.250 87.975 167.530 ;
        RECT 88.095 167.250 88.375 167.530 ;
        RECT 88.495 167.250 88.775 167.530 ;
        RECT 100.865 172.690 101.145 172.970 ;
        RECT 101.265 172.690 101.545 172.970 ;
        RECT 101.665 172.690 101.945 172.970 ;
        RECT 102.065 172.690 102.345 172.970 ;
        RECT 94.080 164.530 94.360 164.810 ;
        RECT 94.480 164.530 94.760 164.810 ;
        RECT 94.880 164.530 95.160 164.810 ;
        RECT 95.280 164.530 95.560 164.810 ;
        RECT 87.295 161.810 87.575 162.090 ;
        RECT 87.695 161.810 87.975 162.090 ;
        RECT 88.095 161.810 88.375 162.090 ;
        RECT 88.495 161.810 88.775 162.090 ;
        RECT 107.650 169.970 107.930 170.250 ;
        RECT 108.050 169.970 108.330 170.250 ;
        RECT 108.450 169.970 108.730 170.250 ;
        RECT 108.850 169.970 109.130 170.250 ;
        RECT 121.130 173.710 121.410 173.990 ;
        RECT 114.435 172.690 114.715 172.970 ;
        RECT 114.835 172.690 115.115 172.970 ;
        RECT 115.235 172.690 115.515 172.970 ;
        RECT 115.635 172.690 115.915 172.970 ;
        RECT 121.220 169.970 121.500 170.250 ;
        RECT 121.620 169.970 121.900 170.250 ;
        RECT 122.020 169.970 122.300 170.250 ;
        RECT 122.420 169.970 122.700 170.250 ;
        RECT 100.865 167.250 101.145 167.530 ;
        RECT 101.265 167.250 101.545 167.530 ;
        RECT 101.665 167.250 101.945 167.530 ;
        RECT 102.065 167.250 102.345 167.530 ;
        RECT 107.650 164.530 107.930 164.810 ;
        RECT 108.050 164.530 108.330 164.810 ;
        RECT 108.450 164.530 108.730 164.810 ;
        RECT 108.850 164.530 109.130 164.810 ;
        RECT 114.435 167.250 114.715 167.530 ;
        RECT 114.835 167.250 115.115 167.530 ;
        RECT 115.235 167.250 115.515 167.530 ;
        RECT 115.635 167.250 115.915 167.530 ;
        RECT 121.220 164.530 121.500 164.810 ;
        RECT 121.620 164.530 121.900 164.810 ;
        RECT 122.020 164.530 122.300 164.810 ;
        RECT 122.420 164.530 122.700 164.810 ;
        RECT 100.865 161.810 101.145 162.090 ;
        RECT 101.265 161.810 101.545 162.090 ;
        RECT 101.665 161.810 101.945 162.090 ;
        RECT 102.065 161.810 102.345 162.090 ;
        RECT 114.435 161.810 114.715 162.090 ;
        RECT 114.835 161.810 115.115 162.090 ;
        RECT 115.235 161.810 115.515 162.090 ;
        RECT 115.635 161.810 115.915 162.090 ;
        RECT 80.510 159.090 80.790 159.370 ;
        RECT 80.910 159.090 81.190 159.370 ;
        RECT 81.310 159.090 81.590 159.370 ;
        RECT 81.710 159.090 81.990 159.370 ;
        RECT 94.080 159.090 94.360 159.370 ;
        RECT 94.480 159.090 94.760 159.370 ;
        RECT 94.880 159.090 95.160 159.370 ;
        RECT 95.280 159.090 95.560 159.370 ;
        RECT 107.650 159.090 107.930 159.370 ;
        RECT 108.050 159.090 108.330 159.370 ;
        RECT 108.450 159.090 108.730 159.370 ;
        RECT 108.850 159.090 109.130 159.370 ;
        RECT 121.220 159.090 121.500 159.370 ;
        RECT 121.620 159.090 121.900 159.370 ;
        RECT 122.020 159.090 122.300 159.370 ;
        RECT 122.420 159.090 122.700 159.370 ;
        RECT 85.740 102.970 86.180 103.390 ;
        RECT 89.410 102.890 89.980 103.450 ;
        RECT 92.810 102.880 93.380 103.440 ;
        RECT 96.570 102.910 97.140 103.470 ;
        RECT 81.830 90.650 83.010 91.800 ;
        RECT 105.360 72.810 105.810 73.210 ;
      LAYER met3 ;
        RECT 131.910 221.660 155.310 222.260 ;
        RECT 131.910 221.170 132.510 221.660 ;
        RECT 59.990 220.570 132.510 221.170 ;
        RECT 59.990 197.950 60.590 220.570 ;
        RECT 151.100 220.110 151.725 220.140 ;
        RECT 151.100 219.485 153.715 220.110 ;
        RECT 151.100 219.455 151.725 219.485 ;
        RECT 80.460 213.465 82.040 213.795 ;
        RECT 94.030 213.465 95.610 213.795 ;
        RECT 107.600 213.465 109.180 213.795 ;
        RECT 121.170 213.465 122.750 213.795 ;
        RECT 73.675 210.745 75.255 211.075 ;
        RECT 87.245 210.745 88.825 211.075 ;
        RECT 100.815 210.745 102.395 211.075 ;
        RECT 114.385 210.745 115.965 211.075 ;
        RECT 80.460 208.025 82.040 208.355 ;
        RECT 94.030 208.025 95.610 208.355 ;
        RECT 107.600 208.025 109.180 208.355 ;
        RECT 121.170 208.025 122.750 208.355 ;
        RECT 73.675 205.305 75.255 205.635 ;
        RECT 87.245 205.305 88.825 205.635 ;
        RECT 100.815 205.305 102.395 205.635 ;
        RECT 114.385 205.305 115.965 205.635 ;
        RECT 80.460 202.585 82.040 202.915 ;
        RECT 94.030 202.585 95.610 202.915 ;
        RECT 107.600 202.585 109.180 202.915 ;
        RECT 121.170 202.585 122.750 202.915 ;
        RECT 73.675 199.865 75.255 200.195 ;
        RECT 87.245 199.865 88.825 200.195 ;
        RECT 100.815 199.865 102.395 200.195 ;
        RECT 114.385 199.865 115.965 200.195 ;
        RECT 59.990 197.800 66.920 197.950 ;
        RECT 78.785 197.800 79.115 197.815 ;
        RECT 59.990 197.500 79.115 197.800 ;
        RECT 59.990 197.350 66.920 197.500 ;
        RECT 78.785 197.485 79.115 197.500 ;
        RECT 80.460 197.145 82.040 197.475 ;
        RECT 94.030 197.145 95.610 197.475 ;
        RECT 107.600 197.145 109.180 197.475 ;
        RECT 121.170 197.145 122.750 197.475 ;
        RECT 73.675 194.425 75.255 194.755 ;
        RECT 87.245 194.425 88.825 194.755 ;
        RECT 100.815 194.425 102.395 194.755 ;
        RECT 114.385 194.425 115.965 194.755 ;
        RECT 80.460 191.705 82.040 192.035 ;
        RECT 94.030 191.705 95.610 192.035 ;
        RECT 107.600 191.705 109.180 192.035 ;
        RECT 121.170 191.705 122.750 192.035 ;
        RECT 73.675 188.985 75.255 189.315 ;
        RECT 87.245 188.985 88.825 189.315 ;
        RECT 100.815 188.985 102.395 189.315 ;
        RECT 114.385 188.985 115.965 189.315 ;
        RECT 80.460 186.265 82.040 186.595 ;
        RECT 94.030 186.265 95.610 186.595 ;
        RECT 107.600 186.265 109.180 186.595 ;
        RECT 121.170 186.265 122.750 186.595 ;
        RECT 73.675 183.545 75.255 183.875 ;
        RECT 87.245 183.545 88.825 183.875 ;
        RECT 100.815 183.545 102.395 183.875 ;
        RECT 114.385 183.545 115.965 183.875 ;
        RECT 80.460 180.825 82.040 181.155 ;
        RECT 94.030 180.825 95.610 181.155 ;
        RECT 107.600 180.825 109.180 181.155 ;
        RECT 121.170 180.825 122.750 181.155 ;
        RECT 73.675 178.105 75.255 178.435 ;
        RECT 87.245 178.105 88.825 178.435 ;
        RECT 100.815 178.105 102.395 178.435 ;
        RECT 114.385 178.105 115.965 178.435 ;
        RECT 80.460 175.385 82.040 175.715 ;
        RECT 94.030 175.385 95.610 175.715 ;
        RECT 107.600 175.385 109.180 175.715 ;
        RECT 121.170 175.385 122.750 175.715 ;
        RECT 153.090 174.150 153.715 219.485 ;
        RECT 121.105 174.000 121.435 174.015 ;
        RECT 122.920 174.000 153.715 174.150 ;
        RECT 121.105 173.700 153.715 174.000 ;
        RECT 121.105 173.685 121.435 173.700 ;
        RECT 122.920 173.550 153.715 173.700 ;
        RECT 153.090 173.540 153.715 173.550 ;
        RECT 73.675 172.665 75.255 172.995 ;
        RECT 87.245 172.665 88.825 172.995 ;
        RECT 100.815 172.665 102.395 172.995 ;
        RECT 114.385 172.665 115.965 172.995 ;
        RECT 80.460 169.945 82.040 170.275 ;
        RECT 94.030 169.945 95.610 170.275 ;
        RECT 107.600 169.945 109.180 170.275 ;
        RECT 121.170 169.945 122.750 170.275 ;
        RECT 85.225 169.240 85.555 169.255 ;
        RECT 92.585 169.240 92.915 169.255 ;
        RECT 85.225 168.940 92.915 169.240 ;
        RECT 85.225 168.925 85.555 168.940 ;
        RECT 92.585 168.925 92.915 168.940 ;
        RECT 73.675 167.225 75.255 167.555 ;
        RECT 87.245 167.225 88.825 167.555 ;
        RECT 100.815 167.225 102.395 167.555 ;
        RECT 114.385 167.225 115.965 167.555 ;
        RECT 80.460 164.505 82.040 164.835 ;
        RECT 94.030 164.505 95.610 164.835 ;
        RECT 107.600 164.505 109.180 164.835 ;
        RECT 121.170 164.505 122.750 164.835 ;
        RECT 73.675 161.785 75.255 162.115 ;
        RECT 87.245 161.785 88.825 162.115 ;
        RECT 100.815 161.785 102.395 162.115 ;
        RECT 114.385 161.785 115.965 162.115 ;
        RECT 80.460 159.065 82.040 159.395 ;
        RECT 94.030 159.065 95.610 159.395 ;
        RECT 107.600 159.065 109.180 159.395 ;
        RECT 121.170 159.065 122.750 159.395 ;
        RECT 39.185 149.090 40.675 149.115 ;
        RECT 73.790 149.090 75.290 153.090 ;
        RECT 87.250 149.090 88.750 153.710 ;
        RECT 101.270 149.090 102.770 154.520 ;
        RECT 114.310 149.090 115.810 154.010 ;
        RECT 39.180 147.590 119.180 149.090 ;
        RECT 39.185 147.565 40.675 147.590 ;
        RECT 85.690 102.945 86.230 103.415 ;
        RECT 89.360 102.865 90.030 103.475 ;
        RECT 92.760 102.855 93.430 103.465 ;
        RECT 96.520 102.885 97.190 103.495 ;
        RECT 81.780 90.625 83.060 91.825 ;
        RECT 105.310 72.785 105.860 73.235 ;
      LAYER via3 ;
        RECT 154.680 221.660 155.280 222.260 ;
        RECT 80.490 213.470 80.810 213.790 ;
        RECT 80.890 213.470 81.210 213.790 ;
        RECT 81.290 213.470 81.610 213.790 ;
        RECT 81.690 213.470 82.010 213.790 ;
        RECT 94.060 213.470 94.380 213.790 ;
        RECT 94.460 213.470 94.780 213.790 ;
        RECT 94.860 213.470 95.180 213.790 ;
        RECT 95.260 213.470 95.580 213.790 ;
        RECT 107.630 213.470 107.950 213.790 ;
        RECT 108.030 213.470 108.350 213.790 ;
        RECT 108.430 213.470 108.750 213.790 ;
        RECT 108.830 213.470 109.150 213.790 ;
        RECT 121.200 213.470 121.520 213.790 ;
        RECT 121.600 213.470 121.920 213.790 ;
        RECT 122.000 213.470 122.320 213.790 ;
        RECT 122.400 213.470 122.720 213.790 ;
        RECT 73.705 210.750 74.025 211.070 ;
        RECT 74.105 210.750 74.425 211.070 ;
        RECT 74.505 210.750 74.825 211.070 ;
        RECT 74.905 210.750 75.225 211.070 ;
        RECT 87.275 210.750 87.595 211.070 ;
        RECT 87.675 210.750 87.995 211.070 ;
        RECT 88.075 210.750 88.395 211.070 ;
        RECT 88.475 210.750 88.795 211.070 ;
        RECT 100.845 210.750 101.165 211.070 ;
        RECT 101.245 210.750 101.565 211.070 ;
        RECT 101.645 210.750 101.965 211.070 ;
        RECT 102.045 210.750 102.365 211.070 ;
        RECT 114.415 210.750 114.735 211.070 ;
        RECT 114.815 210.750 115.135 211.070 ;
        RECT 115.215 210.750 115.535 211.070 ;
        RECT 115.615 210.750 115.935 211.070 ;
        RECT 80.490 208.030 80.810 208.350 ;
        RECT 80.890 208.030 81.210 208.350 ;
        RECT 81.290 208.030 81.610 208.350 ;
        RECT 81.690 208.030 82.010 208.350 ;
        RECT 94.060 208.030 94.380 208.350 ;
        RECT 94.460 208.030 94.780 208.350 ;
        RECT 94.860 208.030 95.180 208.350 ;
        RECT 95.260 208.030 95.580 208.350 ;
        RECT 107.630 208.030 107.950 208.350 ;
        RECT 108.030 208.030 108.350 208.350 ;
        RECT 108.430 208.030 108.750 208.350 ;
        RECT 108.830 208.030 109.150 208.350 ;
        RECT 121.200 208.030 121.520 208.350 ;
        RECT 121.600 208.030 121.920 208.350 ;
        RECT 122.000 208.030 122.320 208.350 ;
        RECT 122.400 208.030 122.720 208.350 ;
        RECT 73.705 205.310 74.025 205.630 ;
        RECT 74.105 205.310 74.425 205.630 ;
        RECT 74.505 205.310 74.825 205.630 ;
        RECT 74.905 205.310 75.225 205.630 ;
        RECT 87.275 205.310 87.595 205.630 ;
        RECT 87.675 205.310 87.995 205.630 ;
        RECT 88.075 205.310 88.395 205.630 ;
        RECT 88.475 205.310 88.795 205.630 ;
        RECT 100.845 205.310 101.165 205.630 ;
        RECT 101.245 205.310 101.565 205.630 ;
        RECT 101.645 205.310 101.965 205.630 ;
        RECT 102.045 205.310 102.365 205.630 ;
        RECT 114.415 205.310 114.735 205.630 ;
        RECT 114.815 205.310 115.135 205.630 ;
        RECT 115.215 205.310 115.535 205.630 ;
        RECT 115.615 205.310 115.935 205.630 ;
        RECT 80.490 202.590 80.810 202.910 ;
        RECT 80.890 202.590 81.210 202.910 ;
        RECT 81.290 202.590 81.610 202.910 ;
        RECT 81.690 202.590 82.010 202.910 ;
        RECT 94.060 202.590 94.380 202.910 ;
        RECT 94.460 202.590 94.780 202.910 ;
        RECT 94.860 202.590 95.180 202.910 ;
        RECT 95.260 202.590 95.580 202.910 ;
        RECT 107.630 202.590 107.950 202.910 ;
        RECT 108.030 202.590 108.350 202.910 ;
        RECT 108.430 202.590 108.750 202.910 ;
        RECT 108.830 202.590 109.150 202.910 ;
        RECT 121.200 202.590 121.520 202.910 ;
        RECT 121.600 202.590 121.920 202.910 ;
        RECT 122.000 202.590 122.320 202.910 ;
        RECT 122.400 202.590 122.720 202.910 ;
        RECT 73.705 199.870 74.025 200.190 ;
        RECT 74.105 199.870 74.425 200.190 ;
        RECT 74.505 199.870 74.825 200.190 ;
        RECT 74.905 199.870 75.225 200.190 ;
        RECT 87.275 199.870 87.595 200.190 ;
        RECT 87.675 199.870 87.995 200.190 ;
        RECT 88.075 199.870 88.395 200.190 ;
        RECT 88.475 199.870 88.795 200.190 ;
        RECT 100.845 199.870 101.165 200.190 ;
        RECT 101.245 199.870 101.565 200.190 ;
        RECT 101.645 199.870 101.965 200.190 ;
        RECT 102.045 199.870 102.365 200.190 ;
        RECT 114.415 199.870 114.735 200.190 ;
        RECT 114.815 199.870 115.135 200.190 ;
        RECT 115.215 199.870 115.535 200.190 ;
        RECT 115.615 199.870 115.935 200.190 ;
        RECT 80.490 197.150 80.810 197.470 ;
        RECT 80.890 197.150 81.210 197.470 ;
        RECT 81.290 197.150 81.610 197.470 ;
        RECT 81.690 197.150 82.010 197.470 ;
        RECT 94.060 197.150 94.380 197.470 ;
        RECT 94.460 197.150 94.780 197.470 ;
        RECT 94.860 197.150 95.180 197.470 ;
        RECT 95.260 197.150 95.580 197.470 ;
        RECT 107.630 197.150 107.950 197.470 ;
        RECT 108.030 197.150 108.350 197.470 ;
        RECT 108.430 197.150 108.750 197.470 ;
        RECT 108.830 197.150 109.150 197.470 ;
        RECT 121.200 197.150 121.520 197.470 ;
        RECT 121.600 197.150 121.920 197.470 ;
        RECT 122.000 197.150 122.320 197.470 ;
        RECT 122.400 197.150 122.720 197.470 ;
        RECT 73.705 194.430 74.025 194.750 ;
        RECT 74.105 194.430 74.425 194.750 ;
        RECT 74.505 194.430 74.825 194.750 ;
        RECT 74.905 194.430 75.225 194.750 ;
        RECT 87.275 194.430 87.595 194.750 ;
        RECT 87.675 194.430 87.995 194.750 ;
        RECT 88.075 194.430 88.395 194.750 ;
        RECT 88.475 194.430 88.795 194.750 ;
        RECT 100.845 194.430 101.165 194.750 ;
        RECT 101.245 194.430 101.565 194.750 ;
        RECT 101.645 194.430 101.965 194.750 ;
        RECT 102.045 194.430 102.365 194.750 ;
        RECT 114.415 194.430 114.735 194.750 ;
        RECT 114.815 194.430 115.135 194.750 ;
        RECT 115.215 194.430 115.535 194.750 ;
        RECT 115.615 194.430 115.935 194.750 ;
        RECT 80.490 191.710 80.810 192.030 ;
        RECT 80.890 191.710 81.210 192.030 ;
        RECT 81.290 191.710 81.610 192.030 ;
        RECT 81.690 191.710 82.010 192.030 ;
        RECT 94.060 191.710 94.380 192.030 ;
        RECT 94.460 191.710 94.780 192.030 ;
        RECT 94.860 191.710 95.180 192.030 ;
        RECT 95.260 191.710 95.580 192.030 ;
        RECT 107.630 191.710 107.950 192.030 ;
        RECT 108.030 191.710 108.350 192.030 ;
        RECT 108.430 191.710 108.750 192.030 ;
        RECT 108.830 191.710 109.150 192.030 ;
        RECT 121.200 191.710 121.520 192.030 ;
        RECT 121.600 191.710 121.920 192.030 ;
        RECT 122.000 191.710 122.320 192.030 ;
        RECT 122.400 191.710 122.720 192.030 ;
        RECT 73.705 188.990 74.025 189.310 ;
        RECT 74.105 188.990 74.425 189.310 ;
        RECT 74.505 188.990 74.825 189.310 ;
        RECT 74.905 188.990 75.225 189.310 ;
        RECT 87.275 188.990 87.595 189.310 ;
        RECT 87.675 188.990 87.995 189.310 ;
        RECT 88.075 188.990 88.395 189.310 ;
        RECT 88.475 188.990 88.795 189.310 ;
        RECT 100.845 188.990 101.165 189.310 ;
        RECT 101.245 188.990 101.565 189.310 ;
        RECT 101.645 188.990 101.965 189.310 ;
        RECT 102.045 188.990 102.365 189.310 ;
        RECT 114.415 188.990 114.735 189.310 ;
        RECT 114.815 188.990 115.135 189.310 ;
        RECT 115.215 188.990 115.535 189.310 ;
        RECT 115.615 188.990 115.935 189.310 ;
        RECT 80.490 186.270 80.810 186.590 ;
        RECT 80.890 186.270 81.210 186.590 ;
        RECT 81.290 186.270 81.610 186.590 ;
        RECT 81.690 186.270 82.010 186.590 ;
        RECT 94.060 186.270 94.380 186.590 ;
        RECT 94.460 186.270 94.780 186.590 ;
        RECT 94.860 186.270 95.180 186.590 ;
        RECT 95.260 186.270 95.580 186.590 ;
        RECT 107.630 186.270 107.950 186.590 ;
        RECT 108.030 186.270 108.350 186.590 ;
        RECT 108.430 186.270 108.750 186.590 ;
        RECT 108.830 186.270 109.150 186.590 ;
        RECT 121.200 186.270 121.520 186.590 ;
        RECT 121.600 186.270 121.920 186.590 ;
        RECT 122.000 186.270 122.320 186.590 ;
        RECT 122.400 186.270 122.720 186.590 ;
        RECT 73.705 183.550 74.025 183.870 ;
        RECT 74.105 183.550 74.425 183.870 ;
        RECT 74.505 183.550 74.825 183.870 ;
        RECT 74.905 183.550 75.225 183.870 ;
        RECT 87.275 183.550 87.595 183.870 ;
        RECT 87.675 183.550 87.995 183.870 ;
        RECT 88.075 183.550 88.395 183.870 ;
        RECT 88.475 183.550 88.795 183.870 ;
        RECT 100.845 183.550 101.165 183.870 ;
        RECT 101.245 183.550 101.565 183.870 ;
        RECT 101.645 183.550 101.965 183.870 ;
        RECT 102.045 183.550 102.365 183.870 ;
        RECT 114.415 183.550 114.735 183.870 ;
        RECT 114.815 183.550 115.135 183.870 ;
        RECT 115.215 183.550 115.535 183.870 ;
        RECT 115.615 183.550 115.935 183.870 ;
        RECT 80.490 180.830 80.810 181.150 ;
        RECT 80.890 180.830 81.210 181.150 ;
        RECT 81.290 180.830 81.610 181.150 ;
        RECT 81.690 180.830 82.010 181.150 ;
        RECT 94.060 180.830 94.380 181.150 ;
        RECT 94.460 180.830 94.780 181.150 ;
        RECT 94.860 180.830 95.180 181.150 ;
        RECT 95.260 180.830 95.580 181.150 ;
        RECT 107.630 180.830 107.950 181.150 ;
        RECT 108.030 180.830 108.350 181.150 ;
        RECT 108.430 180.830 108.750 181.150 ;
        RECT 108.830 180.830 109.150 181.150 ;
        RECT 121.200 180.830 121.520 181.150 ;
        RECT 121.600 180.830 121.920 181.150 ;
        RECT 122.000 180.830 122.320 181.150 ;
        RECT 122.400 180.830 122.720 181.150 ;
        RECT 73.705 178.110 74.025 178.430 ;
        RECT 74.105 178.110 74.425 178.430 ;
        RECT 74.505 178.110 74.825 178.430 ;
        RECT 74.905 178.110 75.225 178.430 ;
        RECT 87.275 178.110 87.595 178.430 ;
        RECT 87.675 178.110 87.995 178.430 ;
        RECT 88.075 178.110 88.395 178.430 ;
        RECT 88.475 178.110 88.795 178.430 ;
        RECT 100.845 178.110 101.165 178.430 ;
        RECT 101.245 178.110 101.565 178.430 ;
        RECT 101.645 178.110 101.965 178.430 ;
        RECT 102.045 178.110 102.365 178.430 ;
        RECT 114.415 178.110 114.735 178.430 ;
        RECT 114.815 178.110 115.135 178.430 ;
        RECT 115.215 178.110 115.535 178.430 ;
        RECT 115.615 178.110 115.935 178.430 ;
        RECT 80.490 175.390 80.810 175.710 ;
        RECT 80.890 175.390 81.210 175.710 ;
        RECT 81.290 175.390 81.610 175.710 ;
        RECT 81.690 175.390 82.010 175.710 ;
        RECT 94.060 175.390 94.380 175.710 ;
        RECT 94.460 175.390 94.780 175.710 ;
        RECT 94.860 175.390 95.180 175.710 ;
        RECT 95.260 175.390 95.580 175.710 ;
        RECT 107.630 175.390 107.950 175.710 ;
        RECT 108.030 175.390 108.350 175.710 ;
        RECT 108.430 175.390 108.750 175.710 ;
        RECT 108.830 175.390 109.150 175.710 ;
        RECT 121.200 175.390 121.520 175.710 ;
        RECT 121.600 175.390 121.920 175.710 ;
        RECT 122.000 175.390 122.320 175.710 ;
        RECT 122.400 175.390 122.720 175.710 ;
        RECT 73.705 172.670 74.025 172.990 ;
        RECT 74.105 172.670 74.425 172.990 ;
        RECT 74.505 172.670 74.825 172.990 ;
        RECT 74.905 172.670 75.225 172.990 ;
        RECT 87.275 172.670 87.595 172.990 ;
        RECT 87.675 172.670 87.995 172.990 ;
        RECT 88.075 172.670 88.395 172.990 ;
        RECT 88.475 172.670 88.795 172.990 ;
        RECT 100.845 172.670 101.165 172.990 ;
        RECT 101.245 172.670 101.565 172.990 ;
        RECT 101.645 172.670 101.965 172.990 ;
        RECT 102.045 172.670 102.365 172.990 ;
        RECT 114.415 172.670 114.735 172.990 ;
        RECT 114.815 172.670 115.135 172.990 ;
        RECT 115.215 172.670 115.535 172.990 ;
        RECT 115.615 172.670 115.935 172.990 ;
        RECT 80.490 169.950 80.810 170.270 ;
        RECT 80.890 169.950 81.210 170.270 ;
        RECT 81.290 169.950 81.610 170.270 ;
        RECT 81.690 169.950 82.010 170.270 ;
        RECT 94.060 169.950 94.380 170.270 ;
        RECT 94.460 169.950 94.780 170.270 ;
        RECT 94.860 169.950 95.180 170.270 ;
        RECT 95.260 169.950 95.580 170.270 ;
        RECT 107.630 169.950 107.950 170.270 ;
        RECT 108.030 169.950 108.350 170.270 ;
        RECT 108.430 169.950 108.750 170.270 ;
        RECT 108.830 169.950 109.150 170.270 ;
        RECT 121.200 169.950 121.520 170.270 ;
        RECT 121.600 169.950 121.920 170.270 ;
        RECT 122.000 169.950 122.320 170.270 ;
        RECT 122.400 169.950 122.720 170.270 ;
        RECT 73.705 167.230 74.025 167.550 ;
        RECT 74.105 167.230 74.425 167.550 ;
        RECT 74.505 167.230 74.825 167.550 ;
        RECT 74.905 167.230 75.225 167.550 ;
        RECT 87.275 167.230 87.595 167.550 ;
        RECT 87.675 167.230 87.995 167.550 ;
        RECT 88.075 167.230 88.395 167.550 ;
        RECT 88.475 167.230 88.795 167.550 ;
        RECT 100.845 167.230 101.165 167.550 ;
        RECT 101.245 167.230 101.565 167.550 ;
        RECT 101.645 167.230 101.965 167.550 ;
        RECT 102.045 167.230 102.365 167.550 ;
        RECT 114.415 167.230 114.735 167.550 ;
        RECT 114.815 167.230 115.135 167.550 ;
        RECT 115.215 167.230 115.535 167.550 ;
        RECT 115.615 167.230 115.935 167.550 ;
        RECT 80.490 164.510 80.810 164.830 ;
        RECT 80.890 164.510 81.210 164.830 ;
        RECT 81.290 164.510 81.610 164.830 ;
        RECT 81.690 164.510 82.010 164.830 ;
        RECT 94.060 164.510 94.380 164.830 ;
        RECT 94.460 164.510 94.780 164.830 ;
        RECT 94.860 164.510 95.180 164.830 ;
        RECT 95.260 164.510 95.580 164.830 ;
        RECT 107.630 164.510 107.950 164.830 ;
        RECT 108.030 164.510 108.350 164.830 ;
        RECT 108.430 164.510 108.750 164.830 ;
        RECT 108.830 164.510 109.150 164.830 ;
        RECT 121.200 164.510 121.520 164.830 ;
        RECT 121.600 164.510 121.920 164.830 ;
        RECT 122.000 164.510 122.320 164.830 ;
        RECT 122.400 164.510 122.720 164.830 ;
        RECT 73.705 161.790 74.025 162.110 ;
        RECT 74.105 161.790 74.425 162.110 ;
        RECT 74.505 161.790 74.825 162.110 ;
        RECT 74.905 161.790 75.225 162.110 ;
        RECT 87.275 161.790 87.595 162.110 ;
        RECT 87.675 161.790 87.995 162.110 ;
        RECT 88.075 161.790 88.395 162.110 ;
        RECT 88.475 161.790 88.795 162.110 ;
        RECT 100.845 161.790 101.165 162.110 ;
        RECT 101.245 161.790 101.565 162.110 ;
        RECT 101.645 161.790 101.965 162.110 ;
        RECT 102.045 161.790 102.365 162.110 ;
        RECT 114.415 161.790 114.735 162.110 ;
        RECT 114.815 161.790 115.135 162.110 ;
        RECT 115.215 161.790 115.535 162.110 ;
        RECT 115.615 161.790 115.935 162.110 ;
        RECT 80.490 159.070 80.810 159.390 ;
        RECT 80.890 159.070 81.210 159.390 ;
        RECT 81.290 159.070 81.610 159.390 ;
        RECT 81.690 159.070 82.010 159.390 ;
        RECT 94.060 159.070 94.380 159.390 ;
        RECT 94.460 159.070 94.780 159.390 ;
        RECT 94.860 159.070 95.180 159.390 ;
        RECT 95.260 159.070 95.580 159.390 ;
        RECT 107.630 159.070 107.950 159.390 ;
        RECT 108.030 159.070 108.350 159.390 ;
        RECT 108.430 159.070 108.750 159.390 ;
        RECT 108.830 159.070 109.150 159.390 ;
        RECT 121.200 159.070 121.520 159.390 ;
        RECT 121.600 159.070 121.920 159.390 ;
        RECT 122.000 159.070 122.320 159.390 ;
        RECT 122.400 159.070 122.720 159.390 ;
        RECT 73.790 151.560 75.290 153.060 ;
        RECT 87.250 152.180 88.750 153.680 ;
        RECT 101.270 152.990 102.770 154.490 ;
        RECT 114.310 152.480 115.810 153.980 ;
        RECT 39.185 147.595 40.675 149.085 ;
        RECT 85.740 102.970 86.180 103.390 ;
        RECT 89.410 102.890 89.980 103.450 ;
        RECT 92.810 102.880 93.380 103.440 ;
        RECT 96.570 102.910 97.140 103.470 ;
        RECT 81.830 90.650 83.010 91.800 ;
        RECT 105.360 72.810 105.810 73.210 ;
      LAYER met4 ;
        RECT 151.100 224.760 151.190 225.230 ;
        RECT 151.490 224.760 151.725 225.230 ;
        RECT 73.665 160.430 75.265 213.870 ;
        RECT 73.665 158.990 75.290 160.430 ;
        RECT 80.450 159.910 82.050 213.870 ;
        RECT 80.450 158.990 82.140 159.910 ;
        RECT 87.235 158.990 88.835 213.870 ;
        RECT 94.020 160.760 95.620 213.870 ;
        RECT 93.890 158.990 95.620 160.760 ;
        RECT 100.805 160.720 102.405 213.870 ;
        RECT 100.805 158.990 102.770 160.720 ;
        RECT 107.590 160.680 109.190 213.870 ;
        RECT 114.375 161.350 115.975 213.870 ;
        RECT 73.790 153.065 75.290 158.990 ;
        RECT 73.785 151.555 75.295 153.065 ;
        RECT 2.500 147.590 40.680 149.090 ;
        RECT 80.470 146.110 82.140 158.990 ;
        RECT 87.250 153.685 88.750 158.990 ;
        RECT 87.245 152.175 88.755 153.685 ;
        RECT 93.890 146.110 95.560 158.990 ;
        RECT 101.270 154.495 102.770 158.990 ;
        RECT 101.265 152.985 102.775 154.495 ;
        RECT 107.560 146.110 109.230 160.680 ;
        RECT 114.310 158.990 115.975 161.350 ;
        RECT 121.160 158.990 122.760 213.870 ;
        RECT 114.310 153.985 115.810 158.990 ;
        RECT 114.305 152.475 115.815 153.985 ;
        RECT 50.500 144.610 116.150 146.110 ;
        RECT 136.470 129.610 136.770 224.760 ;
        RECT 85.810 129.310 136.770 129.610 ;
        RECT 85.810 103.395 86.110 129.310 ;
        RECT 140.150 123.550 140.450 224.760 ;
        RECT 89.560 123.250 140.450 123.550 ;
        RECT 89.560 103.455 89.860 123.250 ;
        RECT 143.830 119.690 144.130 224.760 ;
        RECT 92.940 119.390 144.130 119.690 ;
        RECT 85.735 102.965 86.185 103.395 ;
        RECT 89.405 102.885 89.985 103.455 ;
        RECT 92.940 103.445 93.240 119.390 ;
        RECT 147.510 115.550 147.810 224.760 ;
        RECT 151.100 220.115 151.725 224.760 ;
        RECT 154.700 224.760 154.870 225.280 ;
        RECT 155.170 224.760 155.300 225.280 ;
        RECT 154.700 223.360 155.300 224.760 ;
        RECT 154.680 222.720 155.300 223.360 ;
        RECT 154.680 222.265 155.280 222.720 ;
        RECT 154.675 221.655 155.285 222.265 ;
        RECT 151.095 219.480 151.730 220.115 ;
        RECT 96.670 115.250 147.810 115.550 ;
        RECT 96.670 103.475 96.970 115.250 ;
        RECT 92.805 102.875 93.385 103.445 ;
        RECT 96.565 102.905 97.145 103.475 ;
        RECT 50.500 90.430 83.130 91.930 ;
        RECT 105.170 72.700 157.160 73.300 ;
        RECT 156.560 1.000 157.160 72.700 ;
  END
END tt_um_mattvenn_r2r_dac
END LIBRARY

