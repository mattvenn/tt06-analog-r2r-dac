magic
tech sky130A
magscale 1 2
timestamp 1708508486
<< metal1 >>
rect 22480 31060 22600 31066
rect 23474 31060 23480 31180
rect 23600 31060 23606 31180
rect 22600 30940 22920 31060
rect 22480 30934 22600 30940
rect 21400 29800 21520 29806
rect 21520 29680 22640 29800
rect 21400 29674 21520 29680
rect 21340 29340 21460 29346
rect 21460 29220 22320 29340
rect 21340 29214 21460 29220
rect 22520 29200 22640 29680
rect 22800 29220 22920 30940
rect 23174 30500 23180 30620
rect 23300 30500 23306 30620
rect 23180 29220 23300 30500
rect 23480 29200 23600 31060
rect 23774 31040 23780 31160
rect 23900 31040 23906 31160
rect 23780 29200 23900 31040
rect 24074 31020 24080 31140
rect 24200 31020 24206 31140
rect 24080 29240 24200 31020
rect 24354 30820 24360 30940
rect 24480 30820 24486 30940
rect 24360 29800 24480 30820
rect 24360 29680 24580 29800
rect 24460 29240 24580 29680
rect 24296 27666 25140 27866
rect 24943 6080 25138 27666
rect 24943 5583 25140 6080
rect 25020 5280 25140 5583
rect 26060 5280 26180 5286
rect 25020 5160 26060 5280
rect 26060 5154 26180 5160
<< via1 >>
rect 23480 31060 23600 31180
rect 22480 30940 22600 31060
rect 21400 29680 21520 29800
rect 21340 29220 21460 29340
rect 23180 30500 23300 30620
rect 23780 31040 23900 31160
rect 24080 31020 24200 31140
rect 24360 30820 24480 30940
rect 26060 5160 26180 5280
<< metal2 >>
rect 3948 44538 4008 44547
rect 3948 44469 4008 44478
rect 3950 41864 4006 44469
rect 5250 44339 5310 44341
rect 5243 44283 5252 44339
rect 5308 44283 5317 44339
rect 5250 41703 5310 44283
rect 6515 44089 6524 44149
rect 6584 44089 6593 44149
rect 6526 41737 6582 44089
rect 7809 43931 7869 43933
rect 7802 43875 7811 43931
rect 7867 43875 7876 43931
rect 7809 41727 7869 43875
rect 9096 43700 9152 43707
rect 9094 43698 9154 43700
rect 9094 43642 9096 43698
rect 9152 43642 9154 43698
rect 9094 41815 9154 43642
rect 10388 43452 10448 43461
rect 10388 43383 10448 43392
rect 10390 41801 10446 43383
rect 11680 43202 11740 43204
rect 11673 43146 11682 43202
rect 11738 43146 11747 43202
rect 11680 41767 11740 43146
rect 12964 43012 13024 43021
rect 12964 42943 13024 42952
rect 12966 41857 13022 42943
rect 14242 42786 14302 42788
rect 14235 42730 14244 42786
rect 14300 42730 14309 42786
rect 14242 41759 14302 42730
rect 15540 42594 15600 42603
rect 15540 42525 15600 42534
rect 15542 41897 15598 42525
rect 16826 42397 16886 42399
rect 16819 42341 16828 42397
rect 16884 42341 16893 42397
rect 16826 41835 16886 42341
rect 18107 42144 18116 42204
rect 18176 42144 18185 42204
rect 18118 41872 18174 42144
rect 23480 32335 23600 32340
rect 23476 32225 23485 32335
rect 23595 32225 23604 32335
rect 23180 31475 23300 31480
rect 23176 31365 23185 31475
rect 23295 31365 23304 31475
rect 21285 31060 21395 31064
rect 21280 31055 22480 31060
rect 21280 30945 21285 31055
rect 21395 30945 22480 31055
rect 21280 30940 22480 30945
rect 22600 30940 22606 31060
rect 21285 30936 21395 30940
rect 23180 30620 23300 31365
rect 23480 31180 23600 32225
rect 23780 32035 23900 32040
rect 23776 31925 23785 32035
rect 23895 31925 23904 32035
rect 23480 31054 23600 31060
rect 23780 31160 23900 31925
rect 24080 31815 24200 31820
rect 24076 31705 24085 31815
rect 24195 31705 24204 31815
rect 24360 31795 24480 31800
rect 23780 31034 23900 31040
rect 24080 31140 24200 31705
rect 24356 31685 24365 31795
rect 24475 31685 24484 31795
rect 24080 31014 24200 31020
rect 24360 30940 24480 31685
rect 24360 30814 24480 30820
rect 23180 30494 23300 30500
rect 20945 29800 21055 29804
rect 20940 29795 21400 29800
rect 20940 29685 20945 29795
rect 21055 29685 21400 29795
rect 20940 29680 21400 29685
rect 21520 29680 21526 29800
rect 20945 29676 21055 29680
rect 20945 29340 21055 29344
rect 20940 29335 21340 29340
rect 20940 29225 20945 29335
rect 21055 29225 21340 29335
rect 20940 29220 21340 29225
rect 21460 29220 21466 29340
rect 20945 29216 21055 29220
rect 29465 5280 29575 5284
rect 26054 5160 26060 5280
rect 26180 5275 29580 5280
rect 26180 5165 29465 5275
rect 29575 5165 29580 5275
rect 26180 5160 29580 5165
rect 29465 5156 29575 5160
<< via2 >>
rect 3948 44478 4008 44538
rect 5252 44283 5308 44339
rect 6524 44089 6584 44149
rect 7811 43875 7867 43931
rect 9096 43642 9152 43698
rect 10388 43392 10448 43452
rect 11682 43146 11738 43202
rect 12964 42952 13024 43012
rect 14244 42730 14300 42786
rect 15540 42534 15600 42594
rect 16828 42341 16884 42397
rect 18116 42144 18176 42204
rect 23485 32225 23595 32335
rect 23185 31365 23295 31475
rect 21285 30945 21395 31055
rect 23785 31925 23895 32035
rect 24085 31705 24195 31815
rect 24365 31685 24475 31795
rect 20945 29685 21055 29795
rect 20945 29225 21055 29335
rect 29465 5165 29575 5275
<< metal3 >>
rect 3943 44538 4013 44543
rect 22882 44540 22946 44546
rect 3943 44478 3948 44538
rect 4008 44478 22882 44538
rect 3943 44473 4013 44478
rect 22882 44470 22946 44476
rect 5247 44341 5313 44344
rect 23612 44343 23676 44349
rect 5247 44339 23612 44341
rect 5247 44283 5252 44339
rect 5308 44283 23612 44339
rect 5247 44281 23612 44283
rect 5247 44278 5313 44281
rect 23612 44273 23676 44279
rect 6519 44149 6589 44154
rect 24345 44151 24409 44157
rect 6519 44089 6524 44149
rect 6584 44089 24345 44149
rect 6519 44084 6589 44089
rect 24345 44081 24409 44087
rect 7806 43933 7872 43936
rect 25084 43935 25148 43941
rect 7806 43931 25084 43933
rect 7806 43875 7811 43931
rect 7867 43875 25084 43931
rect 7806 43873 25084 43875
rect 7806 43870 7872 43873
rect 25084 43865 25148 43871
rect 9091 43700 9157 43703
rect 25814 43700 25820 43702
rect 9091 43698 25820 43700
rect 9091 43642 9096 43698
rect 9152 43642 25820 43698
rect 9091 43640 25820 43642
rect 9091 43637 9157 43640
rect 25814 43638 25820 43640
rect 25884 43638 25890 43702
rect 10383 43452 10453 43457
rect 26552 43454 26616 43460
rect 10383 43392 10388 43452
rect 10448 43392 26552 43452
rect 10383 43387 10453 43392
rect 26552 43384 26616 43390
rect 11677 43204 11743 43207
rect 27292 43206 27356 43212
rect 11677 43202 27292 43204
rect 11677 43146 11682 43202
rect 11738 43146 27292 43202
rect 11677 43144 27292 43146
rect 11677 43141 11743 43144
rect 27292 43136 27356 43142
rect 12959 43012 13029 43017
rect 28018 43012 28024 43014
rect 12959 42952 12964 43012
rect 13024 42952 28024 43012
rect 12959 42947 13029 42952
rect 28018 42950 28024 42952
rect 28088 42950 28094 43014
rect 14239 42788 14305 42791
rect 28764 42790 28828 42796
rect 14239 42786 28764 42788
rect 14239 42730 14244 42786
rect 14300 42730 28764 42786
rect 14239 42728 28764 42730
rect 14239 42725 14305 42728
rect 28764 42720 28828 42726
rect 15535 42594 15605 42599
rect 29486 42594 29492 42596
rect 15535 42534 15540 42594
rect 15600 42534 29492 42594
rect 15535 42529 15605 42534
rect 29486 42532 29492 42534
rect 29556 42532 29562 42596
rect 16823 42399 16889 42402
rect 30236 42401 30300 42407
rect 16823 42397 30236 42399
rect 16823 42341 16828 42397
rect 16884 42341 30236 42397
rect 16823 42339 30236 42341
rect 16823 42336 16889 42339
rect 30236 42331 30300 42337
rect 18111 42204 18181 42209
rect 30973 42206 31037 42212
rect 18111 42144 18116 42204
rect 18176 42144 30973 42204
rect 18111 42139 18181 42144
rect 30973 42136 31037 42142
rect 18840 40460 24480 40580
rect 18880 38556 24200 38676
rect 18840 36652 23900 36772
rect 18840 34748 23600 34868
rect 18860 32844 23300 32964
rect 23180 31475 23300 32844
rect 23480 32335 23600 34748
rect 23480 32225 23485 32335
rect 23595 32225 23600 32335
rect 23480 32220 23600 32225
rect 23780 32035 23900 36652
rect 23780 31925 23785 32035
rect 23895 31925 23900 32035
rect 23780 31920 23900 31925
rect 24080 31815 24200 38556
rect 24080 31705 24085 31815
rect 24195 31705 24200 31815
rect 24080 31700 24200 31705
rect 24360 31795 24480 40460
rect 24360 31685 24365 31795
rect 24475 31685 24480 31795
rect 24360 31680 24480 31685
rect 23180 31365 23185 31475
rect 23295 31365 23300 31475
rect 23180 31360 23300 31365
rect 18960 31055 21400 31060
rect 18960 30945 21285 31055
rect 21395 30945 21400 31055
rect 18960 30940 21400 30945
rect 19820 29795 21060 29800
rect 19820 29685 20945 29795
rect 21055 29685 21060 29795
rect 19820 29680 21060 29685
rect 19820 29156 19940 29680
rect 18920 29036 19940 29156
rect 20940 29335 21060 29340
rect 20940 29225 20945 29335
rect 21055 29225 21060 29335
rect 20940 27252 21060 29225
rect 18940 27132 21060 27252
rect 5310 25300 5630 25306
rect 12760 25300 13080 25306
rect 182 24980 188 25300
rect 508 24980 5310 25300
rect 5630 24980 9056 25300
rect 9376 24980 12760 25300
rect 13080 24980 16450 25300
rect 16770 24980 16780 25300
rect 5310 24974 5630 24980
rect 12760 24974 13080 24980
rect 31313 5280 31431 5285
rect 29460 5279 31432 5280
rect 29460 5275 31313 5279
rect 29460 5165 29465 5275
rect 29575 5165 31313 5275
rect 29460 5161 31313 5165
rect 31431 5161 31432 5279
rect 29460 5160 31432 5161
rect 31313 5155 31431 5160
<< via3 >>
rect 22882 44476 22946 44540
rect 23612 44279 23676 44343
rect 24345 44087 24409 44151
rect 25084 43871 25148 43935
rect 25820 43638 25884 43702
rect 26552 43390 26616 43454
rect 27292 43142 27356 43206
rect 28024 42950 28088 43014
rect 28764 42726 28828 42790
rect 29492 42532 29556 42596
rect 30236 42337 30300 42401
rect 30973 42142 31037 42206
rect 188 24980 508 25300
rect 5310 24980 5630 25300
rect 9056 24980 9376 25300
rect 12760 24980 13080 25300
rect 16450 24980 16770 25300
rect 31313 5161 31431 5279
<< metal4 >>
rect 22884 45152 22944 45158
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44723 5274 45152
rect 5950 44723 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22944 45152
rect 3547 44663 6010 44723
rect 200 25301 500 44152
rect 1688 43545 1988 44256
rect 3547 43545 3607 44663
rect 22884 44541 22944 44952
rect 22881 44540 22947 44541
rect 22881 44476 22882 44540
rect 22946 44476 22947 44540
rect 22881 44475 22947 44476
rect 23614 44344 23674 45152
rect 24350 45117 24410 45152
rect 24347 44952 24410 45117
rect 23611 44343 23677 44344
rect 23611 44279 23612 44343
rect 23676 44279 23677 44343
rect 23611 44278 23677 44279
rect 24347 44152 24407 44952
rect 24344 44151 24410 44152
rect 24344 44087 24345 44151
rect 24409 44087 24410 44151
rect 24344 44086 24410 44087
rect 25086 43936 25146 45152
rect 25083 43935 25149 43936
rect 25083 43871 25084 43935
rect 25148 43871 25149 43935
rect 25083 43870 25149 43871
rect 25822 43703 25882 45152
rect 26558 45117 26618 45152
rect 26554 44952 26618 45117
rect 25819 43702 25885 43703
rect 25819 43638 25820 43702
rect 25884 43638 25885 43702
rect 25819 43637 25885 43638
rect 1668 43485 3607 43545
rect 187 25300 509 25301
rect 187 24980 188 25300
rect 508 24980 510 25300
rect 187 24979 509 24980
rect 200 1000 500 24979
rect 1688 24290 1988 43485
rect 26554 43455 26614 44952
rect 26551 43454 26617 43455
rect 26551 43390 26552 43454
rect 26616 43390 26617 43454
rect 26551 43389 26617 43390
rect 27294 43207 27354 45152
rect 28030 45117 28090 45152
rect 28026 44952 28090 45117
rect 27291 43206 27357 43207
rect 27291 43142 27292 43206
rect 27356 43142 27357 43206
rect 27291 43141 27357 43142
rect 28026 43015 28086 44952
rect 28023 43014 28089 43015
rect 28023 42950 28024 43014
rect 28088 42950 28089 43014
rect 28023 42949 28089 42950
rect 28766 42791 28826 45152
rect 29502 45125 29562 45152
rect 29494 44952 29562 45125
rect 28763 42790 28829 42791
rect 28763 42726 28764 42790
rect 28828 42726 28829 42790
rect 28763 42725 28829 42726
rect 29494 42597 29554 44952
rect 29491 42596 29557 42597
rect 29491 42532 29492 42596
rect 29556 42532 29557 42596
rect 29491 42531 29557 42532
rect 30238 42402 30298 45152
rect 30974 45074 31034 45152
rect 30974 44952 31035 45074
rect 31710 44952 31770 45152
rect 30235 42401 30301 42402
rect 30235 42337 30236 42401
rect 30300 42337 30301 42401
rect 30235 42336 30301 42337
rect 30975 42207 31035 44952
rect 30972 42206 31038 42207
rect 30972 42142 30973 42206
rect 31037 42142 31038 42206
rect 30972 42141 31038 42142
rect 5310 25301 5630 27340
rect 5309 25300 5631 25301
rect 5309 24980 5310 25300
rect 5630 24980 5631 25300
rect 5309 24979 5631 24980
rect 7190 24290 7490 27070
rect 9056 25301 9376 27418
rect 9055 25300 9377 25301
rect 9055 24980 9056 25300
rect 9376 24980 9377 25300
rect 9055 24979 9377 24980
rect 10930 24290 11230 27110
rect 12760 25301 13080 27494
rect 12759 25300 13081 25301
rect 12759 24980 12760 25300
rect 13080 24980 13081 25300
rect 12759 24979 13081 24980
rect 14590 24290 14890 27170
rect 16450 25301 16770 27550
rect 16449 25300 16771 25301
rect 16449 24980 16450 25300
rect 16770 24980 16771 25300
rect 16449 24979 16771 24980
rect 1688 23990 18790 24290
rect 1688 1104 1988 23990
rect 31312 5279 31432 5280
rect 31312 5161 31313 5279
rect 31431 5161 31432 5279
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31312 0 31432 5161
use r2r  r2r_0
timestamp 1708461036
transform 1 0 21996 0 1 27306
box 160 -600 2600 2080
use r2r_dac_control  r2r_dac_control_0
timestamp 1708507682
transform 1 0 3104 0 1 26036
box 514 496 16000 16000
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 1688 1104 1988 44256 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
